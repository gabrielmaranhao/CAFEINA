magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< nwell >>
rect 9324 -4370 23581 -2602
rect 9079 -9662 23581 -4370
rect 9079 -18334 18105 -9662
<< locali >>
rect 6981 16254 7043 16432
rect 7221 16254 7275 16432
rect 6981 16209 7275 16254
rect 7480 16254 7542 16432
rect 7720 16254 7774 16432
rect 7480 16209 7774 16254
rect 7978 16254 8040 16432
rect 8218 16254 8272 16432
rect 7978 16209 8272 16254
rect 28407 16254 28469 16432
rect 28647 16254 28701 16432
rect 28407 16209 28701 16254
rect 28905 16254 28967 16432
rect 29145 16254 29199 16432
rect 28905 16209 29199 16254
rect 54121 -4756 54345 -4694
rect 54121 -4934 54166 -4756
rect 54272 -4790 54311 -4756
rect 54272 -4828 54345 -4790
rect 54272 -4862 54311 -4828
rect 54272 -4900 54345 -4862
rect 54272 -4934 54311 -4900
rect 54121 -4988 54345 -4934
rect 54138 -5304 54362 -5242
rect 54138 -5482 54183 -5304
rect 54289 -5338 54328 -5304
rect 54289 -5376 54362 -5338
rect 54289 -5410 54328 -5376
rect 54289 -5448 54362 -5410
rect 54289 -5482 54328 -5448
rect 54138 -5536 54362 -5482
rect 52204 -15074 52428 -15012
rect 52204 -15252 52249 -15074
rect 52355 -15108 52394 -15074
rect 52355 -15146 52428 -15108
rect 52355 -15180 52394 -15146
rect 52355 -15218 52428 -15180
rect 52355 -15252 52394 -15218
rect 52204 -15306 52428 -15252
<< viali >>
rect 6981 16596 7015 16630
rect 7241 16596 7275 16630
rect 7480 16596 7514 16630
rect 7740 16596 7774 16630
rect 7978 16596 8012 16630
rect 8238 16596 8272 16630
rect 28407 16596 28441 16630
rect 28667 16596 28701 16630
rect 28905 16596 28939 16630
rect 29165 16596 29199 16630
rect 6981 16524 7015 16558
rect 7241 16524 7275 16558
rect 7480 16524 7514 16558
rect 7740 16524 7774 16558
rect 7978 16524 8012 16558
rect 8238 16524 8272 16558
rect 28407 16524 28441 16558
rect 28667 16524 28701 16558
rect 28905 16524 28939 16558
rect 29165 16524 29199 16558
rect 7043 16254 7221 16432
rect 7542 16254 7720 16432
rect 8040 16254 8218 16432
rect 28469 16254 28647 16432
rect 28967 16254 29145 16432
rect 54436 -4728 54470 -4694
rect 54509 -4728 54543 -4694
rect 54166 -4934 54272 -4756
rect 54311 -4790 54345 -4756
rect 54311 -4862 54345 -4828
rect 54311 -4934 54345 -4900
rect 54436 -4988 54470 -4954
rect 54509 -4988 54543 -4954
rect 54453 -5276 54487 -5242
rect 54526 -5276 54560 -5242
rect 54183 -5482 54289 -5304
rect 54328 -5338 54362 -5304
rect 54328 -5410 54362 -5376
rect 54328 -5482 54362 -5448
rect 54453 -5536 54487 -5502
rect 54526 -5536 54560 -5502
rect 52519 -15046 52553 -15012
rect 52592 -15046 52626 -15012
rect 52249 -15252 52355 -15074
rect 52394 -15108 52428 -15074
rect 52394 -15180 52428 -15146
rect 52394 -15252 52428 -15218
rect 52519 -15306 52553 -15272
rect 52592 -15306 52626 -15272
<< metal1 >>
rect 6990 17301 7266 17307
rect 6990 17121 7005 17301
rect 7249 17121 7266 17301
rect 6990 17081 7266 17121
rect 6990 16965 7038 17081
rect 7218 16965 7266 17081
rect 6990 16935 7266 16965
rect 7490 17301 7766 17307
rect 7490 17121 7502 17301
rect 7746 17121 7766 17301
rect 7490 17081 7766 17121
rect 7490 16965 7535 17081
rect 7715 16965 7766 17081
rect 7490 16935 7766 16965
rect 7988 17301 8264 17307
rect 7988 17121 7999 17301
rect 8243 17121 8264 17301
rect 7988 17081 8264 17121
rect 7988 16965 8033 17081
rect 8213 16965 8264 17081
rect 7988 16935 8264 16965
rect 28417 17301 28693 17307
rect 28417 17121 28429 17301
rect 28673 17121 28693 17301
rect 28417 17081 28693 17121
rect 28417 16965 28462 17081
rect 28642 16965 28693 17081
rect 28417 16935 28693 16965
rect 28915 17301 29191 17307
rect 28915 17121 28927 17301
rect 29171 17121 29191 17301
rect 28915 17081 29191 17121
rect 28915 16965 28960 17081
rect 29140 16965 29191 17081
rect 28915 16935 29191 16965
rect 7020 16754 7244 16935
rect 7520 16754 7744 16935
rect 8018 16754 8242 16935
rect 28447 16754 28671 16935
rect 28945 16754 29169 16935
rect 6963 16630 7031 16656
rect 6963 16596 6981 16630
rect 7015 16596 7031 16630
rect 6963 16558 7031 16596
rect 6963 16524 6981 16558
rect 7015 16524 7031 16558
rect 7089 16555 7167 16754
rect 7221 16630 7292 16656
rect 7221 16596 7241 16630
rect 7275 16596 7292 16630
rect 7221 16558 7292 16596
rect 6963 16441 7031 16524
rect 7221 16524 7241 16558
rect 7275 16524 7292 16558
rect 7221 16441 7292 16524
rect 6963 16432 7292 16441
rect 6963 16254 7043 16432
rect 7221 16254 7292 16432
rect 6963 16181 7292 16254
rect 7462 16630 7531 16656
rect 7462 16596 7480 16630
rect 7514 16596 7531 16630
rect 7462 16558 7531 16596
rect 7462 16524 7480 16558
rect 7514 16524 7531 16558
rect 7588 16555 7666 16754
rect 7721 16630 7791 16656
rect 7721 16596 7740 16630
rect 7774 16596 7791 16630
rect 7721 16558 7791 16596
rect 7462 16441 7531 16524
rect 7721 16524 7740 16558
rect 7774 16524 7791 16558
rect 7721 16441 7791 16524
rect 7462 16432 7791 16441
rect 7462 16254 7542 16432
rect 7720 16254 7791 16432
rect 7462 16181 7791 16254
rect 7960 16630 8028 16656
rect 7960 16596 7978 16630
rect 8012 16596 8028 16630
rect 7960 16558 8028 16596
rect 7960 16524 7978 16558
rect 8012 16524 8028 16558
rect 8086 16555 8164 16754
rect 8219 16630 8289 16656
rect 8219 16596 8238 16630
rect 8272 16596 8289 16630
rect 8219 16558 8289 16596
rect 7960 16441 8028 16524
rect 8219 16524 8238 16558
rect 8272 16524 8289 16558
rect 8219 16441 8289 16524
rect 7960 16432 8289 16441
rect 7960 16254 8040 16432
rect 8218 16254 8289 16432
rect 7960 16181 8289 16254
rect 28389 16630 28458 16656
rect 28389 16596 28407 16630
rect 28441 16596 28458 16630
rect 28389 16558 28458 16596
rect 28389 16524 28407 16558
rect 28441 16524 28458 16558
rect 28515 16555 28593 16754
rect 28648 16630 28718 16656
rect 28648 16596 28667 16630
rect 28701 16596 28718 16630
rect 28648 16558 28718 16596
rect 28389 16441 28458 16524
rect 28648 16524 28667 16558
rect 28701 16524 28718 16558
rect 28648 16441 28718 16524
rect 28389 16432 28718 16441
rect 28389 16254 28469 16432
rect 28647 16254 28718 16432
rect 28389 16181 28718 16254
rect 28887 16630 28956 16656
rect 28887 16596 28905 16630
rect 28939 16596 28956 16630
rect 28887 16558 28956 16596
rect 28887 16524 28905 16558
rect 28939 16524 28956 16558
rect 29013 16555 29091 16754
rect 29146 16630 29216 16656
rect 29146 16596 29165 16630
rect 29199 16596 29216 16630
rect 29146 16558 29216 16596
rect 28887 16441 28956 16524
rect 29146 16524 29165 16558
rect 29199 16524 29216 16558
rect 29146 16441 29216 16524
rect 28887 16432 29216 16441
rect 28887 16254 28967 16432
rect 29145 16254 29216 16432
rect 28887 16181 29216 16254
rect 6960 16112 52392 16181
rect 6960 15868 35382 16112
rect 35690 15868 35789 16112
rect 36097 15868 36177 16112
rect 36485 15868 36610 16112
rect 36918 15868 37017 16112
rect 37325 15868 37405 16112
rect 37713 15868 37812 16112
rect 38120 15868 38240 16112
rect 38548 15868 38646 16112
rect 38954 15868 39035 16112
rect 39343 15868 39441 16112
rect 39749 15868 39947 16112
rect 40255 15868 40354 16112
rect 40662 15868 40742 16112
rect 41050 15868 41149 16112
rect 41457 15868 41577 16112
rect 41885 15868 41984 16112
rect 42292 15868 42372 16112
rect 42680 15868 42779 16112
rect 43087 15868 43233 16112
rect 43541 15868 43639 16112
rect 43947 15868 44028 16112
rect 44336 15868 44434 16112
rect 44742 15868 44862 16112
rect 45170 15868 45269 16112
rect 45577 15868 45657 16112
rect 45965 15868 46064 16112
rect 46372 15868 46570 16112
rect 46878 15868 46977 16112
rect 47285 15868 47365 16112
rect 47673 15868 47772 16112
rect 48080 15868 48200 16112
rect 48508 15868 48607 16112
rect 48915 15868 48995 16112
rect 49303 15868 49402 16112
rect 49710 15868 49929 16112
rect 50237 15868 50357 16112
rect 50665 15868 50764 16112
rect 51072 15868 51152 16112
rect 51460 15868 51559 16112
rect 51867 15868 51997 16112
rect 52305 15868 52392 16112
rect 6960 15821 52392 15868
rect 9110 15514 51533 15587
rect 9110 15437 35291 15514
rect 35599 15437 35698 15514
rect 36006 15437 36086 15514
rect 36394 15437 36493 15514
rect 36801 15437 36921 15514
rect 37229 15437 37328 15514
rect 37636 15437 37716 15514
rect 38024 15437 38123 15514
rect 38431 15437 38628 15514
rect 38936 15437 39035 15514
rect 39343 15437 39423 15514
rect 39731 15437 39830 15514
rect 40138 15437 40258 15514
rect 40566 15437 40665 15514
rect 40973 15437 41053 15514
rect 41361 15437 41460 15514
rect 41768 15437 41914 15514
rect 42222 15437 42321 15514
rect 42629 15437 42709 15514
rect 43017 15437 43116 15514
rect 43424 15437 43544 15514
rect 43852 15437 43950 15514
rect 44258 15437 44339 15514
rect 44647 15437 44745 15514
rect 45053 15437 45251 15514
rect 45559 15437 45658 15514
rect 45966 15437 46046 15514
rect 46354 15437 46453 15514
rect 46761 15437 46881 15514
rect 47189 15437 47288 15514
rect 47596 15437 47676 15514
rect 47984 15437 48083 15514
rect 48391 15437 48610 15514
rect 48918 15437 49038 15514
rect 49346 15437 49445 15514
rect 49753 15437 49833 15514
rect 50141 15437 50240 15514
rect 50548 15437 51533 15514
rect 9110 -6967 23539 -3934
rect 51894 -4676 52392 15821
rect 51894 -4694 54568 -4676
rect 51894 -4728 54436 -4694
rect 54470 -4728 54509 -4694
rect 54543 -4728 54568 -4694
rect 51894 -4744 54568 -4728
rect 54848 -4715 55220 -4703
rect 54848 -4733 55033 -4715
rect 51894 -4756 54354 -4744
rect 51894 -4934 54166 -4756
rect 54272 -4790 54311 -4756
rect 54345 -4790 54354 -4756
rect 54272 -4828 54354 -4790
rect 54666 -4748 55033 -4733
rect 54666 -4802 54878 -4748
rect 54272 -4862 54311 -4828
rect 54345 -4862 54354 -4828
rect 54272 -4900 54354 -4862
rect 54468 -4880 54878 -4802
rect 54272 -4934 54311 -4900
rect 54345 -4934 54354 -4900
rect 54666 -4928 54878 -4880
rect 54994 -4928 55033 -4748
rect 51894 -4954 54568 -4934
rect 51894 -4988 54436 -4954
rect 54470 -4988 54509 -4954
rect 54543 -4988 54568 -4954
rect 54666 -4957 55033 -4928
rect 54848 -4959 55033 -4957
rect 55213 -4959 55220 -4715
rect 54848 -4979 55220 -4959
rect 51894 -5005 54568 -4988
rect 51894 -5224 52392 -5005
rect 51894 -5242 54585 -5224
rect 51894 -5276 54453 -5242
rect 54487 -5276 54526 -5242
rect 54560 -5276 54585 -5242
rect 51894 -5293 54585 -5276
rect 54865 -5264 55237 -5252
rect 54865 -5282 55050 -5264
rect 51894 -5304 54371 -5293
rect 51894 -5482 54183 -5304
rect 54289 -5338 54328 -5304
rect 54362 -5338 54371 -5304
rect 54289 -5376 54371 -5338
rect 54683 -5297 55050 -5282
rect 54683 -5350 54895 -5297
rect 54289 -5410 54328 -5376
rect 54362 -5410 54371 -5376
rect 54289 -5448 54371 -5410
rect 54485 -5428 54895 -5350
rect 54289 -5482 54328 -5448
rect 54362 -5482 54371 -5448
rect 51894 -5483 54371 -5482
rect 54683 -5477 54895 -5428
rect 55011 -5477 55050 -5297
rect 51894 -5502 54585 -5483
rect 51894 -5536 54453 -5502
rect 54487 -5536 54526 -5502
rect 54560 -5536 54585 -5502
rect 54683 -5506 55050 -5477
rect 54865 -5508 55050 -5506
rect 55230 -5508 55237 -5264
rect 54865 -5528 55237 -5508
rect 51894 -5553 54585 -5536
rect 51894 -5838 52392 -5553
rect 9110 -18307 12319 -6967
rect 24641 -14462 32110 -10798
rect 18726 -14481 32110 -14462
rect 51270 -14481 52392 -5838
rect 18726 -14994 52392 -14481
rect 18726 -15012 52651 -14994
rect 18726 -15046 52519 -15012
rect 52553 -15046 52592 -15012
rect 52626 -15046 52651 -15012
rect 18726 -15062 52651 -15046
rect 52931 -15033 53303 -15021
rect 52931 -15051 53116 -15033
rect 18726 -15074 52437 -15062
rect 18726 -15252 52249 -15074
rect 52355 -15108 52394 -15074
rect 52428 -15108 52437 -15074
rect 52355 -15146 52437 -15108
rect 52749 -15066 53116 -15051
rect 52749 -15120 52961 -15066
rect 52355 -15180 52394 -15146
rect 52428 -15180 52437 -15146
rect 52355 -15218 52437 -15180
rect 52568 -15198 52961 -15120
rect 52355 -15252 52394 -15218
rect 52428 -15252 52437 -15218
rect 52749 -15246 52961 -15198
rect 53077 -15246 53116 -15066
rect 18726 -15272 52651 -15252
rect 18726 -15306 52519 -15272
rect 52553 -15306 52592 -15272
rect 52626 -15306 52651 -15272
rect 52749 -15275 53116 -15246
rect 52931 -15277 53116 -15275
rect 53296 -15277 53303 -15033
rect 52931 -15297 53303 -15277
rect 18726 -15323 52651 -15306
rect 18726 -15324 52392 -15323
rect 18726 -16569 22499 -15324
rect 24621 -16569 52392 -15324
<< via1 >>
rect 7005 17121 7249 17301
rect 7038 16965 7218 17081
rect 7502 17121 7746 17301
rect 7535 16965 7715 17081
rect 7999 17121 8243 17301
rect 8033 16965 8213 17081
rect 28429 17121 28673 17301
rect 28462 16965 28642 17081
rect 28927 17121 29171 17301
rect 28960 16965 29140 17081
rect 35382 15868 35690 16112
rect 35789 15868 36097 16112
rect 36177 15868 36485 16112
rect 36610 15868 36918 16112
rect 37017 15868 37325 16112
rect 37405 15868 37713 16112
rect 37812 15868 38120 16112
rect 38240 15868 38548 16112
rect 38646 15868 38954 16112
rect 39035 15868 39343 16112
rect 39441 15868 39749 16112
rect 39947 15868 40255 16112
rect 40354 15868 40662 16112
rect 40742 15868 41050 16112
rect 41149 15868 41457 16112
rect 41577 15868 41885 16112
rect 41984 15868 42292 16112
rect 42372 15868 42680 16112
rect 42779 15868 43087 16112
rect 43233 15868 43541 16112
rect 43639 15868 43947 16112
rect 44028 15868 44336 16112
rect 44434 15868 44742 16112
rect 44862 15868 45170 16112
rect 45269 15868 45577 16112
rect 45657 15868 45965 16112
rect 46064 15868 46372 16112
rect 46570 15868 46878 16112
rect 46977 15868 47285 16112
rect 47365 15868 47673 16112
rect 47772 15868 48080 16112
rect 48200 15868 48508 16112
rect 48607 15868 48915 16112
rect 48995 15868 49303 16112
rect 49402 15868 49710 16112
rect 49929 15868 50237 16112
rect 50357 15868 50665 16112
rect 50764 15868 51072 16112
rect 51152 15868 51460 16112
rect 51559 15868 51867 16112
rect 51997 15868 52305 16112
rect 35291 15270 35599 15514
rect 35698 15270 36006 15514
rect 36086 15270 36394 15514
rect 36493 15270 36801 15514
rect 36921 15270 37229 15514
rect 37328 15270 37636 15514
rect 37716 15270 38024 15514
rect 38123 15270 38431 15514
rect 38628 15270 38936 15514
rect 39035 15270 39343 15514
rect 39423 15270 39731 15514
rect 39830 15270 40138 15514
rect 40258 15270 40566 15514
rect 40665 15270 40973 15514
rect 41053 15270 41361 15514
rect 41460 15270 41768 15514
rect 41914 15270 42222 15514
rect 42321 15270 42629 15514
rect 42709 15270 43017 15514
rect 43116 15270 43424 15514
rect 43544 15270 43852 15514
rect 43950 15270 44258 15514
rect 44339 15270 44647 15514
rect 44745 15270 45053 15514
rect 45251 15270 45559 15514
rect 45658 15270 45966 15514
rect 46046 15270 46354 15514
rect 46453 15270 46761 15514
rect 46881 15270 47189 15514
rect 47288 15270 47596 15514
rect 47676 15270 47984 15514
rect 48083 15270 48391 15514
rect 48610 15270 48918 15514
rect 49038 15270 49346 15514
rect 49445 15270 49753 15514
rect 49833 15270 50141 15514
rect 50240 15270 50548 15514
rect 54878 -4928 54994 -4748
rect 55033 -4959 55213 -4715
rect 54895 -5477 55011 -5297
rect 55050 -5508 55230 -5264
rect 52961 -15246 53077 -15066
rect 53116 -15277 53296 -15033
<< metal2 >>
rect 6977 17301 7277 17460
rect 6977 17121 7005 17301
rect 7249 17121 7277 17301
rect 6977 17109 7277 17121
rect 6977 17053 7021 17109
rect 7077 17081 7101 17109
rect 7157 17081 7181 17109
rect 7237 17053 7277 17109
rect 6977 17009 7038 17053
rect 7218 17009 7277 17053
rect 6977 16953 7021 17009
rect 7077 16953 7101 16965
rect 7157 16953 7181 16965
rect 7237 16953 7277 17009
rect 6977 16931 7277 16953
rect 7477 17301 7777 17460
rect 7477 17121 7502 17301
rect 7746 17121 7777 17301
rect 7477 17109 7777 17121
rect 7477 17053 7521 17109
rect 7577 17081 7601 17109
rect 7657 17081 7681 17109
rect 7737 17053 7777 17109
rect 7477 17009 7535 17053
rect 7715 17009 7777 17053
rect 7477 16953 7521 17009
rect 7577 16953 7601 16965
rect 7657 16953 7681 16965
rect 7737 16953 7777 17009
rect 7477 16931 7777 16953
rect 7976 17301 8276 17460
rect 7976 17121 7999 17301
rect 8243 17121 8276 17301
rect 7976 17109 8276 17121
rect 7976 17053 8020 17109
rect 8076 17081 8100 17109
rect 8156 17081 8180 17109
rect 8236 17053 8276 17109
rect 7976 17009 8033 17053
rect 8213 17009 8276 17053
rect 7976 16953 8020 17009
rect 8076 16953 8100 16965
rect 8156 16953 8180 16965
rect 8236 16953 8276 17009
rect 7976 16931 8276 16953
rect 28404 17301 28704 17460
rect 28404 17121 28429 17301
rect 28673 17121 28704 17301
rect 28404 17109 28704 17121
rect 28404 17053 28448 17109
rect 28504 17081 28528 17109
rect 28584 17081 28608 17109
rect 28664 17053 28704 17109
rect 28404 17009 28462 17053
rect 28642 17009 28704 17053
rect 28404 16953 28448 17009
rect 28504 16953 28528 16965
rect 28584 16953 28608 16965
rect 28664 16953 28704 17009
rect 28404 16931 28704 16953
rect 28903 17301 29203 17460
rect 28903 17121 28927 17301
rect 29171 17121 29203 17301
rect 28903 17109 29203 17121
rect 28903 17053 28947 17109
rect 29003 17081 29027 17109
rect 29083 17081 29107 17109
rect 29163 17053 29203 17109
rect 28903 17009 28960 17053
rect 29140 17009 29203 17053
rect 28903 16953 28947 17009
rect 29003 16953 29027 16965
rect 29083 16953 29107 16965
rect 29163 16953 29203 17009
rect 28903 16931 29203 16953
rect 35225 16112 52392 16181
rect 35225 15868 35382 16112
rect 35690 15868 35789 16112
rect 36097 15868 36177 16112
rect 36485 15868 36610 16112
rect 36918 15868 37017 16112
rect 37325 15868 37405 16112
rect 37713 15868 37812 16112
rect 38120 15868 38240 16112
rect 38548 15868 38646 16112
rect 38954 15868 39035 16112
rect 39343 15868 39441 16112
rect 39749 15868 39947 16112
rect 40255 15868 40354 16112
rect 40662 15868 40742 16112
rect 41050 15868 41149 16112
rect 41457 15868 41577 16112
rect 41885 15868 41984 16112
rect 42292 15868 42372 16112
rect 42680 15868 42779 16112
rect 43087 15868 43233 16112
rect 43541 15868 43639 16112
rect 43947 15868 44028 16112
rect 44336 15868 44434 16112
rect 44742 15868 44862 16112
rect 45170 15868 45269 16112
rect 45577 15868 45657 16112
rect 45965 15868 46064 16112
rect 46372 15868 46570 16112
rect 46878 15868 46977 16112
rect 47285 15868 47365 16112
rect 47673 15868 47772 16112
rect 48080 15868 48200 16112
rect 48508 15868 48607 16112
rect 48915 15868 48995 16112
rect 49303 15868 49402 16112
rect 49710 15868 49929 16112
rect 50237 15868 50357 16112
rect 50665 15868 50764 16112
rect 51072 15868 51152 16112
rect 51460 15868 51559 16112
rect 51867 15868 51997 16112
rect 52305 15868 52392 16112
rect 35225 15821 52392 15868
rect 35205 15514 53130 15573
rect 35205 15270 35291 15514
rect 35599 15270 35698 15514
rect 36006 15270 36086 15514
rect 36394 15270 36493 15514
rect 36801 15270 36921 15514
rect 37229 15270 37328 15514
rect 37636 15270 37716 15514
rect 38024 15270 38123 15514
rect 38431 15270 38628 15514
rect 38936 15270 39035 15514
rect 39343 15270 39423 15514
rect 39731 15270 39830 15514
rect 40138 15270 40258 15514
rect 40566 15270 40665 15514
rect 40973 15270 41053 15514
rect 41361 15270 41460 15514
rect 41768 15270 41914 15514
rect 42222 15270 42321 15514
rect 42629 15270 42709 15514
rect 43017 15270 43116 15514
rect 43424 15270 43544 15514
rect 43852 15270 43950 15514
rect 44258 15270 44339 15514
rect 44647 15270 44745 15514
rect 45053 15270 45251 15514
rect 45559 15270 45658 15514
rect 45966 15270 46046 15514
rect 46354 15270 46453 15514
rect 46761 15270 46881 15514
rect 47189 15270 47288 15514
rect 47596 15270 47676 15514
rect 47984 15270 48083 15514
rect 48391 15270 48610 15514
rect 48918 15270 49038 15514
rect 49346 15270 49445 15514
rect 49753 15270 49833 15514
rect 50141 15270 50240 15514
rect 50548 15270 53130 15514
rect 35205 15213 53130 15270
rect 41851 -4666 55252 -4644
rect 41851 -4722 42514 -4666
rect 42570 -4722 42594 -4666
rect 42650 -4722 42674 -4666
rect 42730 -4715 55252 -4666
rect 42730 -4722 55033 -4715
rect 41851 -4748 55033 -4722
rect 41851 -4766 54878 -4748
rect 41851 -4822 42514 -4766
rect 42570 -4822 42594 -4766
rect 42650 -4822 42674 -4766
rect 42730 -4822 54878 -4766
rect 41851 -4866 54878 -4822
rect 41851 -4922 42514 -4866
rect 42570 -4922 42594 -4866
rect 42650 -4922 42674 -4866
rect 42730 -4922 54878 -4866
rect 41851 -4928 54878 -4922
rect 54994 -4928 55033 -4748
rect 41851 -4959 55033 -4928
rect 55213 -4959 55252 -4715
rect 41851 -4966 55252 -4959
rect 41851 -5022 42514 -4966
rect 42570 -5022 42594 -4966
rect 42650 -5022 42674 -4966
rect 42730 -5022 55252 -4966
rect 41851 -5044 55252 -5022
rect 49180 -5264 55258 -5193
rect 49180 -5297 55050 -5264
rect 49180 -5477 54895 -5297
rect 55011 -5477 55050 -5297
rect 49180 -5508 55050 -5477
rect 55230 -5508 55258 -5264
rect 49180 -5593 55258 -5508
rect 8750 -5622 28192 -5600
rect 8750 -5678 8794 -5622
rect 8850 -5678 8874 -5622
rect 8930 -5678 8954 -5622
rect 9010 -5678 14166 -5622
rect 14222 -5678 14246 -5622
rect 14302 -5678 14326 -5622
rect 14382 -5678 21181 -5622
rect 21237 -5678 21261 -5622
rect 21317 -5678 21341 -5622
rect 21397 -5678 27936 -5622
rect 27992 -5678 28016 -5622
rect 28072 -5678 28096 -5622
rect 28152 -5678 28192 -5622
rect 8750 -5722 28192 -5678
rect 8750 -5778 8794 -5722
rect 8850 -5778 8874 -5722
rect 8930 -5778 8954 -5722
rect 9010 -5778 14166 -5722
rect 14222 -5778 14246 -5722
rect 14302 -5778 14326 -5722
rect 14382 -5778 21181 -5722
rect 21237 -5778 21261 -5722
rect 21317 -5778 21341 -5722
rect 21397 -5778 27936 -5722
rect 27992 -5778 28016 -5722
rect 28072 -5778 28096 -5722
rect 28152 -5778 28192 -5722
rect 8750 -5822 28192 -5778
rect 8750 -5878 8794 -5822
rect 8850 -5878 8874 -5822
rect 8930 -5878 8954 -5822
rect 9010 -5878 14166 -5822
rect 14222 -5878 14246 -5822
rect 14302 -5878 14326 -5822
rect 14382 -5878 21181 -5822
rect 21237 -5878 21261 -5822
rect 21317 -5878 21341 -5822
rect 21397 -5878 27936 -5822
rect 27992 -5878 28016 -5822
rect 28072 -5878 28096 -5822
rect 28152 -5878 28192 -5822
rect 8750 -5922 28192 -5878
rect 8750 -5978 8794 -5922
rect 8850 -5978 8874 -5922
rect 8930 -5978 8954 -5922
rect 9010 -5978 14166 -5922
rect 14222 -5978 14246 -5922
rect 14302 -5978 14326 -5922
rect 14382 -5978 21181 -5922
rect 21237 -5978 21261 -5922
rect 21317 -5978 21341 -5922
rect 21397 -5978 27936 -5922
rect 27992 -5978 28016 -5922
rect 28072 -5978 28096 -5922
rect 28152 -5978 28192 -5922
rect 8750 -6000 28192 -5978
rect 6977 -6561 20623 -6539
rect 6977 -6617 7021 -6561
rect 7077 -6617 7101 -6561
rect 7157 -6617 7181 -6561
rect 7237 -6617 20363 -6561
rect 20419 -6617 20443 -6561
rect 20499 -6617 20523 -6561
rect 20579 -6617 20623 -6561
rect 6977 -6661 20623 -6617
rect 6977 -6717 7021 -6661
rect 7077 -6717 7101 -6661
rect 7157 -6717 7181 -6661
rect 7237 -6717 20363 -6661
rect 20419 -6717 20443 -6661
rect 20499 -6717 20523 -6661
rect 20579 -6717 20623 -6661
rect 6977 -6761 20623 -6717
rect 6977 -6817 7021 -6761
rect 7077 -6817 7101 -6761
rect 7157 -6817 7181 -6761
rect 7237 -6817 20363 -6761
rect 20419 -6817 20443 -6761
rect 20499 -6817 20523 -6761
rect 20579 -6817 20623 -6761
rect 6977 -6861 20623 -6817
rect 6977 -6917 7021 -6861
rect 7077 -6917 7101 -6861
rect 7157 -6917 7181 -6861
rect 7237 -6917 20363 -6861
rect 20419 -6917 20443 -6861
rect 20499 -6917 20523 -6861
rect 20579 -6917 20623 -6861
rect 6977 -6939 20623 -6917
rect 22917 -7688 30059 -7666
rect 22917 -7744 22961 -7688
rect 23017 -7744 23041 -7688
rect 23097 -7744 23121 -7688
rect 23177 -7744 29803 -7688
rect 29859 -7744 29883 -7688
rect 29939 -7744 29963 -7688
rect 30019 -7744 30059 -7688
rect 22917 -7788 30059 -7744
rect 22917 -7844 22961 -7788
rect 23017 -7844 23041 -7788
rect 23097 -7844 23121 -7788
rect 23177 -7844 29803 -7788
rect 29859 -7844 29883 -7788
rect 29939 -7844 29963 -7788
rect 30019 -7844 30059 -7788
rect 22917 -7888 30059 -7844
rect 22917 -7944 22961 -7888
rect 23017 -7944 23041 -7888
rect 23097 -7944 23121 -7888
rect 23177 -7944 29803 -7888
rect 29859 -7944 29883 -7888
rect 29939 -7944 29963 -7888
rect 30019 -7944 30059 -7888
rect 22917 -7988 30059 -7944
rect 22917 -8044 22961 -7988
rect 23017 -8044 23041 -7988
rect 23097 -8044 23121 -7988
rect 23177 -8044 29803 -7988
rect 29859 -8044 29883 -7988
rect 29939 -8044 29963 -7988
rect 30019 -8044 30059 -7988
rect 22917 -8066 30059 -8044
rect 29034 -8424 33079 -8385
rect 29034 -8480 29078 -8424
rect 29134 -8480 29158 -8424
rect 29214 -8480 29238 -8424
rect 29294 -8480 33079 -8424
rect 29034 -8524 33079 -8480
rect 29034 -8580 29078 -8524
rect 29134 -8580 29158 -8524
rect 29214 -8580 29238 -8524
rect 29294 -8580 33079 -8524
rect 29034 -8624 33079 -8580
rect 29034 -8680 29078 -8624
rect 29134 -8680 29158 -8624
rect 29214 -8680 29238 -8624
rect 29294 -8680 33079 -8624
rect 29034 -8724 33079 -8680
rect 29034 -8780 29078 -8724
rect 29134 -8780 29158 -8724
rect 29214 -8780 29238 -8724
rect 29294 -8780 33079 -8724
rect 29034 -8802 33079 -8780
rect 37669 -8424 41296 -8385
rect 37669 -8480 41036 -8424
rect 41092 -8480 41116 -8424
rect 41172 -8480 41196 -8424
rect 41252 -8480 41296 -8424
rect 37669 -8524 41296 -8480
rect 37669 -8580 41036 -8524
rect 41092 -8580 41116 -8524
rect 41172 -8580 41196 -8524
rect 41252 -8580 41296 -8524
rect 37669 -8624 41296 -8580
rect 37669 -8680 41036 -8624
rect 41092 -8680 41116 -8624
rect 41172 -8680 41196 -8624
rect 41252 -8680 41296 -8624
rect 37669 -8724 41296 -8680
rect 37669 -8780 41036 -8724
rect 41092 -8780 41116 -8724
rect 41172 -8780 41196 -8724
rect 41252 -8780 41296 -8724
rect 37669 -8802 41296 -8780
rect 22917 -10062 30059 -10040
rect 22917 -10118 22961 -10062
rect 23017 -10118 23041 -10062
rect 23097 -10118 23121 -10062
rect 23177 -10118 29803 -10062
rect 29859 -10118 29883 -10062
rect 29939 -10118 29963 -10062
rect 30019 -10118 30059 -10062
rect 22917 -10162 30059 -10118
rect 22917 -10218 22961 -10162
rect 23017 -10218 23041 -10162
rect 23097 -10218 23121 -10162
rect 23177 -10218 29803 -10162
rect 29859 -10218 29883 -10162
rect 29939 -10218 29963 -10162
rect 30019 -10218 30059 -10162
rect 22917 -10262 30059 -10218
rect 22917 -10318 22961 -10262
rect 23017 -10318 23041 -10262
rect 23097 -10318 23121 -10262
rect 23177 -10318 29803 -10262
rect 29859 -10318 29883 -10262
rect 29939 -10318 29963 -10262
rect 30019 -10318 30059 -10262
rect 22917 -10362 30059 -10318
rect 22917 -10418 22961 -10362
rect 23017 -10418 23041 -10362
rect 23097 -10418 23121 -10362
rect 23177 -10418 29803 -10362
rect 29859 -10418 29883 -10362
rect 29939 -10418 29963 -10362
rect 30019 -10418 30059 -10362
rect 22917 -10440 30059 -10418
rect 25575 -14270 51603 -14248
rect 25575 -14326 31057 -14270
rect 31113 -14326 31137 -14270
rect 31193 -14326 31217 -14270
rect 31273 -14326 39447 -14270
rect 39503 -14326 39527 -14270
rect 39583 -14326 39607 -14270
rect 39663 -14326 42957 -14270
rect 43013 -14326 43037 -14270
rect 43093 -14326 43117 -14270
rect 43173 -14326 51347 -14270
rect 51403 -14326 51427 -14270
rect 51483 -14326 51507 -14270
rect 51563 -14326 51603 -14270
rect 25575 -14370 51603 -14326
rect 25575 -14426 31057 -14370
rect 31113 -14426 31137 -14370
rect 31193 -14426 31217 -14370
rect 31273 -14426 39447 -14370
rect 39503 -14426 39527 -14370
rect 39583 -14426 39607 -14370
rect 39663 -14426 42957 -14370
rect 43013 -14426 43037 -14370
rect 43093 -14426 43117 -14370
rect 43173 -14426 51347 -14370
rect 51403 -14426 51427 -14370
rect 51483 -14426 51507 -14370
rect 51563 -14426 51603 -14370
rect 25575 -14470 51603 -14426
rect 25575 -14526 31057 -14470
rect 31113 -14526 31137 -14470
rect 31193 -14526 31217 -14470
rect 31273 -14526 39447 -14470
rect 39503 -14526 39527 -14470
rect 39583 -14526 39607 -14470
rect 39663 -14526 42957 -14470
rect 43013 -14526 43037 -14470
rect 43093 -14526 43117 -14470
rect 43173 -14526 51347 -14470
rect 51403 -14526 51427 -14470
rect 51483 -14526 51507 -14470
rect 51563 -14526 51603 -14470
rect 25575 -14570 51603 -14526
rect 25575 -14626 31057 -14570
rect 31113 -14626 31137 -14570
rect 31193 -14626 31217 -14570
rect 31273 -14626 39447 -14570
rect 39503 -14626 39527 -14570
rect 39583 -14626 39607 -14570
rect 39663 -14626 42957 -14570
rect 43013 -14626 43037 -14570
rect 43093 -14626 43117 -14570
rect 43173 -14626 51347 -14570
rect 51403 -14626 51427 -14570
rect 51483 -14626 51507 -14570
rect 51563 -14626 51603 -14570
rect 25575 -14648 51603 -14626
rect 25575 -14683 26336 -14648
rect 22026 -14705 26336 -14683
rect 22026 -14761 22070 -14705
rect 22126 -14761 22150 -14705
rect 22206 -14761 22230 -14705
rect 22286 -14761 26336 -14705
rect 22026 -14805 26336 -14761
rect 22026 -14861 22070 -14805
rect 22126 -14861 22150 -14805
rect 22206 -14861 22230 -14805
rect 22286 -14861 26336 -14805
rect 22026 -14905 26336 -14861
rect 22026 -14961 22070 -14905
rect 22126 -14961 22150 -14905
rect 22206 -14961 22230 -14905
rect 22286 -14961 26336 -14905
rect 22026 -15005 26336 -14961
rect 22026 -15061 22070 -15005
rect 22126 -15061 22150 -15005
rect 22206 -15061 22230 -15005
rect 22286 -15061 26336 -15005
rect 22026 -15083 26336 -15061
rect 29759 -14982 40562 -14960
rect 29759 -15038 29803 -14982
rect 29859 -15038 29883 -14982
rect 29939 -15038 29963 -14982
rect 30019 -15038 40306 -14982
rect 40362 -15038 40386 -14982
rect 40442 -15038 40466 -14982
rect 40522 -15038 40562 -14982
rect 29759 -15082 40562 -15038
rect 29759 -15138 29803 -15082
rect 29859 -15138 29883 -15082
rect 29939 -15138 29963 -15082
rect 30019 -15138 40306 -15082
rect 40362 -15138 40386 -15082
rect 40442 -15138 40466 -15082
rect 40522 -15138 40562 -15082
rect 29759 -15182 40562 -15138
rect 29759 -15238 29803 -15182
rect 29859 -15238 29883 -15182
rect 29939 -15238 29963 -15182
rect 30019 -15238 40306 -15182
rect 40362 -15238 40386 -15182
rect 40442 -15238 40466 -15182
rect 40522 -15238 40562 -15182
rect 29759 -15282 40562 -15238
rect 29759 -15338 29803 -15282
rect 29859 -15338 29883 -15282
rect 29939 -15338 29963 -15282
rect 30019 -15338 40306 -15282
rect 40362 -15338 40386 -15282
rect 40442 -15338 40466 -15282
rect 40522 -15338 40562 -15282
rect 29759 -15360 40562 -15338
rect 41986 -14982 53365 -14960
rect 41986 -15038 42030 -14982
rect 42086 -15038 42110 -14982
rect 42166 -15038 42190 -14982
rect 42246 -15038 52360 -14982
rect 52416 -15038 52440 -14982
rect 52496 -15038 52520 -14982
rect 52576 -15033 53365 -14982
rect 52576 -15038 53116 -15033
rect 41986 -15066 53116 -15038
rect 41986 -15082 52961 -15066
rect 41986 -15138 42030 -15082
rect 42086 -15138 42110 -15082
rect 42166 -15138 42190 -15082
rect 42246 -15138 52360 -15082
rect 52416 -15138 52440 -15082
rect 52496 -15138 52520 -15082
rect 52576 -15138 52961 -15082
rect 41986 -15182 52961 -15138
rect 41986 -15238 42030 -15182
rect 42086 -15238 42110 -15182
rect 42166 -15238 42190 -15182
rect 42246 -15238 52360 -15182
rect 52416 -15238 52440 -15182
rect 52496 -15238 52520 -15182
rect 52576 -15238 52961 -15182
rect 41986 -15246 52961 -15238
rect 53077 -15246 53116 -15066
rect 41986 -15277 53116 -15246
rect 53296 -15277 53365 -15033
rect 41986 -15282 53365 -15277
rect 41986 -15338 42030 -15282
rect 42086 -15338 42110 -15282
rect 42166 -15338 42190 -15282
rect 42246 -15338 52360 -15282
rect 52416 -15338 52440 -15282
rect 52496 -15338 52520 -15282
rect 52576 -15338 53365 -15282
rect 41986 -15360 53365 -15338
rect 23076 -15700 41296 -15678
rect 23076 -15756 24906 -15700
rect 24962 -15756 24986 -15700
rect 25042 -15756 25066 -15700
rect 25122 -15756 29078 -15700
rect 29134 -15756 29158 -15700
rect 29214 -15756 29238 -15700
rect 29294 -15756 41040 -15700
rect 41096 -15756 41120 -15700
rect 41176 -15756 41200 -15700
rect 41256 -15756 41296 -15700
rect 23076 -15800 41296 -15756
rect 18543 -15856 18843 -15842
rect 16577 -15864 18843 -15856
rect 16577 -15920 18587 -15864
rect 18643 -15920 18667 -15864
rect 18723 -15920 18747 -15864
rect 18803 -15920 18843 -15864
rect 16577 -15926 18843 -15920
rect 18543 -15942 18843 -15926
rect 23076 -15856 24906 -15800
rect 24962 -15856 24986 -15800
rect 25042 -15856 25066 -15800
rect 25122 -15856 29078 -15800
rect 29134 -15856 29158 -15800
rect 29214 -15856 29238 -15800
rect 29294 -15856 41040 -15800
rect 41096 -15856 41120 -15800
rect 41176 -15856 41200 -15800
rect 41256 -15856 41296 -15800
rect 23076 -15900 41296 -15856
rect 23076 -15956 24906 -15900
rect 24962 -15956 24986 -15900
rect 25042 -15956 25066 -15900
rect 25122 -15956 29078 -15900
rect 29134 -15956 29158 -15900
rect 29214 -15956 29238 -15900
rect 29294 -15956 41040 -15900
rect 41096 -15956 41120 -15900
rect 41176 -15956 41200 -15900
rect 41256 -15956 41296 -15900
rect 23076 -16000 41296 -15956
rect 23076 -16056 24906 -16000
rect 24962 -16056 24986 -16000
rect 25042 -16056 25066 -16000
rect 25122 -16056 29078 -16000
rect 29134 -16056 29158 -16000
rect 29214 -16056 29238 -16000
rect 29294 -16056 41040 -16000
rect 41096 -16056 41120 -16000
rect 41176 -16056 41200 -16000
rect 41256 -16056 41296 -16000
rect 23076 -16078 41296 -16056
rect 16577 -16300 18843 -16275
rect 16577 -16345 18583 -16300
rect 18543 -16356 18583 -16345
rect 18639 -16356 18663 -16300
rect 18719 -16356 18743 -16300
rect 18799 -16356 18843 -16300
rect 18543 -16378 18843 -16356
rect 18542 -17275 25162 -17253
rect 18542 -17331 18583 -17275
rect 18639 -17331 18663 -17275
rect 18719 -17331 18743 -17275
rect 18799 -17331 24902 -17275
rect 24958 -17331 24982 -17275
rect 25038 -17331 25062 -17275
rect 25118 -17331 25162 -17275
rect 18542 -17360 25162 -17331
rect 16577 -17375 25162 -17360
rect 16577 -17430 18583 -17375
rect 18542 -17431 18583 -17430
rect 18639 -17431 18663 -17375
rect 18719 -17431 18743 -17375
rect 18799 -17431 24902 -17375
rect 24958 -17431 24982 -17375
rect 25038 -17431 25062 -17375
rect 25118 -17431 25162 -17375
rect 18542 -17475 25162 -17431
rect 18542 -17531 18583 -17475
rect 18639 -17531 18663 -17475
rect 18719 -17531 18743 -17475
rect 18799 -17531 24902 -17475
rect 24958 -17531 24982 -17475
rect 25038 -17531 25062 -17475
rect 25118 -17531 25162 -17475
rect 18542 -17553 25162 -17531
<< via2 >>
rect 7021 17153 7077 17209
rect 7101 17153 7157 17209
rect 7181 17153 7237 17209
rect 7021 17081 7077 17109
rect 7101 17081 7157 17109
rect 7181 17081 7237 17109
rect 7021 17053 7038 17081
rect 7038 17053 7077 17081
rect 7101 17053 7157 17081
rect 7181 17053 7218 17081
rect 7218 17053 7237 17081
rect 7021 16965 7038 17009
rect 7038 16965 7077 17009
rect 7101 16965 7157 17009
rect 7181 16965 7218 17009
rect 7218 16965 7237 17009
rect 7021 16953 7077 16965
rect 7101 16953 7157 16965
rect 7181 16953 7237 16965
rect 7521 17153 7577 17209
rect 7601 17153 7657 17209
rect 7681 17153 7737 17209
rect 7521 17081 7577 17109
rect 7601 17081 7657 17109
rect 7681 17081 7737 17109
rect 7521 17053 7535 17081
rect 7535 17053 7577 17081
rect 7601 17053 7657 17081
rect 7681 17053 7715 17081
rect 7715 17053 7737 17081
rect 7521 16965 7535 17009
rect 7535 16965 7577 17009
rect 7601 16965 7657 17009
rect 7681 16965 7715 17009
rect 7715 16965 7737 17009
rect 7521 16953 7577 16965
rect 7601 16953 7657 16965
rect 7681 16953 7737 16965
rect 8020 17153 8076 17209
rect 8100 17153 8156 17209
rect 8180 17153 8236 17209
rect 8020 17081 8076 17109
rect 8100 17081 8156 17109
rect 8180 17081 8236 17109
rect 8020 17053 8033 17081
rect 8033 17053 8076 17081
rect 8100 17053 8156 17081
rect 8180 17053 8213 17081
rect 8213 17053 8236 17081
rect 8020 16965 8033 17009
rect 8033 16965 8076 17009
rect 8100 16965 8156 17009
rect 8180 16965 8213 17009
rect 8213 16965 8236 17009
rect 8020 16953 8076 16965
rect 8100 16953 8156 16965
rect 8180 16953 8236 16965
rect 28448 17153 28504 17209
rect 28528 17153 28584 17209
rect 28608 17153 28664 17209
rect 28448 17081 28504 17109
rect 28528 17081 28584 17109
rect 28608 17081 28664 17109
rect 28448 17053 28462 17081
rect 28462 17053 28504 17081
rect 28528 17053 28584 17081
rect 28608 17053 28642 17081
rect 28642 17053 28664 17081
rect 28448 16965 28462 17009
rect 28462 16965 28504 17009
rect 28528 16965 28584 17009
rect 28608 16965 28642 17009
rect 28642 16965 28664 17009
rect 28448 16953 28504 16965
rect 28528 16953 28584 16965
rect 28608 16953 28664 16965
rect 28947 17153 29003 17209
rect 29027 17153 29083 17209
rect 29107 17153 29163 17209
rect 28947 17081 29003 17109
rect 29027 17081 29083 17109
rect 29107 17081 29163 17109
rect 28947 17053 28960 17081
rect 28960 17053 29003 17081
rect 29027 17053 29083 17081
rect 29107 17053 29140 17081
rect 29140 17053 29163 17081
rect 28947 16965 28960 17009
rect 28960 16965 29003 17009
rect 29027 16965 29083 17009
rect 29107 16965 29140 17009
rect 29140 16965 29163 17009
rect 28947 16953 29003 16965
rect 29027 16953 29083 16965
rect 29107 16953 29163 16965
rect 42514 -4722 42570 -4666
rect 42594 -4722 42650 -4666
rect 42674 -4722 42730 -4666
rect 42514 -4822 42570 -4766
rect 42594 -4822 42650 -4766
rect 42674 -4822 42730 -4766
rect 42514 -4922 42570 -4866
rect 42594 -4922 42650 -4866
rect 42674 -4922 42730 -4866
rect 42514 -5022 42570 -4966
rect 42594 -5022 42650 -4966
rect 42674 -5022 42730 -4966
rect 8794 -5678 8850 -5622
rect 8874 -5678 8930 -5622
rect 8954 -5678 9010 -5622
rect 14166 -5678 14222 -5622
rect 14246 -5678 14302 -5622
rect 14326 -5678 14382 -5622
rect 21181 -5678 21237 -5622
rect 21261 -5678 21317 -5622
rect 21341 -5678 21397 -5622
rect 27936 -5678 27992 -5622
rect 28016 -5678 28072 -5622
rect 28096 -5678 28152 -5622
rect 8794 -5778 8850 -5722
rect 8874 -5778 8930 -5722
rect 8954 -5778 9010 -5722
rect 14166 -5778 14222 -5722
rect 14246 -5778 14302 -5722
rect 14326 -5778 14382 -5722
rect 21181 -5778 21237 -5722
rect 21261 -5778 21317 -5722
rect 21341 -5778 21397 -5722
rect 27936 -5778 27992 -5722
rect 28016 -5778 28072 -5722
rect 28096 -5778 28152 -5722
rect 8794 -5878 8850 -5822
rect 8874 -5878 8930 -5822
rect 8954 -5878 9010 -5822
rect 14166 -5878 14222 -5822
rect 14246 -5878 14302 -5822
rect 14326 -5878 14382 -5822
rect 21181 -5878 21237 -5822
rect 21261 -5878 21317 -5822
rect 21341 -5878 21397 -5822
rect 27936 -5878 27992 -5822
rect 28016 -5878 28072 -5822
rect 28096 -5878 28152 -5822
rect 8794 -5978 8850 -5922
rect 8874 -5978 8930 -5922
rect 8954 -5978 9010 -5922
rect 14166 -5978 14222 -5922
rect 14246 -5978 14302 -5922
rect 14326 -5978 14382 -5922
rect 21181 -5978 21237 -5922
rect 21261 -5978 21317 -5922
rect 21341 -5978 21397 -5922
rect 27936 -5978 27992 -5922
rect 28016 -5978 28072 -5922
rect 28096 -5978 28152 -5922
rect 7021 -6617 7077 -6561
rect 7101 -6617 7157 -6561
rect 7181 -6617 7237 -6561
rect 20363 -6617 20419 -6561
rect 20443 -6617 20499 -6561
rect 20523 -6617 20579 -6561
rect 7021 -6717 7077 -6661
rect 7101 -6717 7157 -6661
rect 7181 -6717 7237 -6661
rect 20363 -6717 20419 -6661
rect 20443 -6717 20499 -6661
rect 20523 -6717 20579 -6661
rect 7021 -6817 7077 -6761
rect 7101 -6817 7157 -6761
rect 7181 -6817 7237 -6761
rect 20363 -6817 20419 -6761
rect 20443 -6817 20499 -6761
rect 20523 -6817 20579 -6761
rect 7021 -6917 7077 -6861
rect 7101 -6917 7157 -6861
rect 7181 -6917 7237 -6861
rect 20363 -6917 20419 -6861
rect 20443 -6917 20499 -6861
rect 20523 -6917 20579 -6861
rect 22961 -7744 23017 -7688
rect 23041 -7744 23097 -7688
rect 23121 -7744 23177 -7688
rect 29803 -7744 29859 -7688
rect 29883 -7744 29939 -7688
rect 29963 -7744 30019 -7688
rect 22961 -7844 23017 -7788
rect 23041 -7844 23097 -7788
rect 23121 -7844 23177 -7788
rect 29803 -7844 29859 -7788
rect 29883 -7844 29939 -7788
rect 29963 -7844 30019 -7788
rect 22961 -7944 23017 -7888
rect 23041 -7944 23097 -7888
rect 23121 -7944 23177 -7888
rect 29803 -7944 29859 -7888
rect 29883 -7944 29939 -7888
rect 29963 -7944 30019 -7888
rect 22961 -8044 23017 -7988
rect 23041 -8044 23097 -7988
rect 23121 -8044 23177 -7988
rect 29803 -8044 29859 -7988
rect 29883 -8044 29939 -7988
rect 29963 -8044 30019 -7988
rect 29078 -8480 29134 -8424
rect 29158 -8480 29214 -8424
rect 29238 -8480 29294 -8424
rect 29078 -8580 29134 -8524
rect 29158 -8580 29214 -8524
rect 29238 -8580 29294 -8524
rect 29078 -8680 29134 -8624
rect 29158 -8680 29214 -8624
rect 29238 -8680 29294 -8624
rect 29078 -8780 29134 -8724
rect 29158 -8780 29214 -8724
rect 29238 -8780 29294 -8724
rect 41036 -8480 41092 -8424
rect 41116 -8480 41172 -8424
rect 41196 -8480 41252 -8424
rect 41036 -8580 41092 -8524
rect 41116 -8580 41172 -8524
rect 41196 -8580 41252 -8524
rect 41036 -8680 41092 -8624
rect 41116 -8680 41172 -8624
rect 41196 -8680 41252 -8624
rect 41036 -8780 41092 -8724
rect 41116 -8780 41172 -8724
rect 41196 -8780 41252 -8724
rect 22961 -10118 23017 -10062
rect 23041 -10118 23097 -10062
rect 23121 -10118 23177 -10062
rect 29803 -10118 29859 -10062
rect 29883 -10118 29939 -10062
rect 29963 -10118 30019 -10062
rect 22961 -10218 23017 -10162
rect 23041 -10218 23097 -10162
rect 23121 -10218 23177 -10162
rect 29803 -10218 29859 -10162
rect 29883 -10218 29939 -10162
rect 29963 -10218 30019 -10162
rect 22961 -10318 23017 -10262
rect 23041 -10318 23097 -10262
rect 23121 -10318 23177 -10262
rect 29803 -10318 29859 -10262
rect 29883 -10318 29939 -10262
rect 29963 -10318 30019 -10262
rect 22961 -10418 23017 -10362
rect 23041 -10418 23097 -10362
rect 23121 -10418 23177 -10362
rect 29803 -10418 29859 -10362
rect 29883 -10418 29939 -10362
rect 29963 -10418 30019 -10362
rect 31057 -14326 31113 -14270
rect 31137 -14326 31193 -14270
rect 31217 -14326 31273 -14270
rect 39447 -14326 39503 -14270
rect 39527 -14326 39583 -14270
rect 39607 -14326 39663 -14270
rect 42957 -14326 43013 -14270
rect 43037 -14326 43093 -14270
rect 43117 -14326 43173 -14270
rect 51347 -14326 51403 -14270
rect 51427 -14326 51483 -14270
rect 51507 -14326 51563 -14270
rect 31057 -14426 31113 -14370
rect 31137 -14426 31193 -14370
rect 31217 -14426 31273 -14370
rect 39447 -14426 39503 -14370
rect 39527 -14426 39583 -14370
rect 39607 -14426 39663 -14370
rect 42957 -14426 43013 -14370
rect 43037 -14426 43093 -14370
rect 43117 -14426 43173 -14370
rect 51347 -14426 51403 -14370
rect 51427 -14426 51483 -14370
rect 51507 -14426 51563 -14370
rect 31057 -14526 31113 -14470
rect 31137 -14526 31193 -14470
rect 31217 -14526 31273 -14470
rect 39447 -14526 39503 -14470
rect 39527 -14526 39583 -14470
rect 39607 -14526 39663 -14470
rect 42957 -14526 43013 -14470
rect 43037 -14526 43093 -14470
rect 43117 -14526 43173 -14470
rect 51347 -14526 51403 -14470
rect 51427 -14526 51483 -14470
rect 51507 -14526 51563 -14470
rect 31057 -14626 31113 -14570
rect 31137 -14626 31193 -14570
rect 31217 -14626 31273 -14570
rect 39447 -14626 39503 -14570
rect 39527 -14626 39583 -14570
rect 39607 -14626 39663 -14570
rect 42957 -14626 43013 -14570
rect 43037 -14626 43093 -14570
rect 43117 -14626 43173 -14570
rect 51347 -14626 51403 -14570
rect 51427 -14626 51483 -14570
rect 51507 -14626 51563 -14570
rect 22070 -14761 22126 -14705
rect 22150 -14761 22206 -14705
rect 22230 -14761 22286 -14705
rect 22070 -14861 22126 -14805
rect 22150 -14861 22206 -14805
rect 22230 -14861 22286 -14805
rect 22070 -14961 22126 -14905
rect 22150 -14961 22206 -14905
rect 22230 -14961 22286 -14905
rect 22070 -15061 22126 -15005
rect 22150 -15061 22206 -15005
rect 22230 -15061 22286 -15005
rect 29803 -15038 29859 -14982
rect 29883 -15038 29939 -14982
rect 29963 -15038 30019 -14982
rect 40306 -15038 40362 -14982
rect 40386 -15038 40442 -14982
rect 40466 -15038 40522 -14982
rect 29803 -15138 29859 -15082
rect 29883 -15138 29939 -15082
rect 29963 -15138 30019 -15082
rect 40306 -15138 40362 -15082
rect 40386 -15138 40442 -15082
rect 40466 -15138 40522 -15082
rect 29803 -15238 29859 -15182
rect 29883 -15238 29939 -15182
rect 29963 -15238 30019 -15182
rect 40306 -15238 40362 -15182
rect 40386 -15238 40442 -15182
rect 40466 -15238 40522 -15182
rect 29803 -15338 29859 -15282
rect 29883 -15338 29939 -15282
rect 29963 -15338 30019 -15282
rect 40306 -15338 40362 -15282
rect 40386 -15338 40442 -15282
rect 40466 -15338 40522 -15282
rect 42030 -15038 42086 -14982
rect 42110 -15038 42166 -14982
rect 42190 -15038 42246 -14982
rect 52360 -15038 52416 -14982
rect 52440 -15038 52496 -14982
rect 52520 -15038 52576 -14982
rect 42030 -15138 42086 -15082
rect 42110 -15138 42166 -15082
rect 42190 -15138 42246 -15082
rect 52360 -15138 52416 -15082
rect 52440 -15138 52496 -15082
rect 52520 -15138 52576 -15082
rect 42030 -15238 42086 -15182
rect 42110 -15238 42166 -15182
rect 42190 -15238 42246 -15182
rect 52360 -15238 52416 -15182
rect 52440 -15238 52496 -15182
rect 52520 -15238 52576 -15182
rect 42030 -15338 42086 -15282
rect 42110 -15338 42166 -15282
rect 42190 -15338 42246 -15282
rect 52360 -15338 52416 -15282
rect 52440 -15338 52496 -15282
rect 52520 -15338 52576 -15282
rect 24906 -15756 24962 -15700
rect 24986 -15756 25042 -15700
rect 25066 -15756 25122 -15700
rect 29078 -15756 29134 -15700
rect 29158 -15756 29214 -15700
rect 29238 -15756 29294 -15700
rect 41040 -15756 41096 -15700
rect 41120 -15756 41176 -15700
rect 41200 -15756 41256 -15700
rect 18587 -15920 18643 -15864
rect 18667 -15920 18723 -15864
rect 18747 -15920 18803 -15864
rect 24906 -15856 24962 -15800
rect 24986 -15856 25042 -15800
rect 25066 -15856 25122 -15800
rect 29078 -15856 29134 -15800
rect 29158 -15856 29214 -15800
rect 29238 -15856 29294 -15800
rect 41040 -15856 41096 -15800
rect 41120 -15856 41176 -15800
rect 41200 -15856 41256 -15800
rect 24906 -15956 24962 -15900
rect 24986 -15956 25042 -15900
rect 25066 -15956 25122 -15900
rect 29078 -15956 29134 -15900
rect 29158 -15956 29214 -15900
rect 29238 -15956 29294 -15900
rect 41040 -15956 41096 -15900
rect 41120 -15956 41176 -15900
rect 41200 -15956 41256 -15900
rect 24906 -16056 24962 -16000
rect 24986 -16056 25042 -16000
rect 25066 -16056 25122 -16000
rect 29078 -16056 29134 -16000
rect 29158 -16056 29214 -16000
rect 29238 -16056 29294 -16000
rect 41040 -16056 41096 -16000
rect 41120 -16056 41176 -16000
rect 41200 -16056 41256 -16000
rect 18583 -16356 18639 -16300
rect 18663 -16356 18719 -16300
rect 18743 -16356 18799 -16300
rect 18583 -17331 18639 -17275
rect 18663 -17331 18719 -17275
rect 18743 -17331 18799 -17275
rect 24902 -17331 24958 -17275
rect 24982 -17331 25038 -17275
rect 25062 -17331 25118 -17275
rect 18583 -17431 18639 -17375
rect 18663 -17431 18719 -17375
rect 18743 -17431 18799 -17375
rect 24902 -17431 24958 -17375
rect 24982 -17431 25038 -17375
rect 25062 -17431 25118 -17375
rect 18583 -17531 18639 -17475
rect 18663 -17531 18719 -17475
rect 18743 -17531 18799 -17475
rect 24902 -17531 24958 -17475
rect 24982 -17531 25038 -17475
rect 25062 -17531 25118 -17475
<< metal3 >>
rect 6977 17209 7277 17295
rect 6977 17153 7021 17209
rect 7077 17153 7101 17209
rect 7157 17153 7181 17209
rect 7237 17153 7277 17209
rect 6977 17109 7277 17153
rect 6977 17053 7021 17109
rect 7077 17053 7101 17109
rect 7157 17053 7181 17109
rect 7237 17053 7277 17109
rect 6977 17009 7277 17053
rect 6977 16953 7021 17009
rect 7077 16953 7101 17009
rect 7157 16953 7181 17009
rect 7237 16953 7277 17009
rect 6977 -6561 7277 16953
rect 7477 17209 7777 17295
rect 7477 17153 7521 17209
rect 7577 17153 7601 17209
rect 7657 17153 7681 17209
rect 7737 17153 7777 17209
rect 7477 17109 7777 17153
rect 7477 17053 7521 17109
rect 7577 17053 7601 17109
rect 7657 17053 7681 17109
rect 7737 17053 7777 17109
rect 7477 17009 7777 17053
rect 7477 16953 7521 17009
rect 7577 16953 7601 17009
rect 7657 16953 7681 17009
rect 7737 16953 7777 17009
rect 7477 -1436 7777 16953
rect 7976 17209 8276 17295
rect 7976 17153 8020 17209
rect 8076 17153 8100 17209
rect 8156 17153 8180 17209
rect 8236 17153 8276 17209
rect 7976 17109 8276 17153
rect 7976 17053 8020 17109
rect 8076 17053 8100 17109
rect 8156 17053 8180 17109
rect 8236 17053 8276 17109
rect 7976 17009 8276 17053
rect 7976 16953 8020 17009
rect 8076 16953 8100 17009
rect 8156 16953 8180 17009
rect 8236 16953 8276 17009
rect 7976 -1436 8276 16953
rect 28404 17209 28704 17231
rect 28404 17153 28448 17209
rect 28504 17153 28528 17209
rect 28584 17153 28608 17209
rect 28664 17153 28704 17209
rect 28404 17109 28704 17153
rect 28404 17053 28448 17109
rect 28504 17053 28528 17109
rect 28584 17053 28608 17109
rect 28664 17053 28704 17109
rect 28404 17009 28704 17053
rect 28404 16953 28448 17009
rect 28504 16953 28528 17009
rect 28584 16953 28608 17009
rect 28664 16953 28704 17009
rect 8750 -5622 9050 11594
rect 8750 -5678 8794 -5622
rect 8850 -5678 8874 -5622
rect 8930 -5678 8954 -5622
rect 9010 -5678 9050 -5622
rect 8750 -5722 9050 -5678
rect 8750 -5778 8794 -5722
rect 8850 -5778 8874 -5722
rect 8930 -5778 8954 -5722
rect 9010 -5778 9050 -5722
rect 8750 -5822 9050 -5778
rect 8750 -5878 8794 -5822
rect 8850 -5878 8874 -5822
rect 8930 -5878 8954 -5822
rect 9010 -5878 9050 -5822
rect 8750 -5922 9050 -5878
rect 8750 -5978 8794 -5922
rect 8850 -5978 8874 -5922
rect 8930 -5978 8954 -5922
rect 9010 -5978 9050 -5922
rect 8750 -6000 9050 -5978
rect 14126 -5622 14426 -5600
rect 14126 -5678 14166 -5622
rect 14222 -5678 14246 -5622
rect 14302 -5678 14326 -5622
rect 14382 -5678 14426 -5622
rect 14126 -5722 14426 -5678
rect 14126 -5778 14166 -5722
rect 14222 -5778 14246 -5722
rect 14302 -5778 14326 -5722
rect 14382 -5778 14426 -5722
rect 14126 -5822 14426 -5778
rect 14126 -5878 14166 -5822
rect 14222 -5878 14246 -5822
rect 14302 -5878 14326 -5822
rect 14382 -5878 14426 -5822
rect 14126 -5922 14426 -5878
rect 14126 -5978 14166 -5922
rect 14222 -5978 14246 -5922
rect 14302 -5978 14326 -5922
rect 14382 -5978 14426 -5922
rect 6977 -6617 7021 -6561
rect 7077 -6617 7101 -6561
rect 7157 -6617 7181 -6561
rect 7237 -6617 7277 -6561
rect 6977 -6661 7277 -6617
rect 6977 -6717 7021 -6661
rect 7077 -6717 7101 -6661
rect 7157 -6717 7181 -6661
rect 7237 -6717 7277 -6661
rect 6977 -6761 7277 -6717
rect 6977 -6817 7021 -6761
rect 7077 -6817 7101 -6761
rect 7157 -6817 7181 -6761
rect 7237 -6817 7277 -6761
rect 6977 -6861 7277 -6817
rect 6977 -6917 7021 -6861
rect 7077 -6917 7101 -6861
rect 7157 -6917 7181 -6861
rect 7237 -6917 7277 -6861
rect 6977 -6939 7277 -6917
rect 14126 -8285 14426 -5978
rect 21141 -5622 21442 -5600
rect 21141 -5678 21181 -5622
rect 21237 -5678 21261 -5622
rect 21317 -5678 21341 -5622
rect 21397 -5678 21442 -5622
rect 21141 -5722 21442 -5678
rect 21141 -5778 21181 -5722
rect 21237 -5778 21261 -5722
rect 21317 -5778 21341 -5722
rect 21397 -5778 21442 -5722
rect 21141 -5822 21442 -5778
rect 21141 -5878 21181 -5822
rect 21237 -5878 21261 -5822
rect 21317 -5878 21341 -5822
rect 21397 -5878 21442 -5822
rect 21141 -5922 21442 -5878
rect 21141 -5978 21181 -5922
rect 21237 -5978 21261 -5922
rect 21317 -5978 21341 -5922
rect 21397 -5978 21442 -5922
rect 20323 -6561 20623 -6539
rect 20323 -6617 20363 -6561
rect 20419 -6617 20443 -6561
rect 20499 -6617 20523 -6561
rect 20579 -6617 20623 -6561
rect 20323 -6661 20623 -6617
rect 20323 -6717 20363 -6661
rect 20419 -6717 20443 -6661
rect 20499 -6717 20523 -6661
rect 20579 -6717 20623 -6661
rect 20323 -6761 20623 -6717
rect 20323 -6817 20363 -6761
rect 20419 -6817 20443 -6761
rect 20499 -6817 20523 -6761
rect 20579 -6817 20623 -6761
rect 20323 -6861 20623 -6817
rect 20323 -6917 20363 -6861
rect 20419 -6917 20443 -6861
rect 20499 -6917 20523 -6861
rect 20579 -6917 20623 -6861
rect 20323 -14065 20623 -6917
rect 21141 -13126 21442 -5978
rect 27892 -5622 28192 11540
rect 28404 -2633 28704 16953
rect 28903 17209 29203 17231
rect 28903 17153 28947 17209
rect 29003 17153 29027 17209
rect 29083 17153 29107 17209
rect 29163 17153 29203 17209
rect 28903 17109 29203 17153
rect 28903 17053 28947 17109
rect 29003 17053 29027 17109
rect 29083 17053 29107 17109
rect 29163 17053 29203 17109
rect 28903 17009 29203 17053
rect 28903 16953 28947 17009
rect 29003 16953 29027 17009
rect 29083 16953 29107 17009
rect 29163 16953 29203 17009
rect 28903 -2633 29203 16953
rect 27892 -5678 27936 -5622
rect 27992 -5678 28016 -5622
rect 28072 -5678 28096 -5622
rect 28152 -5678 28192 -5622
rect 27892 -5722 28192 -5678
rect 27892 -5778 27936 -5722
rect 27992 -5778 28016 -5722
rect 28072 -5778 28096 -5722
rect 28152 -5778 28192 -5722
rect 27892 -5822 28192 -5778
rect 27892 -5878 27936 -5822
rect 27992 -5878 28016 -5822
rect 28072 -5878 28096 -5822
rect 28152 -5878 28192 -5822
rect 27892 -5922 28192 -5878
rect 27892 -5978 27936 -5922
rect 27992 -5978 28016 -5922
rect 28072 -5978 28096 -5922
rect 28152 -5978 28192 -5922
rect 27892 -6000 28192 -5978
rect 22917 -7688 23217 -7666
rect 22917 -7744 22961 -7688
rect 23017 -7744 23041 -7688
rect 23097 -7744 23121 -7688
rect 23177 -7744 23217 -7688
rect 22917 -7788 23217 -7744
rect 22917 -7844 22961 -7788
rect 23017 -7844 23041 -7788
rect 23097 -7844 23121 -7788
rect 23177 -7844 23217 -7788
rect 22917 -7888 23217 -7844
rect 22917 -7944 22961 -7888
rect 23017 -7944 23041 -7888
rect 23097 -7944 23121 -7888
rect 23177 -7944 23217 -7888
rect 22917 -7988 23217 -7944
rect 22917 -8044 22961 -7988
rect 23017 -8044 23041 -7988
rect 23097 -8044 23121 -7988
rect 23177 -8044 23217 -7988
rect 22917 -8066 23217 -8044
rect 29759 -7688 30059 -1868
rect 29759 -7744 29803 -7688
rect 29859 -7744 29883 -7688
rect 29939 -7744 29963 -7688
rect 30019 -7744 30059 -7688
rect 29759 -7788 30059 -7744
rect 29759 -7844 29803 -7788
rect 29859 -7844 29883 -7788
rect 29939 -7844 29963 -7788
rect 30019 -7844 30059 -7788
rect 29759 -7888 30059 -7844
rect 29759 -7944 29803 -7888
rect 29859 -7944 29883 -7888
rect 29939 -7944 29963 -7888
rect 30019 -7944 30059 -7888
rect 29759 -7988 30059 -7944
rect 29759 -8044 29803 -7988
rect 29859 -8044 29883 -7988
rect 29939 -8044 29963 -7988
rect 30019 -8044 30059 -7988
rect 29034 -8424 29334 -8402
rect 29034 -8480 29078 -8424
rect 29134 -8480 29158 -8424
rect 29214 -8480 29238 -8424
rect 29294 -8480 29334 -8424
rect 29034 -8524 29334 -8480
rect 29034 -8580 29078 -8524
rect 29134 -8580 29158 -8524
rect 29214 -8580 29238 -8524
rect 29294 -8580 29334 -8524
rect 29034 -8624 29334 -8580
rect 29034 -8680 29078 -8624
rect 29134 -8680 29158 -8624
rect 29214 -8680 29238 -8624
rect 29294 -8680 29334 -8624
rect 29034 -8724 29334 -8680
rect 29034 -8780 29078 -8724
rect 29134 -8780 29158 -8724
rect 29214 -8780 29238 -8724
rect 29294 -8780 29334 -8724
rect 22917 -10062 23217 -10040
rect 22917 -10118 22961 -10062
rect 23017 -10118 23041 -10062
rect 23097 -10118 23121 -10062
rect 23177 -10118 23217 -10062
rect 22917 -10162 23217 -10118
rect 22917 -10218 22961 -10162
rect 23017 -10218 23041 -10162
rect 23097 -10218 23121 -10162
rect 23177 -10218 23217 -10162
rect 22917 -10262 23217 -10218
rect 22917 -10318 22961 -10262
rect 23017 -10318 23041 -10262
rect 23097 -10318 23121 -10262
rect 23177 -10318 23217 -10262
rect 22917 -10362 23217 -10318
rect 22917 -10418 22961 -10362
rect 23017 -10418 23041 -10362
rect 23097 -10418 23121 -10362
rect 23177 -10418 23217 -10362
rect 22917 -10440 23217 -10418
rect 22026 -14705 22326 -14683
rect 22026 -14761 22070 -14705
rect 22126 -14761 22150 -14705
rect 22206 -14761 22230 -14705
rect 22286 -14761 22326 -14705
rect 22026 -14805 22326 -14761
rect 22026 -14861 22070 -14805
rect 22126 -14861 22150 -14805
rect 22206 -14861 22230 -14805
rect 22286 -14861 22326 -14805
rect 22026 -14905 22326 -14861
rect 22026 -14961 22070 -14905
rect 22126 -14961 22150 -14905
rect 22206 -14961 22230 -14905
rect 22286 -14961 22326 -14905
rect 22026 -15005 22326 -14961
rect 22026 -15061 22070 -15005
rect 22126 -15061 22150 -15005
rect 22206 -15061 22230 -15005
rect 22286 -15061 22326 -15005
rect 22026 -15083 22326 -15061
rect 24861 -15700 25162 -15678
rect 24861 -15756 24906 -15700
rect 24962 -15756 24986 -15700
rect 25042 -15756 25066 -15700
rect 25122 -15756 25162 -15700
rect 24861 -15800 25162 -15756
rect 18542 -15864 18843 -15842
rect 18542 -15920 18587 -15864
rect 18643 -15920 18667 -15864
rect 18723 -15920 18747 -15864
rect 18803 -15920 18843 -15864
rect 18542 -16300 18843 -15920
rect 18542 -16356 18583 -16300
rect 18639 -16356 18663 -16300
rect 18719 -16356 18743 -16300
rect 18799 -16356 18843 -16300
rect 18542 -17275 18843 -16356
rect 18542 -17331 18583 -17275
rect 18639 -17331 18663 -17275
rect 18719 -17331 18743 -17275
rect 18799 -17331 18843 -17275
rect 18542 -17375 18843 -17331
rect 18542 -17431 18583 -17375
rect 18639 -17431 18663 -17375
rect 18719 -17431 18743 -17375
rect 18799 -17431 18843 -17375
rect 18542 -17475 18843 -17431
rect 18542 -17531 18583 -17475
rect 18639 -17531 18663 -17475
rect 18719 -17531 18743 -17475
rect 18799 -17531 18843 -17475
rect 18542 -17553 18843 -17531
rect 24861 -15856 24906 -15800
rect 24962 -15856 24986 -15800
rect 25042 -15856 25066 -15800
rect 25122 -15856 25162 -15800
rect 24861 -15900 25162 -15856
rect 24861 -15956 24906 -15900
rect 24962 -15956 24986 -15900
rect 25042 -15956 25066 -15900
rect 25122 -15956 25162 -15900
rect 24861 -16000 25162 -15956
rect 24861 -16056 24906 -16000
rect 24962 -16056 24986 -16000
rect 25042 -16056 25066 -16000
rect 25122 -16056 25162 -16000
rect 24861 -17275 25162 -16056
rect 29034 -15700 29334 -8780
rect 29759 -10062 30059 -8044
rect 29759 -10118 29803 -10062
rect 29859 -10118 29883 -10062
rect 29939 -10118 29963 -10062
rect 30019 -10118 30059 -10062
rect 29759 -10162 30059 -10118
rect 29759 -10218 29803 -10162
rect 29859 -10218 29883 -10162
rect 29939 -10218 29963 -10162
rect 30019 -10218 30059 -10162
rect 29759 -10262 30059 -10218
rect 29759 -10318 29803 -10262
rect 29859 -10318 29883 -10262
rect 29939 -10318 29963 -10262
rect 30019 -10318 30059 -10262
rect 29759 -10362 30059 -10318
rect 29759 -10418 29803 -10362
rect 29859 -10418 29883 -10362
rect 29939 -10418 29963 -10362
rect 30019 -10418 30059 -10362
rect 29759 -14982 30059 -10418
rect 31012 -14270 31313 -12834
rect 31012 -14326 31057 -14270
rect 31113 -14326 31137 -14270
rect 31193 -14326 31217 -14270
rect 31273 -14326 31313 -14270
rect 31012 -14370 31313 -14326
rect 31012 -14426 31057 -14370
rect 31113 -14426 31137 -14370
rect 31193 -14426 31217 -14370
rect 31273 -14426 31313 -14370
rect 31012 -14470 31313 -14426
rect 31012 -14526 31057 -14470
rect 31113 -14526 31137 -14470
rect 31193 -14526 31217 -14470
rect 31273 -14526 31313 -14470
rect 31012 -14570 31313 -14526
rect 31012 -14626 31057 -14570
rect 31113 -14626 31137 -14570
rect 31193 -14626 31217 -14570
rect 31273 -14626 31313 -14570
rect 31012 -14648 31313 -14626
rect 39403 -14270 39703 -12834
rect 39403 -14326 39447 -14270
rect 39503 -14326 39527 -14270
rect 39583 -14326 39607 -14270
rect 39663 -14326 39703 -14270
rect 39403 -14370 39703 -14326
rect 39403 -14426 39447 -14370
rect 39503 -14426 39527 -14370
rect 39583 -14426 39607 -14370
rect 39663 -14426 39703 -14370
rect 39403 -14470 39703 -14426
rect 39403 -14526 39447 -14470
rect 39503 -14526 39527 -14470
rect 39583 -14526 39607 -14470
rect 39663 -14526 39703 -14470
rect 39403 -14570 39703 -14526
rect 39403 -14626 39447 -14570
rect 39503 -14626 39527 -14570
rect 39583 -14626 39607 -14570
rect 39663 -14626 39703 -14570
rect 39403 -14648 39703 -14626
rect 29759 -15038 29803 -14982
rect 29859 -15038 29883 -14982
rect 29939 -15038 29963 -14982
rect 30019 -15038 30059 -14982
rect 29759 -15082 30059 -15038
rect 29759 -15138 29803 -15082
rect 29859 -15138 29883 -15082
rect 29939 -15138 29963 -15082
rect 30019 -15138 30059 -15082
rect 29759 -15182 30059 -15138
rect 29759 -15238 29803 -15182
rect 29859 -15238 29883 -15182
rect 29939 -15238 29963 -15182
rect 30019 -15238 30059 -15182
rect 29759 -15282 30059 -15238
rect 29759 -15338 29803 -15282
rect 29859 -15338 29883 -15282
rect 29939 -15338 29963 -15282
rect 30019 -15338 30059 -15282
rect 29759 -15360 30059 -15338
rect 40262 -14982 40562 -1868
rect 42474 -4666 42774 -4644
rect 42474 -4722 42514 -4666
rect 42570 -4722 42594 -4666
rect 42650 -4722 42674 -4666
rect 42730 -4722 42774 -4666
rect 42474 -4766 42774 -4722
rect 42474 -4822 42514 -4766
rect 42570 -4822 42594 -4766
rect 42650 -4822 42674 -4766
rect 42730 -4822 42774 -4766
rect 42474 -4866 42774 -4822
rect 42474 -4922 42514 -4866
rect 42570 -4922 42594 -4866
rect 42650 -4922 42674 -4866
rect 42730 -4922 42774 -4866
rect 42474 -4966 42774 -4922
rect 42474 -5022 42514 -4966
rect 42570 -5022 42594 -4966
rect 42650 -5022 42674 -4966
rect 42730 -5022 42774 -4966
rect 42474 -5044 42774 -5022
rect 40262 -15038 40306 -14982
rect 40362 -15038 40386 -14982
rect 40442 -15038 40466 -14982
rect 40522 -15038 40562 -14982
rect 40262 -15082 40562 -15038
rect 40262 -15138 40306 -15082
rect 40362 -15138 40386 -15082
rect 40442 -15138 40466 -15082
rect 40522 -15138 40562 -15082
rect 40262 -15182 40562 -15138
rect 40262 -15238 40306 -15182
rect 40362 -15238 40386 -15182
rect 40442 -15238 40466 -15182
rect 40522 -15238 40562 -15182
rect 40262 -15282 40562 -15238
rect 40262 -15338 40306 -15282
rect 40362 -15338 40386 -15282
rect 40442 -15338 40466 -15282
rect 40522 -15338 40562 -15282
rect 40262 -15360 40562 -15338
rect 40996 -8424 41296 -8402
rect 40996 -8480 41036 -8424
rect 41092 -8480 41116 -8424
rect 41172 -8480 41196 -8424
rect 41252 -8480 41296 -8424
rect 40996 -8524 41296 -8480
rect 40996 -8580 41036 -8524
rect 41092 -8580 41116 -8524
rect 41172 -8580 41196 -8524
rect 41252 -8580 41296 -8524
rect 40996 -8624 41296 -8580
rect 40996 -8680 41036 -8624
rect 41092 -8680 41116 -8624
rect 41172 -8680 41196 -8624
rect 41252 -8680 41296 -8624
rect 40996 -8724 41296 -8680
rect 40996 -8780 41036 -8724
rect 41092 -8780 41116 -8724
rect 41172 -8780 41196 -8724
rect 41252 -8780 41296 -8724
rect 29034 -15756 29078 -15700
rect 29134 -15756 29158 -15700
rect 29214 -15756 29238 -15700
rect 29294 -15756 29334 -15700
rect 29034 -15800 29334 -15756
rect 29034 -15856 29078 -15800
rect 29134 -15856 29158 -15800
rect 29214 -15856 29238 -15800
rect 29294 -15856 29334 -15800
rect 29034 -15900 29334 -15856
rect 29034 -15956 29078 -15900
rect 29134 -15956 29158 -15900
rect 29214 -15956 29238 -15900
rect 29294 -15956 29334 -15900
rect 29034 -16000 29334 -15956
rect 29034 -16056 29078 -16000
rect 29134 -16056 29158 -16000
rect 29214 -16056 29238 -16000
rect 29294 -16056 29334 -16000
rect 29034 -16078 29334 -16056
rect 40996 -15700 41296 -8780
rect 41986 -14982 42286 -7834
rect 42913 -14270 43213 -12834
rect 42913 -14326 42957 -14270
rect 43013 -14326 43037 -14270
rect 43093 -14326 43117 -14270
rect 43173 -14326 43213 -14270
rect 42913 -14370 43213 -14326
rect 42913 -14426 42957 -14370
rect 43013 -14426 43037 -14370
rect 43093 -14426 43117 -14370
rect 43173 -14426 43213 -14370
rect 42913 -14470 43213 -14426
rect 42913 -14526 42957 -14470
rect 43013 -14526 43037 -14470
rect 43093 -14526 43117 -14470
rect 43173 -14526 43213 -14470
rect 42913 -14570 43213 -14526
rect 42913 -14626 42957 -14570
rect 43013 -14626 43037 -14570
rect 43093 -14626 43117 -14570
rect 43173 -14626 43213 -14570
rect 42913 -14648 43213 -14626
rect 51303 -14270 51603 -12834
rect 51303 -14326 51347 -14270
rect 51403 -14326 51427 -14270
rect 51483 -14326 51507 -14270
rect 51563 -14326 51603 -14270
rect 51303 -14370 51603 -14326
rect 51303 -14426 51347 -14370
rect 51403 -14426 51427 -14370
rect 51483 -14426 51507 -14370
rect 51563 -14426 51603 -14370
rect 51303 -14470 51603 -14426
rect 51303 -14526 51347 -14470
rect 51403 -14526 51427 -14470
rect 51483 -14526 51507 -14470
rect 51563 -14526 51603 -14470
rect 51303 -14570 51603 -14526
rect 51303 -14626 51347 -14570
rect 51403 -14626 51427 -14570
rect 51483 -14626 51507 -14570
rect 51563 -14626 51603 -14570
rect 51303 -14648 51603 -14626
rect 41986 -15038 42030 -14982
rect 42086 -15038 42110 -14982
rect 42166 -15038 42190 -14982
rect 42246 -15038 42286 -14982
rect 41986 -15082 42286 -15038
rect 41986 -15138 42030 -15082
rect 42086 -15138 42110 -15082
rect 42166 -15138 42190 -15082
rect 42246 -15138 42286 -15082
rect 41986 -15182 42286 -15138
rect 41986 -15238 42030 -15182
rect 42086 -15238 42110 -15182
rect 42166 -15238 42190 -15182
rect 42246 -15238 42286 -15182
rect 41986 -15282 42286 -15238
rect 41986 -15338 42030 -15282
rect 42086 -15338 42110 -15282
rect 42166 -15338 42190 -15282
rect 42246 -15338 42286 -15282
rect 41986 -15360 42286 -15338
rect 52316 -14982 52617 -7834
rect 52316 -15038 52360 -14982
rect 52416 -15038 52440 -14982
rect 52496 -15038 52520 -14982
rect 52576 -15038 52617 -14982
rect 52316 -15082 52617 -15038
rect 52316 -15138 52360 -15082
rect 52416 -15138 52440 -15082
rect 52496 -15138 52520 -15082
rect 52576 -15138 52617 -15082
rect 52316 -15182 52617 -15138
rect 52316 -15238 52360 -15182
rect 52416 -15238 52440 -15182
rect 52496 -15238 52520 -15182
rect 52576 -15238 52617 -15182
rect 52316 -15282 52617 -15238
rect 52316 -15338 52360 -15282
rect 52416 -15338 52440 -15282
rect 52496 -15338 52520 -15282
rect 52576 -15338 52617 -15282
rect 52316 -15360 52617 -15338
rect 40996 -15756 41040 -15700
rect 41096 -15756 41120 -15700
rect 41176 -15756 41200 -15700
rect 41256 -15756 41296 -15700
rect 40996 -15800 41296 -15756
rect 40996 -15856 41040 -15800
rect 41096 -15856 41120 -15800
rect 41176 -15856 41200 -15800
rect 41256 -15856 41296 -15800
rect 40996 -15900 41296 -15856
rect 40996 -15956 41040 -15900
rect 41096 -15956 41120 -15900
rect 41176 -15956 41200 -15900
rect 41256 -15956 41296 -15900
rect 40996 -16000 41296 -15956
rect 40996 -16056 41040 -16000
rect 41096 -16056 41120 -16000
rect 41176 -16056 41200 -16000
rect 41256 -16056 41296 -16000
rect 40996 -16078 41296 -16056
rect 24861 -17331 24902 -17275
rect 24958 -17331 24982 -17275
rect 25038 -17331 25062 -17275
rect 25118 -17331 25162 -17275
rect 24861 -17375 25162 -17331
rect 24861 -17431 24902 -17375
rect 24958 -17431 24982 -17375
rect 25038 -17431 25062 -17375
rect 25118 -17431 25162 -17375
rect 24861 -17475 25162 -17431
rect 24861 -17531 24902 -17475
rect 24958 -17531 24982 -17475
rect 25038 -17531 25062 -17475
rect 25118 -17531 25162 -17475
rect 24861 -17553 25162 -17531
use bias  bias_0
timestamp 1698888477
transform 1 0 11885 0 1 -14246
box 290 -4088 13796 7675
use dda  dda_0
timestamp 1698888477
transform 1 0 34509 0 1 3684
box -27032 -18271 18695 11936
use diode  diode_0
timestamp 1698888477
transform 0 -1 7509 1 0 17069
box -701 208 -355 554
use diode  diode_1
timestamp 1698888477
transform 0 -1 8008 1 0 17069
box -701 208 -355 554
use diode  diode_2
timestamp 1698888477
transform 0 -1 8506 1 0 17069
box -701 208 -355 554
use diode  diode_3
timestamp 1698888477
transform 0 -1 28935 1 0 17069
box -701 208 -355 554
use diode  diode_4
timestamp 1698888477
transform 0 -1 29433 1 0 17069
box -701 208 -355 554
use diode  diode_5
timestamp 1698888477
transform 1 0 54981 0 1 -5222
box -701 208 -355 554
use diode  diode_6
timestamp 1698888477
transform -1 0 52013 0 -1 -14778
box -701 208 -355 554
use diode  diode_7
timestamp 1698888477
transform 1 0 54998 0 1 -5770
box -701 208 -355 554
<< labels >>
flabel metal2 s 27735 -14463 27735 -14463 2 FreeSans 3126 0 0 0 VB2
flabel metal2 s 33748 -15180 33748 -15180 2 FreeSans 3126 0 0 0 VB4
flabel metal2 s 34024 -15896 34024 -15896 2 FreeSans 3126 0 0 0 VB3
flabel metal2 s 18228 -5911 18228 -5911 2 FreeSans 3126 0 0 0 VB1
flabel metal2 s 53433 -5555 54650 -5218 2 FreeSans 3126 0 0 0 VO2
port 1 nsew
flabel metal2 s 54041 -5386 54041 -5386 2 FreeSans 3126 0 0 0 VO2
flabel metal2 s 28907 17282 29197 17402 2 FreeSans 3126 0 0 0 VI_2A
port 2 nsew
flabel metal2 s 28435 17249 28680 17402 2 FreeSans 3126 0 0 0 VI_2B
port 3 nsew
flabel metal2 s 7991 17317 8262 17439 2 FreeSans 3126 0 0 0 VI_1B
port 4 nsew
flabel metal2 s 7519 17321 7743 17437 2 FreeSans 3126 0 0 0 VI_1A
port 5 nsew
flabel metal2 s 7015 17331 7233 17428 2 FreeSans 3126 0 0 0 IREF
port 6 nsew
flabel metal2 s 42965 -15318 51605 -14983 2 FreeSans 3126 0 0 0 VCM
port 7 nsew
flabel metal2 s 53422 -5012 54634 -4670 2 FreeSans 3126 0 0 0 VO1
port 8 nsew
flabel metal2 s 52185 15258 53090 15540 2 FreeSans 3126 0 0 0 AVDD
port 9 nsew
flabel metal2 s 39277 15922 50288 16168 2 FreeSans 3126 0 0 0 AVSS
port 10 nsew
<< end >>
