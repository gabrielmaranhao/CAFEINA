magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< pwell >>
rect 2121 -118 2747 134
<< nmos >>
rect 2205 -92 2405 108
rect 2463 -92 2663 108
<< ndiff >>
rect 2147 93 2205 108
rect 2147 59 2159 93
rect 2193 59 2205 93
rect 2147 25 2205 59
rect 2147 -9 2159 25
rect 2193 -9 2205 25
rect 2147 -43 2205 -9
rect 2147 -77 2159 -43
rect 2193 -77 2205 -43
rect 2147 -92 2205 -77
rect 2405 93 2463 108
rect 2405 59 2417 93
rect 2451 59 2463 93
rect 2405 25 2463 59
rect 2405 -9 2417 25
rect 2451 -9 2463 25
rect 2405 -43 2463 -9
rect 2405 -77 2417 -43
rect 2451 -77 2463 -43
rect 2405 -92 2463 -77
rect 2663 93 2721 108
rect 2663 59 2675 93
rect 2709 59 2721 93
rect 2663 25 2721 59
rect 2663 -9 2675 25
rect 2709 -9 2721 25
rect 2663 -43 2721 -9
rect 2663 -77 2675 -43
rect 2709 -77 2721 -43
rect 2663 -92 2721 -77
<< ndiffc >>
rect 2159 59 2193 93
rect 2159 -9 2193 25
rect 2159 -77 2193 -43
rect 2417 59 2451 93
rect 2417 -9 2451 25
rect 2417 -77 2451 -43
rect 2675 59 2709 93
rect 2675 -9 2709 25
rect 2675 -77 2709 -43
<< poly >>
rect 2205 180 2405 196
rect 2205 146 2254 180
rect 2288 146 2322 180
rect 2356 146 2405 180
rect 2205 108 2405 146
rect 2463 180 2663 196
rect 2463 146 2512 180
rect 2546 146 2580 180
rect 2614 146 2663 180
rect 2463 108 2663 146
rect 2205 -118 2405 -92
rect 2463 -118 2663 -92
<< polycont >>
rect 2254 146 2288 180
rect 2322 146 2356 180
rect 2512 146 2546 180
rect 2580 146 2614 180
<< locali >>
rect 2205 146 2252 180
rect 2288 146 2322 180
rect 2358 146 2405 180
rect 2463 146 2510 180
rect 2546 146 2580 180
rect 2616 146 2663 180
rect 2159 93 2193 112
rect 2159 25 2193 27
rect 2159 -11 2193 -9
rect 2159 -96 2193 -77
rect 2417 93 2451 112
rect 2417 25 2451 27
rect 2417 -11 2451 -9
rect 2417 -96 2451 -77
rect 2675 93 2709 112
rect 2675 25 2709 27
rect 2675 -11 2709 -9
rect 2675 -96 2709 -77
<< viali >>
rect 2252 146 2254 180
rect 2254 146 2286 180
rect 2324 146 2356 180
rect 2356 146 2358 180
rect 2510 146 2512 180
rect 2512 146 2544 180
rect 2582 146 2614 180
rect 2614 146 2616 180
rect 2159 59 2193 61
rect 2159 27 2193 59
rect 2159 -43 2193 -11
rect 2159 -45 2193 -43
rect 2417 59 2451 61
rect 2417 27 2451 59
rect 2417 -43 2451 -11
rect 2417 -45 2451 -43
rect 2675 59 2709 61
rect 2675 27 2709 59
rect 2675 -43 2709 -11
rect 2675 -45 2709 -43
<< metal1 >>
rect 2209 180 2659 186
rect 2209 146 2252 180
rect 2286 146 2324 180
rect 2358 146 2510 180
rect 2544 146 2582 180
rect 2616 146 2659 180
rect 2209 140 2659 146
rect 2153 61 2199 108
rect 2153 27 2159 61
rect 2193 27 2199 61
rect 2153 -11 2199 27
rect 2153 -45 2159 -11
rect 2193 -45 2199 -11
rect 2153 -92 2199 -45
rect 2411 61 2457 108
rect 2411 27 2417 61
rect 2451 27 2457 61
rect 2411 -11 2457 27
rect 2411 -45 2417 -11
rect 2451 -45 2457 -11
rect 2411 -92 2457 -45
rect 2669 61 2715 108
rect 2669 27 2675 61
rect 2709 27 2715 61
rect 2669 -11 2715 27
rect 2669 -45 2675 -11
rect 2709 -45 2715 -11
rect 2669 -92 2715 -45
<< end >>
