magic
tech sky130A
magscale 1 2
timestamp 1698351692
<< pwell >>
rect -952 -448 952 448
<< mvnmos >>
rect -734 -200 -574 200
rect -516 -200 -356 200
rect -298 -200 -138 200
rect -80 -200 80 200
rect 138 -200 298 200
rect 356 -200 516 200
rect 574 -200 734 200
<< mvndiff >>
rect -792 187 -734 200
rect -792 153 -780 187
rect -746 153 -734 187
rect -792 119 -734 153
rect -792 85 -780 119
rect -746 85 -734 119
rect -792 51 -734 85
rect -792 17 -780 51
rect -746 17 -734 51
rect -792 -17 -734 17
rect -792 -51 -780 -17
rect -746 -51 -734 -17
rect -792 -85 -734 -51
rect -792 -119 -780 -85
rect -746 -119 -734 -85
rect -792 -153 -734 -119
rect -792 -187 -780 -153
rect -746 -187 -734 -153
rect -792 -200 -734 -187
rect -574 187 -516 200
rect -574 153 -562 187
rect -528 153 -516 187
rect -574 119 -516 153
rect -574 85 -562 119
rect -528 85 -516 119
rect -574 51 -516 85
rect -574 17 -562 51
rect -528 17 -516 51
rect -574 -17 -516 17
rect -574 -51 -562 -17
rect -528 -51 -516 -17
rect -574 -85 -516 -51
rect -574 -119 -562 -85
rect -528 -119 -516 -85
rect -574 -153 -516 -119
rect -574 -187 -562 -153
rect -528 -187 -516 -153
rect -574 -200 -516 -187
rect -356 187 -298 200
rect -356 153 -344 187
rect -310 153 -298 187
rect -356 119 -298 153
rect -356 85 -344 119
rect -310 85 -298 119
rect -356 51 -298 85
rect -356 17 -344 51
rect -310 17 -298 51
rect -356 -17 -298 17
rect -356 -51 -344 -17
rect -310 -51 -298 -17
rect -356 -85 -298 -51
rect -356 -119 -344 -85
rect -310 -119 -298 -85
rect -356 -153 -298 -119
rect -356 -187 -344 -153
rect -310 -187 -298 -153
rect -356 -200 -298 -187
rect -138 187 -80 200
rect -138 153 -126 187
rect -92 153 -80 187
rect -138 119 -80 153
rect -138 85 -126 119
rect -92 85 -80 119
rect -138 51 -80 85
rect -138 17 -126 51
rect -92 17 -80 51
rect -138 -17 -80 17
rect -138 -51 -126 -17
rect -92 -51 -80 -17
rect -138 -85 -80 -51
rect -138 -119 -126 -85
rect -92 -119 -80 -85
rect -138 -153 -80 -119
rect -138 -187 -126 -153
rect -92 -187 -80 -153
rect -138 -200 -80 -187
rect 80 187 138 200
rect 80 153 92 187
rect 126 153 138 187
rect 80 119 138 153
rect 80 85 92 119
rect 126 85 138 119
rect 80 51 138 85
rect 80 17 92 51
rect 126 17 138 51
rect 80 -17 138 17
rect 80 -51 92 -17
rect 126 -51 138 -17
rect 80 -85 138 -51
rect 80 -119 92 -85
rect 126 -119 138 -85
rect 80 -153 138 -119
rect 80 -187 92 -153
rect 126 -187 138 -153
rect 80 -200 138 -187
rect 298 187 356 200
rect 298 153 310 187
rect 344 153 356 187
rect 298 119 356 153
rect 298 85 310 119
rect 344 85 356 119
rect 298 51 356 85
rect 298 17 310 51
rect 344 17 356 51
rect 298 -17 356 17
rect 298 -51 310 -17
rect 344 -51 356 -17
rect 298 -85 356 -51
rect 298 -119 310 -85
rect 344 -119 356 -85
rect 298 -153 356 -119
rect 298 -187 310 -153
rect 344 -187 356 -153
rect 298 -200 356 -187
rect 516 187 574 200
rect 516 153 528 187
rect 562 153 574 187
rect 516 119 574 153
rect 516 85 528 119
rect 562 85 574 119
rect 516 51 574 85
rect 516 17 528 51
rect 562 17 574 51
rect 516 -17 574 17
rect 516 -51 528 -17
rect 562 -51 574 -17
rect 516 -85 574 -51
rect 516 -119 528 -85
rect 562 -119 574 -85
rect 516 -153 574 -119
rect 516 -187 528 -153
rect 562 -187 574 -153
rect 516 -200 574 -187
rect 734 187 792 200
rect 734 153 746 187
rect 780 153 792 187
rect 734 119 792 153
rect 734 85 746 119
rect 780 85 792 119
rect 734 51 792 85
rect 734 17 746 51
rect 780 17 792 51
rect 734 -17 792 17
rect 734 -51 746 -17
rect 780 -51 792 -17
rect 734 -85 792 -51
rect 734 -119 746 -85
rect 780 -119 792 -85
rect 734 -153 792 -119
rect 734 -187 746 -153
rect 780 -187 792 -153
rect 734 -200 792 -187
<< mvndiffc >>
rect -780 153 -746 187
rect -780 85 -746 119
rect -780 17 -746 51
rect -780 -51 -746 -17
rect -780 -119 -746 -85
rect -780 -187 -746 -153
rect -562 153 -528 187
rect -562 85 -528 119
rect -562 17 -528 51
rect -562 -51 -528 -17
rect -562 -119 -528 -85
rect -562 -187 -528 -153
rect -344 153 -310 187
rect -344 85 -310 119
rect -344 17 -310 51
rect -344 -51 -310 -17
rect -344 -119 -310 -85
rect -344 -187 -310 -153
rect -126 153 -92 187
rect -126 85 -92 119
rect -126 17 -92 51
rect -126 -51 -92 -17
rect -126 -119 -92 -85
rect -126 -187 -92 -153
rect 92 153 126 187
rect 92 85 126 119
rect 92 17 126 51
rect 92 -51 126 -17
rect 92 -119 126 -85
rect 92 -187 126 -153
rect 310 153 344 187
rect 310 85 344 119
rect 310 17 344 51
rect 310 -51 344 -17
rect 310 -119 344 -85
rect 310 -187 344 -153
rect 528 153 562 187
rect 528 85 562 119
rect 528 17 562 51
rect 528 -51 562 -17
rect 528 -119 562 -85
rect 528 -187 562 -153
rect 746 153 780 187
rect 746 85 780 119
rect 746 17 780 51
rect 746 -51 780 -17
rect 746 -119 780 -85
rect 746 -187 780 -153
<< mvpsubdiff >>
rect -926 410 926 422
rect -926 376 -799 410
rect -765 376 -731 410
rect -697 376 -663 410
rect -629 376 -595 410
rect -561 376 -527 410
rect -493 376 -459 410
rect -425 376 -391 410
rect -357 376 -323 410
rect -289 376 -255 410
rect -221 376 -187 410
rect -153 376 -119 410
rect -85 376 -51 410
rect -17 376 17 410
rect 51 376 85 410
rect 119 376 153 410
rect 187 376 221 410
rect 255 376 289 410
rect 323 376 357 410
rect 391 376 425 410
rect 459 376 493 410
rect 527 376 561 410
rect 595 376 629 410
rect 663 376 697 410
rect 731 376 765 410
rect 799 376 926 410
rect -926 364 926 376
rect -926 289 -868 364
rect -926 255 -914 289
rect -880 255 -868 289
rect 868 289 926 364
rect -926 221 -868 255
rect -926 187 -914 221
rect -880 187 -868 221
rect 868 255 880 289
rect 914 255 926 289
rect 868 221 926 255
rect -926 153 -868 187
rect -926 119 -914 153
rect -880 119 -868 153
rect -926 85 -868 119
rect -926 51 -914 85
rect -880 51 -868 85
rect -926 17 -868 51
rect -926 -17 -914 17
rect -880 -17 -868 17
rect -926 -51 -868 -17
rect -926 -85 -914 -51
rect -880 -85 -868 -51
rect -926 -119 -868 -85
rect -926 -153 -914 -119
rect -880 -153 -868 -119
rect -926 -187 -868 -153
rect -926 -221 -914 -187
rect -880 -221 -868 -187
rect 868 187 880 221
rect 914 187 926 221
rect 868 153 926 187
rect 868 119 880 153
rect 914 119 926 153
rect 868 85 926 119
rect 868 51 880 85
rect 914 51 926 85
rect 868 17 926 51
rect 868 -17 880 17
rect 914 -17 926 17
rect 868 -51 926 -17
rect 868 -85 880 -51
rect 914 -85 926 -51
rect 868 -119 926 -85
rect 868 -153 880 -119
rect 914 -153 926 -119
rect 868 -187 926 -153
rect -926 -255 -868 -221
rect -926 -289 -914 -255
rect -880 -289 -868 -255
rect 868 -221 880 -187
rect 914 -221 926 -187
rect 868 -255 926 -221
rect -926 -364 -868 -289
rect 868 -289 880 -255
rect 914 -289 926 -255
rect 868 -364 926 -289
rect -926 -376 926 -364
rect -926 -410 -799 -376
rect -765 -410 -731 -376
rect -697 -410 -663 -376
rect -629 -410 -595 -376
rect -561 -410 -527 -376
rect -493 -410 -459 -376
rect -425 -410 -391 -376
rect -357 -410 -323 -376
rect -289 -410 -255 -376
rect -221 -410 -187 -376
rect -153 -410 -119 -376
rect -85 -410 -51 -376
rect -17 -410 17 -376
rect 51 -410 85 -376
rect 119 -410 153 -376
rect 187 -410 221 -376
rect 255 -410 289 -376
rect 323 -410 357 -376
rect 391 -410 425 -376
rect 459 -410 493 -376
rect 527 -410 561 -376
rect 595 -410 629 -376
rect 663 -410 697 -376
rect 731 -410 765 -376
rect 799 -410 926 -376
rect -926 -422 926 -410
<< mvpsubdiffcont >>
rect -799 376 -765 410
rect -731 376 -697 410
rect -663 376 -629 410
rect -595 376 -561 410
rect -527 376 -493 410
rect -459 376 -425 410
rect -391 376 -357 410
rect -323 376 -289 410
rect -255 376 -221 410
rect -187 376 -153 410
rect -119 376 -85 410
rect -51 376 -17 410
rect 17 376 51 410
rect 85 376 119 410
rect 153 376 187 410
rect 221 376 255 410
rect 289 376 323 410
rect 357 376 391 410
rect 425 376 459 410
rect 493 376 527 410
rect 561 376 595 410
rect 629 376 663 410
rect 697 376 731 410
rect 765 376 799 410
rect -914 255 -880 289
rect -914 187 -880 221
rect 880 255 914 289
rect -914 119 -880 153
rect -914 51 -880 85
rect -914 -17 -880 17
rect -914 -85 -880 -51
rect -914 -153 -880 -119
rect -914 -221 -880 -187
rect 880 187 914 221
rect 880 119 914 153
rect 880 51 914 85
rect 880 -17 914 17
rect 880 -85 914 -51
rect 880 -153 914 -119
rect -914 -289 -880 -255
rect 880 -221 914 -187
rect 880 -289 914 -255
rect -799 -410 -765 -376
rect -731 -410 -697 -376
rect -663 -410 -629 -376
rect -595 -410 -561 -376
rect -527 -410 -493 -376
rect -459 -410 -425 -376
rect -391 -410 -357 -376
rect -323 -410 -289 -376
rect -255 -410 -221 -376
rect -187 -410 -153 -376
rect -119 -410 -85 -376
rect -51 -410 -17 -376
rect 17 -410 51 -376
rect 85 -410 119 -376
rect 153 -410 187 -376
rect 221 -410 255 -376
rect 289 -410 323 -376
rect 357 -410 391 -376
rect 425 -410 459 -376
rect 493 -410 527 -376
rect 561 -410 595 -376
rect 629 -410 663 -376
rect 697 -410 731 -376
rect 765 -410 799 -376
<< poly >>
rect -734 272 -574 288
rect -734 238 -705 272
rect -671 238 -637 272
rect -603 238 -574 272
rect -734 200 -574 238
rect -516 272 -356 288
rect -516 238 -487 272
rect -453 238 -419 272
rect -385 238 -356 272
rect -516 200 -356 238
rect -298 272 -138 288
rect -298 238 -269 272
rect -235 238 -201 272
rect -167 238 -138 272
rect -298 200 -138 238
rect -80 272 80 288
rect -80 238 -51 272
rect -17 238 17 272
rect 51 238 80 272
rect -80 200 80 238
rect 138 272 298 288
rect 138 238 167 272
rect 201 238 235 272
rect 269 238 298 272
rect 138 200 298 238
rect 356 272 516 288
rect 356 238 385 272
rect 419 238 453 272
rect 487 238 516 272
rect 356 200 516 238
rect 574 272 734 288
rect 574 238 603 272
rect 637 238 671 272
rect 705 238 734 272
rect 574 200 734 238
rect -734 -238 -574 -200
rect -734 -272 -705 -238
rect -671 -272 -637 -238
rect -603 -272 -574 -238
rect -734 -288 -574 -272
rect -516 -238 -356 -200
rect -516 -272 -487 -238
rect -453 -272 -419 -238
rect -385 -272 -356 -238
rect -516 -288 -356 -272
rect -298 -238 -138 -200
rect -298 -272 -269 -238
rect -235 -272 -201 -238
rect -167 -272 -138 -238
rect -298 -288 -138 -272
rect -80 -238 80 -200
rect -80 -272 -51 -238
rect -17 -272 17 -238
rect 51 -272 80 -238
rect -80 -288 80 -272
rect 138 -238 298 -200
rect 138 -272 167 -238
rect 201 -272 235 -238
rect 269 -272 298 -238
rect 138 -288 298 -272
rect 356 -238 516 -200
rect 356 -272 385 -238
rect 419 -272 453 -238
rect 487 -272 516 -238
rect 356 -288 516 -272
rect 574 -238 734 -200
rect 574 -272 603 -238
rect 637 -272 671 -238
rect 705 -272 734 -238
rect 574 -288 734 -272
<< polycont >>
rect -705 238 -671 272
rect -637 238 -603 272
rect -487 238 -453 272
rect -419 238 -385 272
rect -269 238 -235 272
rect -201 238 -167 272
rect -51 238 -17 272
rect 17 238 51 272
rect 167 238 201 272
rect 235 238 269 272
rect 385 238 419 272
rect 453 238 487 272
rect 603 238 637 272
rect 671 238 705 272
rect -705 -272 -671 -238
rect -637 -272 -603 -238
rect -487 -272 -453 -238
rect -419 -272 -385 -238
rect -269 -272 -235 -238
rect -201 -272 -167 -238
rect -51 -272 -17 -238
rect 17 -272 51 -238
rect 167 -272 201 -238
rect 235 -272 269 -238
rect 385 -272 419 -238
rect 453 -272 487 -238
rect 603 -272 637 -238
rect 671 -272 705 -238
<< locali >>
rect -914 376 -799 410
rect -765 376 -731 410
rect -697 376 -663 410
rect -629 376 -595 410
rect -561 376 -527 410
rect -493 376 -459 410
rect -425 376 -391 410
rect -357 376 -323 410
rect -289 376 -255 410
rect -221 376 -187 410
rect -153 376 -119 410
rect -85 376 -51 410
rect -17 376 17 410
rect 51 376 85 410
rect 119 376 153 410
rect 187 376 221 410
rect 255 376 289 410
rect 323 376 357 410
rect 391 376 425 410
rect 459 376 493 410
rect 527 376 561 410
rect 595 376 629 410
rect 663 376 697 410
rect 731 376 765 410
rect 799 376 914 410
rect -914 289 -880 376
rect 880 289 914 376
rect -914 233 -880 255
rect -734 238 -707 272
rect -671 238 -637 272
rect -601 238 -574 272
rect -516 238 -489 272
rect -453 238 -419 272
rect -383 238 -356 272
rect -298 238 -271 272
rect -235 238 -201 272
rect -165 238 -138 272
rect -80 238 -53 272
rect -17 238 17 272
rect 53 238 80 272
rect 138 238 165 272
rect 201 238 235 272
rect 271 238 298 272
rect 356 238 383 272
rect 419 238 453 272
rect 489 238 516 272
rect 574 238 601 272
rect 637 238 671 272
rect 707 238 734 272
rect 880 221 914 255
rect -914 161 -880 187
rect -914 89 -880 119
rect -914 17 -880 51
rect -914 -51 -880 -17
rect -914 -119 -880 -89
rect -914 -187 -880 -161
rect -780 187 -746 204
rect -780 149 -746 153
rect -780 77 -746 85
rect -780 -17 -746 17
rect -780 -85 -746 -51
rect -780 -153 -746 -119
rect -780 -204 -746 -187
rect -562 187 -528 204
rect -562 119 -528 153
rect -562 51 -528 85
rect -562 -17 -528 17
rect -562 -85 -528 -77
rect -562 -153 -528 -149
rect -562 -204 -528 -187
rect -344 187 -310 204
rect -344 149 -310 153
rect -344 77 -310 85
rect -344 -17 -310 17
rect -344 -85 -310 -51
rect -344 -153 -310 -119
rect -344 -204 -310 -187
rect -126 187 -92 204
rect -126 119 -92 153
rect -126 51 -92 85
rect -126 -17 -92 17
rect -126 -85 -92 -77
rect -126 -153 -92 -149
rect -126 -204 -92 -187
rect 92 187 126 204
rect 92 149 126 153
rect 92 77 126 85
rect 92 -17 126 17
rect 92 -85 126 -51
rect 92 -153 126 -119
rect 92 -204 126 -187
rect 310 187 344 204
rect 310 119 344 153
rect 310 51 344 85
rect 310 -17 344 17
rect 310 -85 344 -77
rect 310 -153 344 -149
rect 310 -204 344 -187
rect 528 187 562 204
rect 528 149 562 153
rect 528 77 562 85
rect 528 -17 562 17
rect 528 -85 562 -51
rect 528 -153 562 -119
rect 528 -204 562 -187
rect 746 187 780 204
rect 746 119 780 153
rect 746 51 780 85
rect 746 -17 780 17
rect 746 -85 780 -77
rect 746 -153 780 -149
rect 746 -204 780 -187
rect 880 153 914 187
rect 880 85 914 119
rect 880 17 914 51
rect 880 -51 914 -17
rect 880 -119 914 -85
rect 880 -187 914 -153
rect -914 -255 -880 -233
rect -734 -272 -707 -238
rect -671 -272 -637 -238
rect -601 -272 -574 -238
rect -516 -272 -489 -238
rect -453 -272 -419 -238
rect -383 -272 -356 -238
rect -298 -272 -271 -238
rect -235 -272 -201 -238
rect -165 -272 -138 -238
rect -80 -272 -53 -238
rect -17 -272 17 -238
rect 53 -272 80 -238
rect 138 -272 165 -238
rect 201 -272 235 -238
rect 271 -272 298 -238
rect 356 -272 383 -238
rect 419 -272 453 -238
rect 489 -272 516 -238
rect 574 -272 601 -238
rect 637 -272 671 -238
rect 707 -272 734 -238
rect 880 -255 914 -221
rect -914 -376 -880 -289
rect 880 -376 914 -289
rect -914 -410 -799 -376
rect -765 -410 -731 -376
rect -697 -410 -663 -376
rect -629 -410 -595 -376
rect -561 -410 -527 -376
rect -493 -410 -459 -376
rect -425 -410 -391 -376
rect -357 -410 -323 -376
rect -289 -410 -255 -376
rect -221 -410 -187 -376
rect -153 -410 -119 -376
rect -85 -410 -51 -376
rect -17 -410 17 -376
rect 51 -410 85 -376
rect 119 -410 153 -376
rect 187 -410 221 -376
rect 255 -410 289 -376
rect 323 -410 357 -376
rect 391 -410 425 -376
rect 459 -410 493 -376
rect 527 -410 561 -376
rect 595 -410 629 -376
rect 663 -410 697 -376
rect 731 -410 765 -376
rect 799 -410 914 -376
<< viali >>
rect -707 238 -705 272
rect -705 238 -673 272
rect -635 238 -603 272
rect -603 238 -601 272
rect -489 238 -487 272
rect -487 238 -455 272
rect -417 238 -385 272
rect -385 238 -383 272
rect -271 238 -269 272
rect -269 238 -237 272
rect -199 238 -167 272
rect -167 238 -165 272
rect -53 238 -51 272
rect -51 238 -19 272
rect 19 238 51 272
rect 51 238 53 272
rect 165 238 167 272
rect 167 238 199 272
rect 237 238 269 272
rect 269 238 271 272
rect 383 238 385 272
rect 385 238 417 272
rect 455 238 487 272
rect 487 238 489 272
rect 601 238 603 272
rect 603 238 635 272
rect 673 238 705 272
rect 705 238 707 272
rect -914 221 -880 233
rect -914 199 -880 221
rect -914 153 -880 161
rect -914 127 -880 153
rect -914 85 -880 89
rect -914 55 -880 85
rect -914 -17 -880 17
rect -914 -85 -880 -55
rect -914 -89 -880 -85
rect -914 -153 -880 -127
rect -914 -161 -880 -153
rect -914 -221 -880 -199
rect -780 119 -746 149
rect -780 115 -746 119
rect -780 51 -746 77
rect -780 43 -746 51
rect -562 -51 -528 -43
rect -562 -77 -528 -51
rect -562 -119 -528 -115
rect -562 -149 -528 -119
rect -344 119 -310 149
rect -344 115 -310 119
rect -344 51 -310 77
rect -344 43 -310 51
rect -126 -51 -92 -43
rect -126 -77 -92 -51
rect -126 -119 -92 -115
rect -126 -149 -92 -119
rect 92 119 126 149
rect 92 115 126 119
rect 92 51 126 77
rect 92 43 126 51
rect 310 -51 344 -43
rect 310 -77 344 -51
rect 310 -119 344 -115
rect 310 -149 344 -119
rect 528 119 562 149
rect 528 115 562 119
rect 528 51 562 77
rect 528 43 562 51
rect 746 -51 780 -43
rect 746 -77 780 -51
rect 746 -119 780 -115
rect 746 -149 780 -119
rect -914 -233 -880 -221
rect -707 -272 -705 -238
rect -705 -272 -673 -238
rect -635 -272 -603 -238
rect -603 -272 -601 -238
rect -489 -272 -487 -238
rect -487 -272 -455 -238
rect -417 -272 -385 -238
rect -385 -272 -383 -238
rect -271 -272 -269 -238
rect -269 -272 -237 -238
rect -199 -272 -167 -238
rect -167 -272 -165 -238
rect -53 -272 -51 -238
rect -51 -272 -19 -238
rect 19 -272 51 -238
rect 51 -272 53 -238
rect 165 -272 167 -238
rect 167 -272 199 -238
rect 237 -272 269 -238
rect 269 -272 271 -238
rect 383 -272 385 -238
rect 385 -272 417 -238
rect 455 -272 487 -238
rect 487 -272 489 -238
rect 601 -272 603 -238
rect 603 -272 635 -238
rect 673 -272 705 -238
rect 705 -272 707 -238
<< metal1 >>
rect -920 233 -874 275
rect -920 199 -914 233
rect -880 199 -874 233
rect -730 272 -578 278
rect -730 238 -707 272
rect -673 238 -635 272
rect -601 238 -578 272
rect -730 232 -578 238
rect -512 272 -360 278
rect -512 238 -489 272
rect -455 238 -417 272
rect -383 238 -360 272
rect -512 232 -360 238
rect -294 272 -142 278
rect -294 238 -271 272
rect -237 238 -199 272
rect -165 238 -142 272
rect -294 232 -142 238
rect -76 272 76 278
rect -76 238 -53 272
rect -19 238 19 272
rect 53 238 76 272
rect -76 232 76 238
rect 142 272 294 278
rect 142 238 165 272
rect 199 238 237 272
rect 271 238 294 272
rect 142 232 294 238
rect 360 272 512 278
rect 360 238 383 272
rect 417 238 455 272
rect 489 238 512 272
rect 360 232 512 238
rect 578 272 730 278
rect 578 238 601 272
rect 635 238 673 272
rect 707 238 730 272
rect 578 232 730 238
rect -920 161 -874 199
rect -920 127 -914 161
rect -880 127 -874 161
rect -920 89 -874 127
rect -920 55 -914 89
rect -880 55 -874 89
rect -920 17 -874 55
rect -920 -17 -914 17
rect -880 -17 -874 17
rect -786 149 -740 183
rect -786 115 -780 149
rect -746 115 -740 149
rect -786 77 -740 115
rect -786 43 -780 77
rect -746 43 -740 77
rect -786 9 -740 43
rect -350 149 -304 183
rect -350 115 -344 149
rect -310 115 -304 149
rect -350 77 -304 115
rect -350 43 -344 77
rect -310 43 -304 77
rect -350 9 -304 43
rect 86 149 132 183
rect 86 115 92 149
rect 126 115 132 149
rect 86 77 132 115
rect 86 43 92 77
rect 126 43 132 77
rect 86 9 132 43
rect 522 149 568 183
rect 522 115 528 149
rect 562 115 568 149
rect 522 77 568 115
rect 522 43 528 77
rect 562 43 568 77
rect 522 9 568 43
rect -920 -55 -874 -17
rect -920 -89 -914 -55
rect -880 -89 -874 -55
rect -920 -127 -874 -89
rect -920 -161 -914 -127
rect -880 -161 -874 -127
rect -920 -199 -874 -161
rect -568 -43 -522 -9
rect -568 -77 -562 -43
rect -528 -77 -522 -43
rect -568 -115 -522 -77
rect -568 -149 -562 -115
rect -528 -149 -522 -115
rect -568 -183 -522 -149
rect -132 -43 -86 -9
rect -132 -77 -126 -43
rect -92 -77 -86 -43
rect -132 -115 -86 -77
rect -132 -149 -126 -115
rect -92 -149 -86 -115
rect -132 -183 -86 -149
rect 304 -43 350 -9
rect 304 -77 310 -43
rect 344 -77 350 -43
rect 304 -115 350 -77
rect 304 -149 310 -115
rect 344 -149 350 -115
rect 304 -183 350 -149
rect 740 -43 786 -9
rect 740 -77 746 -43
rect 780 -77 786 -43
rect 740 -115 786 -77
rect 740 -149 746 -115
rect 780 -149 786 -115
rect 740 -183 786 -149
rect -920 -233 -914 -199
rect -880 -233 -874 -199
rect -920 -275 -874 -233
rect -730 -238 -578 -232
rect -730 -272 -707 -238
rect -673 -272 -635 -238
rect -601 -272 -578 -238
rect -730 -278 -578 -272
rect -512 -238 -360 -232
rect -512 -272 -489 -238
rect -455 -272 -417 -238
rect -383 -272 -360 -238
rect -512 -278 -360 -272
rect -294 -238 -142 -232
rect -294 -272 -271 -238
rect -237 -272 -199 -238
rect -165 -272 -142 -238
rect -294 -278 -142 -272
rect -76 -238 76 -232
rect -76 -272 -53 -238
rect -19 -272 19 -238
rect 53 -272 76 -238
rect -76 -278 76 -272
rect 142 -238 294 -232
rect 142 -272 165 -238
rect 199 -272 237 -238
rect 271 -272 294 -238
rect 142 -278 294 -272
rect 360 -238 512 -232
rect 360 -272 383 -238
rect 417 -272 455 -238
rect 489 -272 512 -238
rect 360 -278 512 -272
rect 578 -238 730 -232
rect 578 -272 601 -238
rect 635 -272 673 -238
rect 707 -272 730 -238
rect 578 -278 730 -272
<< properties >>
string FIXED_BBOX -897 -393 897 393
<< end >>
