magic
tech sky130A
timestamp 1697634299
<< pwell >>
rect -752 -586 752 586
<< mvpsubdiff >>
rect -734 562 -498 568
rect -734 545 -680 562
rect -552 545 -498 562
rect -734 539 -498 545
rect -734 514 -705 539
rect -734 -514 -728 514
rect -711 -514 -705 514
rect -527 514 -498 539
rect -734 -539 -705 -514
rect -527 -514 -521 514
rect -504 -514 -498 514
rect -527 -539 -498 -514
rect -734 -545 -498 -539
rect -734 -562 -680 -545
rect -552 -562 -498 -545
rect -734 -568 -498 -562
rect -426 562 -190 568
rect -426 545 -372 562
rect -244 545 -190 562
rect -426 539 -190 545
rect -426 514 -397 539
rect -426 -514 -420 514
rect -403 -514 -397 514
rect -219 514 -190 539
rect -426 -539 -397 -514
rect -219 -514 -213 514
rect -196 -514 -190 514
rect -219 -539 -190 -514
rect -426 -545 -190 -539
rect -426 -562 -372 -545
rect -244 -562 -190 -545
rect -426 -568 -190 -562
rect -118 562 118 568
rect -118 545 -64 562
rect 64 545 118 562
rect -118 539 118 545
rect -118 514 -89 539
rect -118 -514 -112 514
rect -95 -514 -89 514
rect 89 514 118 539
rect -118 -539 -89 -514
rect 89 -514 95 514
rect 112 -514 118 514
rect 89 -539 118 -514
rect -118 -545 118 -539
rect -118 -562 -64 -545
rect 64 -562 118 -545
rect -118 -568 118 -562
rect 190 562 426 568
rect 190 545 244 562
rect 372 545 426 562
rect 190 539 426 545
rect 190 514 219 539
rect 190 -514 196 514
rect 213 -514 219 514
rect 397 514 426 539
rect 190 -539 219 -514
rect 397 -514 403 514
rect 420 -514 426 514
rect 397 -539 426 -514
rect 190 -545 426 -539
rect 190 -562 244 -545
rect 372 -562 426 -545
rect 190 -568 426 -562
rect 498 562 734 568
rect 498 545 552 562
rect 680 545 734 562
rect 498 539 734 545
rect 498 514 527 539
rect 498 -514 504 514
rect 521 -514 527 514
rect 705 514 734 539
rect 498 -539 527 -514
rect 705 -514 711 514
rect 728 -514 734 514
rect 705 -539 734 -514
rect 498 -545 734 -539
rect 498 -562 552 -545
rect 680 -562 734 -545
rect 498 -568 734 -562
<< mvpsubdiffcont >>
rect -680 545 -552 562
rect -728 -514 -711 514
rect -521 -514 -504 514
rect -680 -562 -552 -545
rect -372 545 -244 562
rect -420 -514 -403 514
rect -213 -514 -196 514
rect -372 -562 -244 -545
rect -64 545 64 562
rect -112 -514 -95 514
rect 95 -514 112 514
rect -64 -562 64 -545
rect 244 545 372 562
rect 196 -514 213 514
rect 403 -514 420 514
rect 244 -562 372 -545
rect 552 545 680 562
rect 504 -514 521 514
rect 711 -514 728 514
rect 552 -562 680 -545
<< mvndiode >>
rect -666 494 -566 500
rect -666 -494 -660 494
rect -572 -494 -566 494
rect -666 -500 -566 -494
rect -358 494 -258 500
rect -358 -494 -352 494
rect -264 -494 -258 494
rect -358 -500 -258 -494
rect -50 494 50 500
rect -50 -494 -44 494
rect 44 -494 50 494
rect -50 -500 50 -494
rect 258 494 358 500
rect 258 -494 264 494
rect 352 -494 358 494
rect 258 -500 358 -494
rect 566 494 666 500
rect 566 -494 572 494
rect 660 -494 666 494
rect 566 -500 666 -494
<< mvndiodec >>
rect -660 -494 -572 494
rect -352 -494 -264 494
rect -44 -494 44 494
rect 264 -494 352 494
rect 572 -494 660 494
<< locali >>
rect -728 545 -680 562
rect -552 545 -504 562
rect -728 514 -711 545
rect -521 514 -504 545
rect -660 494 -572 502
rect -660 -502 -572 -494
rect -728 -545 -711 -514
rect -521 -545 -504 -514
rect -728 -562 -680 -545
rect -552 -562 -504 -545
rect -420 545 -372 562
rect -244 545 -196 562
rect -420 514 -403 545
rect -213 514 -196 545
rect -352 494 -264 502
rect -352 -502 -264 -494
rect -420 -545 -403 -514
rect -213 -545 -196 -514
rect -420 -562 -372 -545
rect -244 -562 -196 -545
rect -112 545 -64 562
rect 64 545 112 562
rect -112 514 -95 545
rect 95 514 112 545
rect -44 494 44 502
rect -44 -502 44 -494
rect -112 -545 -95 -514
rect 95 -545 112 -514
rect -112 -562 -64 -545
rect 64 -562 112 -545
rect 196 545 244 562
rect 372 545 420 562
rect 196 514 213 545
rect 403 514 420 545
rect 264 494 352 502
rect 264 -502 352 -494
rect 196 -545 213 -514
rect 403 -545 420 -514
rect 196 -562 244 -545
rect 372 -562 420 -545
rect 504 545 552 562
rect 680 545 728 562
rect 504 514 521 545
rect 711 514 728 545
rect 572 494 660 502
rect 572 -502 660 -494
rect 504 -545 521 -514
rect 711 -545 728 -514
rect 504 -562 552 -545
rect 680 -562 728 -545
<< viali >>
rect -660 -494 -572 494
rect -352 -494 -264 494
rect -44 -494 44 494
rect 264 -494 352 494
rect 572 -494 660 494
<< metal1 >>
rect -663 494 -569 500
rect -663 -494 -660 494
rect -572 -494 -569 494
rect -663 -500 -569 -494
rect -355 494 -261 500
rect -355 -494 -352 494
rect -264 -494 -261 494
rect -355 -500 -261 -494
rect -47 494 47 500
rect -47 -494 -44 494
rect 44 -494 47 494
rect -47 -500 47 -494
rect 261 494 355 500
rect 261 -494 264 494
rect 352 -494 355 494
rect 261 -500 355 -494
rect 569 494 663 500
rect 569 -494 572 494
rect 660 -494 663 494
rect 569 -500 663 -494
<< properties >>
string FIXED_BBOX 512 -553 719 553
string gencell sky130_fd_pr__diode_pw2nd_11v0
string library sky130
string parameters w 1 l 10 area 10.0 peri 22.0 nx 5 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
