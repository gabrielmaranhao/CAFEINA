magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< pwell >>
rect -831 78 -485 424
<< psubdiff >>
rect -805 364 -709 398
rect -675 364 -641 398
rect -607 364 -511 398
rect -805 302 -771 364
rect -545 302 -511 364
rect -805 234 -771 268
rect -545 234 -511 268
rect -805 138 -771 200
rect -545 138 -511 200
rect -805 104 -709 138
rect -675 104 -641 138
rect -607 104 -511 138
<< psubdiffcont >>
rect -709 364 -675 398
rect -641 364 -607 398
rect -805 268 -771 302
rect -805 200 -771 234
rect -545 268 -511 302
rect -545 200 -511 234
rect -709 104 -675 138
rect -641 104 -607 138
<< ndiode >>
rect -703 268 -613 296
rect -703 234 -675 268
rect -641 234 -613 268
rect -703 206 -613 234
<< ndiodec >>
rect -675 234 -641 268
<< locali >>
rect -805 364 -709 398
rect -675 364 -641 398
rect -607 364 -511 398
rect -805 302 -771 364
rect -545 302 -511 364
rect -805 234 -771 268
rect -707 268 -609 284
rect -707 234 -675 268
rect -641 234 -609 268
rect -707 218 -609 234
rect -545 234 -511 268
rect -805 138 -771 200
rect -545 138 -511 200
rect -805 104 -709 138
rect -675 104 -641 138
rect -607 104 -511 138
<< viali >>
rect -675 234 -641 268
<< metal1 >>
rect -703 268 -613 290
rect -703 234 -675 268
rect -641 234 -613 268
rect -703 212 -613 234
<< properties >>
string FIXED_BBOX -788 121 -528 381
<< end >>
