** sch_path: /home/gmaranhao/Desktop/sky130_work/user_wrapper_caravan/user_analog_project_wrapper.sch
.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1] wbs_sel_i[0] wbs_dat_i[31]
+ wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26] wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23]
+ wbs_dat_i[22] wbs_dat_i[21] wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16] wbs_dat_i[15]
+ wbs_dat_i[14] wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8] wbs_dat_i[7]
+ wbs_dat_i[6] wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1] wbs_dat_i[0] wbs_adr_i[31]
+ wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28] wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23]
+ wbs_adr_i[22] wbs_adr_i[21] wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18] wbs_adr_i[17] wbs_adr_i[16] wbs_adr_i[15]
+ wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10] wbs_adr_i[9] wbs_adr_i[8] wbs_adr_i[7]
+ wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3] wbs_adr_i[2] wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o
+ wbs_dat_o[31] wbs_dat_o[30] wbs_dat_o[29] wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24]
+ wbs_dat_o[23] wbs_dat_o[22] wbs_dat_o[21] wbs_dat_o[20] wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16]
+ wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10] wbs_dat_o[9] wbs_dat_o[8]
+ wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4] wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0]
+ la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121]
+ la_data_in[120] la_data_in[119] la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114]
+ la_data_in[113] la_data_in[112] la_data_in[111] la_data_in[110] la_data_in[109] la_data_in[108] la_data_in[107]
+ la_data_in[106] la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102] la_data_in[101] la_data_in[100]
+ la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93]
+ la_data_in[92] la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86]
+ la_data_in[85] la_data_in[84] la_data_in[83] la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79]
+ la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75] la_data_in[74] la_data_in[73] la_data_in[72]
+ la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66] la_data_in[65]
+ la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58]
+ la_data_in[57] la_data_in[56] la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51]
+ la_data_in[50] la_data_in[49] la_data_in[48] la_data_in[47] la_data_in[46] la_data_in[45] la_data_in[44]
+ la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39] la_data_in[38] la_data_in[37]
+ la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30]
+ la_data_in[29] la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23]
+ la_data_in[22] la_data_in[21] la_data_in[20] la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16]
+ la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12] la_data_in[11] la_data_in[10] la_data_in[9]
+ la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2] la_data_in[1]
+ la_data_in[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124] la_data_out[123]
+ la_data_out[122] la_data_out[121] la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117]
+ la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113] la_data_out[112] la_data_out[111]
+ la_data_out[110] la_data_out[109] la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105]
+ la_data_out[104] la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98]
+ la_data_out[97] la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92] la_data_out[91]
+ la_data_out[90] la_data_out[89] la_data_out[88] la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84]
+ la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79] la_data_out[78] la_data_out[77]
+ la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70]
+ la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64] la_data_out[63]
+ la_data_out[62] la_data_out[61] la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56]
+ la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52] la_data_out[51] la_data_out[50] la_data_out[49]
+ la_data_out[48] la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43] la_data_out[42]
+ la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35]
+ la_data_out[34] la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28]
+ la_data_out[27] la_data_out[26] la_data_out[25] la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21]
+ la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17] la_data_out[16] la_data_out[15] la_data_out[14]
+ la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7]
+ la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1] la_data_out[0] io_in[26]
+ io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19] io_in[18] io_in[17] io_in[16] io_in[15]
+ io_in[14] io_in[13] io_in[12] io_in[11] io_in[10] io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4]
+ io_in[3] io_in[2] io_in[1] io_in[0] io_in_3v3[26] io_in_3v3[25] io_in_3v3[24] io_in_3v3[23] io_in_3v3[22]
+ io_in_3v3[21] io_in_3v3[20] io_in_3v3[19] io_in_3v3[18] io_in_3v3[17] io_in_3v3[16] io_in_3v3[15] io_in_3v3[14]
+ io_in_3v3[13] io_in_3v3[12] io_in_3v3[11] io_in_3v3[10] io_in_3v3[9] io_in_3v3[8] io_in_3v3[7] io_in_3v3[6]
+ io_in_3v3[5] io_in_3v3[4] io_in_3v3[3] io_in_3v3[2] io_in_3v3[1] io_in_3v3[0] user_clock2 io_out[26] io_out[25]
+ io_out[24] io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15]
+ io_out[14] io_out[13] io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7] io_out[6] io_out[5]
+ io_out[4] io_out[3] io_out[2] io_out[1] io_out[0] io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22]
+ io_oeb[21] io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12]
+ io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2]
+ io_oeb[1] io_oeb[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14] gpio_analog[13]
+ gpio_analog[12] gpio_analog[11] gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7] gpio_analog[6]
+ gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2] gpio_analog[1] gpio_analog[0] gpio_noesd[17]
+ gpio_noesd[16] gpio_noesd[15] gpio_noesd[14] gpio_noesd[13] gpio_noesd[12] gpio_noesd[11] gpio_noesd[10]
+ gpio_noesd[9] gpio_noesd[8] gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2]
+ gpio_noesd[1] gpio_noesd[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7] io_analog[6] io_analog[5]
+ io_analog[4] io_analog[3] io_analog[2] io_analog[1] io_analog[0] io_clamp_high[2] io_clamp_high[1]
+ io_clamp_high[0] io_clamp_low[2] io_clamp_low[1] io_clamp_low[0] user_irq[2] user_irq[1] user_irq[0] la_oenb[127]
+ la_oenb[126] la_oenb[125] la_oenb[124] la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119]
+ la_oenb[118] la_oenb[117] la_oenb[116] la_oenb[115] la_oenb[114] la_oenb[113] la_oenb[112] la_oenb[111]
+ la_oenb[110] la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104] la_oenb[103]
+ la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97] la_oenb[96] la_oenb[95] la_oenb[94]
+ la_oenb[93] la_oenb[92] la_oenb[91] la_oenb[90] la_oenb[89] la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85]
+ la_oenb[84] la_oenb[83] la_oenb[82] la_oenb[81] la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76]
+ la_oenb[75] la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70] la_oenb[69] la_oenb[68] la_oenb[67]
+ la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62] la_oenb[61] la_oenb[60] la_oenb[59] la_oenb[58]
+ la_oenb[57] la_oenb[56] la_oenb[55] la_oenb[54] la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49]
+ la_oenb[48] la_oenb[47] la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41] la_oenb[40]
+ la_oenb[39] la_oenb[38] la_oenb[37] la_oenb[36] la_oenb[35] la_oenb[34] la_oenb[33] la_oenb[32] la_oenb[31]
+ la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27] la_oenb[26] la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22]
+ la_oenb[21] la_oenb[20] la_oenb[19] la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15] la_oenb[14] la_oenb[13]
+ la_oenb[12] la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6] la_oenb[5] la_oenb[4]
+ la_oenb[3] la_oenb[2] la_oenb[1] la_oenb[0]
*.PININFO vdda1:B vdda2:B vssa1:B vssa2:B vccd1:B vccd2:B vssd1:B vssd2:B wb_clk_i:I wb_rst_i:I
*+ wbs_stb_i:I wbs_cyc_i:I wbs_we_i:I wbs_sel_i[3:0]:I wbs_dat_i[31:0]:I wbs_adr_i[31:0]:I wbs_ack_o:O
*+ wbs_dat_o[31:0]:O la_data_in[127:0]:I la_data_out[127:0]:O io_in[26:0]:I io_in_3v3[26:0]:I user_clock2:I
*+ io_out[26:0]:O io_oeb[26:0]:O gpio_analog[17:0]:B gpio_noesd[17:0]:B io_analog[10:0]:B io_clamp_high[2:0]:B
*+ io_clamp_low[2:0]:B user_irq[2:0]:O la_oenb[127:0]:I
x1 io_analog[0] vssa1 io_analog[4] io_analog[3] gpio_noesd[5] gpio_noesd[6] gpio_noesd[4]
+ io_analog[5] io_analog[1] io_analog[2] ina_top
.ends

* expanding   symbol:  INA_layout_v2/ina_top.sym # of pins=10
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/ina_top.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/ina_top.sch
.subckt ina_top AVDD AVSS VI_1A VI_1B VO2 VO1 VCM IREF VI_2A VI_2B
*.PININFO IREF:B VI_1A:B VI_1B:B VI_2A:B VI_2B:B VO2:B VO1:B VCM:B AVDD:B AVSS:B
x1 AVDD AVSS VI_1A VI_1B VO2 VO1 VCM VB1 VB2 VB3 VB4 VI_2A VI_2B dda
x2 IREF VB1 AVDD AVSS VB2 VB3 VB4 bias
D3 AVSS VI_2A sky130_fd_pr__diode_pw2nd_05v5 area=0.2025e12 pj=1.8e6
D4 AVSS VI_2B sky130_fd_pr__diode_pw2nd_05v5 area=0.2025e12 pj=1.8e6
D5 AVSS VI_1B sky130_fd_pr__diode_pw2nd_05v5 area=0.2025e12 pj=1.8e6
D6 AVSS VI_1A sky130_fd_pr__diode_pw2nd_05v5 area=0.2025e12 pj=1.8e6
D7 AVSS IREF sky130_fd_pr__diode_pw2nd_05v5 area=0.2025e12 pj=1.8e6
D2 AVSS VO1 sky130_fd_pr__diode_pw2nd_05v5 area=0.2025e12 pj=1.8e6
D1 AVSS VO2 sky130_fd_pr__diode_pw2nd_05v5 area=0.2025e12 pj=1.8e6
D8 AVSS VCM sky130_fd_pr__diode_pw2nd_05v5 area=0.2025e12 pj=1.8e6
.ends


* expanding   symbol:  INA_layout_v2/dda.sym # of pins=13
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/dda.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/dda.sch
.subckt dda AVDD AVSS VI_1A VI_1B VO2 VO1 VCM VB1 VB2 VB3 VB4 VI_2A VI_2B
*.PININFO AVDD:B VI_1A:B VI_1B:B VI_2A:B VI_2B:B VO1:B VO2:B VB1:B VB2:B VB3:B VB4:B VCM:B AVSS:B
x1 AVDD AVDD VB1 AVDD VB1 VIT_P2 VIT_P1 pfets_8x
x2 VIT_P1 VIT_P1 VI_1B AVDD VI_1A SUM_N SUM_P pfets_4x
x3 VIT_P2 VIT_P2 VI_2B AVDD VI_2A SUM_P SUM_N pfets_4x
x6 VD5 VD6 VB4 AVDD VB4 VO2 VO1 pfets_4x
x7 AVDD AVDD VCMFB AVDD VCMFB VD6 VD5 pfets_4x
x9 AVDD AVDD VD2 AVDD VD1 VD2 VD1 pfets_4x
x5 VO1 VO2 VB3 VB3 AVSS SUM_N SUM_P nfets_2x
x10 VD1 VCMFB VCM VO1 AVSS VIT_N1 VIT_N1 nfets_2x
x11 VD2 VCMFB VCM VO2 AVSS VIT_N2 VIT_N2 nfets_2x
x12 VIT_N1 VIT_N2 VB2 VB2 AVSS AVSS AVSS nfets_4x
x4 SUM_P SUM_N VB2 VB2 AVSS AVSS AVSS nfets_4x
x8 AVDD AVDD VCMFB AVDD VCMFB VCMFB VCMFB pfets_4x
.ends


* expanding   symbol:  INA_layout_v2/bias/bias.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/bias.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/bias.sch
.subckt bias IREF VB1 AVDD AVSS VB2 VB3 VB4
*.PININFO IREF:B VB1:B VB2:B VB3:B VB4:B AVDD:B AVSS:B
x1 IREF VB2 VB1 VB4 AVSS nbias_vb124
x2 VB3 VB1 VB2 AVDD pbias_vb123
x4 AVDD VB4 pbias_vb4
x3 VB3 AVSS nbias_vb3
.ends


* expanding   symbol:  INA_layout_v2/pfets_8x.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets_8x.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets_8x.sch
.subckt pfets_8x VS1 VS2 VG2 VB VG1 VD2 VD1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
x1[2] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets_4x
x1[1] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets_4x
.ends


* expanding   symbol:  INA_layout_v2/pfets_4x.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets_4x.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets_4x.sch
.subckt pfets_4x VS1 VS2 VG2 VB VG1 VD2 VD1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
x1[4] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets
x1[3] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets
x1[2] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets
x1[1] VS1 VS2 VG2 VB VG1 VD2 VD1 pfets
.ends


* expanding   symbol:  INA_layout_v2/nfets_2x.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets_2x.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets_2x.sch
.subckt nfets_2x VD1 VD2 VG2 VG1 VB VS2 VS1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
XM3[1] VB VB VB VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=9
XM3[0] VB VB VB VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=9
x1[2] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets
x1[1] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets
.ends


* expanding   symbol:  INA_layout_v2/nfets_4x.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets_4x.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets_4x.sch
.subckt nfets_4x VD1 VD2 VG2 VG1 VB VS2 VS1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
x1[2] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets_2x
x1[1] VD1 VD2 VG2 VG1 VB VS2 VS1 nfets_2x
.ends


* expanding   symbol:  INA_layout_v2/bias/nbias_vb124.sym # of pins=5
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nbias_vb124.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nbias_vb124.sch
.subckt nbias_vb124 IREF VB2 VB1 VB4 AVSS
*.PININFO IREF:B VB1:B VB2:B VB4:B AVSS:B
x1[5] AVSS AVSS IREF IREF nfet_2series
x1[4] AVSS AVSS IREF IREF nfet_2series
x1[3] AVSS AVSS IREF IREF nfet_2series
x1[2] AVSS AVSS IREF IREF nfet_2series
x1[1] AVSS AVSS IREF IREF nfet_2series
x2[5] AVSS AVSS IREF VB1 nfet_2series
x2[4] AVSS AVSS IREF VB1 nfet_2series
x2[3] AVSS AVSS IREF VB1 nfet_2series
x2[2] AVSS AVSS IREF VB1 nfet_2series
x2[1] AVSS AVSS IREF VB1 nfet_2series
x3[5] AVSS AVSS VB2 VB2 nfet_2series
x3[4] AVSS AVSS VB2 VB2 nfet_2series
x3[3] AVSS AVSS VB2 VB2 nfet_2series
x3[2] AVSS AVSS VB2 VB2 nfet_2series
x3[1] AVSS AVSS VB2 VB2 nfet_2series
x4[5] AVSS AVSS VB2 VB4 nfet_2series
x4[4] AVSS AVSS VB2 VB4 nfet_2series
x4[3] AVSS AVSS VB2 VB4 nfet_2series
x4[2] AVSS AVSS VB2 VB4 nfet_2series
x4[1] AVSS AVSS VB2 VB4 nfet_2series
XM1 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=44
.ends


* expanding   symbol:  INA_layout_v2/bias/pbias_vb123.sym # of pins=4
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pbias_vb123.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pbias_vb123.sch
.subckt pbias_vb123 VB3 VB1 VB2 AVDD
*.PININFO VB1:B VB2:B VB3:B AVDD:B
x1[35] AVDD AVDD VB1 VB1 pfet_2series
x1[34] AVDD AVDD VB1 VB1 pfet_2series
x1[33] AVDD AVDD VB1 VB1 pfet_2series
x1[32] AVDD AVDD VB1 VB1 pfet_2series
x1[31] AVDD AVDD VB1 VB1 pfet_2series
x1[30] AVDD AVDD VB1 VB1 pfet_2series
x1[29] AVDD AVDD VB1 VB1 pfet_2series
x1[28] AVDD AVDD VB1 VB1 pfet_2series
x1[27] AVDD AVDD VB1 VB1 pfet_2series
x1[26] AVDD AVDD VB1 VB1 pfet_2series
x1[25] AVDD AVDD VB1 VB1 pfet_2series
x1[24] AVDD AVDD VB1 VB1 pfet_2series
x1[23] AVDD AVDD VB1 VB1 pfet_2series
x1[22] AVDD AVDD VB1 VB1 pfet_2series
x1[21] AVDD AVDD VB1 VB1 pfet_2series
x1[20] AVDD AVDD VB1 VB1 pfet_2series
x1[19] AVDD AVDD VB1 VB1 pfet_2series
x1[18] AVDD AVDD VB1 VB1 pfet_2series
x1[17] AVDD AVDD VB1 VB1 pfet_2series
x1[16] AVDD AVDD VB1 VB1 pfet_2series
x1[15] AVDD AVDD VB1 VB1 pfet_2series
x1[14] AVDD AVDD VB1 VB1 pfet_2series
x1[13] AVDD AVDD VB1 VB1 pfet_2series
x1[12] AVDD AVDD VB1 VB1 pfet_2series
x1[11] AVDD AVDD VB1 VB1 pfet_2series
x1[10] AVDD AVDD VB1 VB1 pfet_2series
x1[9] AVDD AVDD VB1 VB1 pfet_2series
x1[8] AVDD AVDD VB1 VB1 pfet_2series
x1[7] AVDD AVDD VB1 VB1 pfet_2series
x1[6] AVDD AVDD VB1 VB1 pfet_2series
x1[5] AVDD AVDD VB1 VB1 pfet_2series
x1[4] AVDD AVDD VB1 VB1 pfet_2series
x1[3] AVDD AVDD VB1 VB1 pfet_2series
x1[2] AVDD AVDD VB1 VB1 pfet_2series
x1[1] AVDD AVDD VB1 VB1 pfet_2series
x2[35] AVDD AVDD VB1 VB3 pfet_2series
x2[34] AVDD AVDD VB1 VB3 pfet_2series
x2[33] AVDD AVDD VB1 VB3 pfet_2series
x2[32] AVDD AVDD VB1 VB3 pfet_2series
x2[31] AVDD AVDD VB1 VB3 pfet_2series
x2[30] AVDD AVDD VB1 VB3 pfet_2series
x2[29] AVDD AVDD VB1 VB3 pfet_2series
x2[28] AVDD AVDD VB1 VB3 pfet_2series
x2[27] AVDD AVDD VB1 VB3 pfet_2series
x2[26] AVDD AVDD VB1 VB3 pfet_2series
x2[25] AVDD AVDD VB1 VB3 pfet_2series
x2[24] AVDD AVDD VB1 VB3 pfet_2series
x2[23] AVDD AVDD VB1 VB3 pfet_2series
x2[22] AVDD AVDD VB1 VB3 pfet_2series
x2[21] AVDD AVDD VB1 VB3 pfet_2series
x2[20] AVDD AVDD VB1 VB3 pfet_2series
x2[19] AVDD AVDD VB1 VB3 pfet_2series
x2[18] AVDD AVDD VB1 VB3 pfet_2series
x2[17] AVDD AVDD VB1 VB3 pfet_2series
x2[16] AVDD AVDD VB1 VB3 pfet_2series
x2[15] AVDD AVDD VB1 VB3 pfet_2series
x2[14] AVDD AVDD VB1 VB3 pfet_2series
x2[13] AVDD AVDD VB1 VB3 pfet_2series
x2[12] AVDD AVDD VB1 VB3 pfet_2series
x2[11] AVDD AVDD VB1 VB3 pfet_2series
x2[10] AVDD AVDD VB1 VB3 pfet_2series
x2[9] AVDD AVDD VB1 VB3 pfet_2series
x2[8] AVDD AVDD VB1 VB3 pfet_2series
x2[7] AVDD AVDD VB1 VB3 pfet_2series
x2[6] AVDD AVDD VB1 VB3 pfet_2series
x2[5] AVDD AVDD VB1 VB3 pfet_2series
x2[4] AVDD AVDD VB1 VB3 pfet_2series
x2[3] AVDD AVDD VB1 VB3 pfet_2series
x2[2] AVDD AVDD VB1 VB3 pfet_2series
x2[1] AVDD AVDD VB1 VB3 pfet_2series
x3[35] AVDD AVDD VB1 VB2 pfet_2series
x3[34] AVDD AVDD VB1 VB2 pfet_2series
x3[33] AVDD AVDD VB1 VB2 pfet_2series
x3[32] AVDD AVDD VB1 VB2 pfet_2series
x3[31] AVDD AVDD VB1 VB2 pfet_2series
x3[30] AVDD AVDD VB1 VB2 pfet_2series
x3[29] AVDD AVDD VB1 VB2 pfet_2series
x3[28] AVDD AVDD VB1 VB2 pfet_2series
x3[27] AVDD AVDD VB1 VB2 pfet_2series
x3[26] AVDD AVDD VB1 VB2 pfet_2series
x3[25] AVDD AVDD VB1 VB2 pfet_2series
x3[24] AVDD AVDD VB1 VB2 pfet_2series
x3[23] AVDD AVDD VB1 VB2 pfet_2series
x3[22] AVDD AVDD VB1 VB2 pfet_2series
x3[21] AVDD AVDD VB1 VB2 pfet_2series
x3[20] AVDD AVDD VB1 VB2 pfet_2series
x3[19] AVDD AVDD VB1 VB2 pfet_2series
x3[18] AVDD AVDD VB1 VB2 pfet_2series
x3[17] AVDD AVDD VB1 VB2 pfet_2series
x3[16] AVDD AVDD VB1 VB2 pfet_2series
x3[15] AVDD AVDD VB1 VB2 pfet_2series
x3[14] AVDD AVDD VB1 VB2 pfet_2series
x3[13] AVDD AVDD VB1 VB2 pfet_2series
x3[12] AVDD AVDD VB1 VB2 pfet_2series
x3[11] AVDD AVDD VB1 VB2 pfet_2series
x3[10] AVDD AVDD VB1 VB2 pfet_2series
x3[9] AVDD AVDD VB1 VB2 pfet_2series
x3[8] AVDD AVDD VB1 VB2 pfet_2series
x3[7] AVDD AVDD VB1 VB2 pfet_2series
x3[6] AVDD AVDD VB1 VB2 pfet_2series
x3[5] AVDD AVDD VB1 VB2 pfet_2series
x3[4] AVDD AVDD VB1 VB2 pfet_2series
x3[3] AVDD AVDD VB1 VB2 pfet_2series
x3[2] AVDD AVDD VB1 VB2 pfet_2series
x3[1] AVDD AVDD VB1 VB2 pfet_2series
XM1 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=96
.ends


* expanding   symbol:  INA_layout_v2/bias/pbias_vb4.sym # of pins=2
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pbias_vb4.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pbias_vb4.sch
.subckt pbias_vb4 AVDD VB4
*.PININFO VB4:B AVDD:B
XM1 net1 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM2 net2 VB4 net1 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM3 VB4 VB4 net2 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM4 net3 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM5 net4 VB4 net3 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM6 VB4 VB4 net4 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM7 net5 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM8 net6 VB4 net5 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM9 VB4 VB4 net6 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM10 net7 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM11 net8 VB4 net7 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM12 VB4 VB4 net8 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM13 net9 VB4 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM14 net10 VB4 net9 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM15 VB4 VB4 net10 AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[20] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[19] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[18] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[17] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[16] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[15] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[14] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[13] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[12] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[11] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[10] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[9] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[8] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[7] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[6] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[5] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[4] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[3] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[2] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM16[1] AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  INA_layout_v2/bias/nbias_vb3.sym # of pins=2
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nbias_vb3.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nbias_vb3.sch
.subckt nbias_vb3 VB3 AVSS
*.PININFO AVSS:B VB3:B
x1 AVSS AVSS VB3 net1 nfet_2series
x2 net1 AVSS VB3 VB3 nfet_2series
XM1[14] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[13] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[12] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[11] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[10] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[9] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[8] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[7] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[6] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[5] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[4] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[3] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[2] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM1[1] AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  INA_layout_v2/pfets.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/pfets.sch
.subckt pfets VS1 VS2 VG2 VB VG1 VD2 VD1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
XM1 VD1 VG1 VS1 VB sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=22
XM2 VD2 VG2 VS2 VB sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=22
XM3 VB VB VB VB sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=34
.ends


* expanding   symbol:  INA_layout_v2/nfets.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/nfets.sch
.subckt nfets VD1 VD2 VG2 VG1 VB VS2 VS1
*.PININFO VS1:B VS2:B VB:B VG1:B VG2:B VD1:B VD2:B
XM1 VD1 VG1 VS1 VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=7
XM2 VD2 VG2 VS2 VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=7
XM3 VB VB VB VB sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=4
.ends


* expanding   symbol:  INA_layout_v2/bias/nfet_2series.sym # of pins=4
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nfet_2series.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/nfet_2series.sch
.subckt nfet_2series S B G D
*.PININFO S:B B:B G:B D:B
XM1 D G net1 B sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM2 net1 G S B sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  INA_layout_v2/bias/pfet_2series.sym # of pins=4
** sym_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pfet_2series.sym
** sch_path: /home/gmaranhao/Desktop/sky130_work/INA_layout_v2/bias/pfet_2series.sch
.subckt pfet_2series S B G D
*.PININFO S:B B:B G:B D:B
XM1 net1 G S B sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
XM2 D G net1 B sky130_fd_pr__pfet_01v8_hvt L=1 W=1 nf=1 m=1
.ends

.end
