* NGSPICE file created from pbias_vb123.ext - technology: sky130A

.subckt pbias_vb123 VB3 VB2 AVDD VB1
X0 VB3 VB1 a_3228_3476# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 a_2712_1968# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X3 a_5228_2589# VB1 a_4970_2589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X4 a_1486_599# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X5 a_4002_4980# VB1 a_3744_4980# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X6 a_3228_599# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X7 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X8 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X9 a_2712_4093# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X10 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X11 a_4970_1968# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X12 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X13 a_3228_n962# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 a_3744_4980# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X15 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X16 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X17 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X18 a_2002_n495# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X20 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X21 a_2260_n3972# VB1 a_2002_n3972# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X22 a_5228_n3085# VB1 a_4970_n3085# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X23 VB2 VB1 a_3228_n3085# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X24 a_4970_n2468# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X25 VB3 VB1 a_3228_4980# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 a_4002_599# VB1 a_3744_599# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X27 VB1 VB1 a_1486_n495# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X28 a_4970_4093# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 a_4454_134# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X30 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X31 a_5228_1968# VB1 a_4970_1968# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X32 a_1486_n495# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X33 a_4002_n2468# VB1 a_3744_n2468# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X34 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X35 VB2 VB1 a_4454_n2468# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X36 AVDD VB1 a_2712_n2468# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 a_3228_n3085# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X38 a_1486_n3085# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X39 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X40 a_2002_3476# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X41 a_2260_2589# VB1 a_2002_2589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X42 AVDD VB1 a_2712_2589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X43 a_4002_1220# VB1 a_3744_1220# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X44 a_3744_n4589# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X45 a_4970_n3972# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X46 a_2002_n2468# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X47 a_5228_4093# VB1 a_4970_4093# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X48 a_4454_n4589# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X49 a_2712_n2468# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X50 VB2 VB1 a_1486_3476# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X51 a_3744_1220# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X52 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X53 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X54 VB1 VB1 a_1486_134# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X55 a_4002_n3972# VB1 a_3744_n3972# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X56 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X57 a_1486_3476# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X58 VB1 VB1 a_3228_1220# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X59 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X60 VB2 VB1 a_4454_n3972# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X61 AVDD VB1 a_2712_n3972# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X62 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X63 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X64 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X65 VB3 VB1 a_1486_n4589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X66 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X67 a_3228_2589# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X68 a_2260_134# VB1 a_2002_134# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X69 a_2002_4980# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X70 VB1 VB1 a_4454_n495# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X71 a_2260_1968# VB1 a_2002_1968# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X72 AVDD VB1 a_2712_1968# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X73 a_2002_n3972# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X74 a_2712_n3972# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X75 VB2 VB1 a_1486_4980# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X76 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X77 a_4454_n495# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X78 a_4002_n962# VB1 a_3744_n962# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X79 VB2 VB1 a_3228_n1581# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X80 a_5228_n1581# VB1 a_4970_n1581# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X81 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X82 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X83 a_1486_4980# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X84 a_3744_n962# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X85 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X86 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X87 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X88 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X89 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X90 a_2260_4093# VB1 a_2002_4093# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X91 AVDD VB1 a_2712_4093# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X92 VB1 VB1 a_3228_n962# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X93 a_3228_n1581# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X94 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X95 a_3228_1968# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X96 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X97 a_1486_n1581# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X98 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X99 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X100 VB2 VB1 a_4454_3476# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X101 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X102 a_4454_3476# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X103 a_3744_599# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X104 a_2002_1220# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X105 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X106 a_3228_4093# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X107 a_2260_n4589# VB1 a_2002_n4589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X108 VB1 VB1 a_1486_1220# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X109 a_2712_134# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X110 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X111 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X112 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X113 a_1486_1220# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X114 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X115 a_3744_n3085# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X116 VB2 VB1 a_4454_4980# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X117 a_4970_134# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X118 a_4454_n3085# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X119 a_4454_4980# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X120 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X121 a_4002_2589# VB1 a_3744_2589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X122 a_2712_n495# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X123 a_1486_134# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X124 a_3228_134# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X125 a_4970_n4589# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X126 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X127 VB3 VB1 a_1486_n3085# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X128 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X129 a_3744_2589# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X130 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X131 a_2002_n962# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X132 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X133 VB2 VB1 a_3228_2589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X134 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X135 VB1 VB1 a_1486_n962# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X136 a_4002_n4589# VB1 a_3744_n4589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X137 a_4970_n495# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X138 VB3 VB1 a_4454_n4589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X139 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X140 a_4002_134# VB1 a_3744_134# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X141 a_1486_n962# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X142 AVDD VB1 a_2712_n4589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X143 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X144 a_4002_1968# VB1 a_3744_1968# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X145 AVDD VB1 a_2712_599# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X146 a_2712_3476# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X147 VB1 VB1 a_4454_1220# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X148 VB1 VB1 a_4454_599# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X149 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X150 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X151 a_3744_1968# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X152 a_2002_n4589# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X153 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X154 a_2712_n4589# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X155 a_5228_n2468# VB1 a_4970_n2468# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X156 a_4454_1220# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X157 a_5228_n495# VB1 a_4970_n495# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X158 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X159 VB3 VB1 a_3228_n2468# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X160 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X161 VB3 VB1 a_3228_1968# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X162 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X163 a_4002_4093# VB1 a_3744_4093# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X164 a_4970_3476# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X165 a_3744_n1581# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X166 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X167 a_3744_4093# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X168 VB1 VB1 a_3228_599# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X169 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X170 a_3228_n2468# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X171 a_4454_n1581# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X172 a_5228_599# VB1 a_4970_599# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X173 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X174 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X175 a_2260_n3085# VB1 a_2002_n3085# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X176 a_1486_n2468# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X177 a_2712_4980# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X178 VB2 VB1 a_3228_4093# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X179 a_2002_599# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X180 a_2002_2589# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X181 VB1 VB1 a_4454_n962# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X182 a_5228_n3972# VB1 a_4970_n3972# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X183 a_5228_3476# VB1 a_4970_3476# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X184 VB3 VB1 a_1486_n1581# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X185 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X186 VB3 VB1 a_3228_n3972# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X187 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X188 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X189 VB3 VB1 a_1486_2589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X190 a_4454_n962# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X191 a_4970_4980# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X192 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X193 a_1486_2589# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X194 a_3228_n3972# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X195 a_1486_n3972# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X196 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X197 a_2260_n495# VB1 a_2002_n495# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X198 AVDD VB1 a_2712_n495# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X199 a_4970_n3085# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X200 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X201 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X202 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X203 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X204 a_2002_1968# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X205 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X206 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X207 a_5228_4980# VB1 a_4970_4980# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X208 a_2712_1220# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X209 a_4002_n3085# VB1 a_3744_n3085# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X210 VB3 VB1 a_4454_n3085# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X211 VB2 VB1 a_1486_1968# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X212 AVDD VB1 a_2712_n3085# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X213 a_1486_1968# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X214 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X215 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X216 a_3744_134# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X217 a_3228_n495# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X218 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X219 a_2002_4093# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X220 a_2260_3476# VB1 a_2002_3476# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X221 AVDD VB1 a_2712_3476# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X222 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X223 a_2002_n3085# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X224 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X225 a_4970_1220# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X226 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X227 a_4454_599# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X228 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X229 a_2712_n3085# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X230 VB3 VB1 a_1486_4093# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X231 a_2260_n1581# VB1 a_2002_n1581# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X232 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X233 VB3 VB1 a_4454_2589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X234 a_1486_4093# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X235 a_4454_2589# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X236 a_2712_n962# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X237 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X238 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X239 a_3228_3476# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X240 a_5228_1220# VB1 a_4970_1220# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X241 a_2260_4980# VB1 a_2002_4980# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X242 AVDD VB1 a_2712_4980# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X243 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X244 VB1 VB1 a_1486_599# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X245 a_3744_n2468# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X246 a_4970_n1581# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X247 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X248 VB2 VB1 a_4454_1968# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X249 a_4970_n962# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X250 a_4454_n2468# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X251 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X252 a_2260_599# VB1 a_2002_599# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X253 a_4454_1968# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X254 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X255 a_4002_n1581# VB1 a_3744_n1581# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X256 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X257 VB3 VB1 a_4454_n1581# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X258 a_3228_4980# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X259 AVDD VB1 a_2712_n1581# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X260 a_5228_n4589# VB1 a_4970_n4589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X261 VB2 VB1 a_3228_n4589# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X262 VB2 VB1 a_1486_n2468# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X263 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X264 AVDD VB1 a_2712_134# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X265 VB1 VB1 a_4454_134# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X266 VB3 VB1 a_4454_4093# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X267 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X268 a_5228_n962# VB1 a_4970_n962# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X269 a_4454_4093# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X270 a_4002_n495# VB1 a_3744_n495# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X271 a_2002_n1581# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X272 a_3744_n3972# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X273 a_2712_n1581# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X274 a_3228_n4589# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X275 a_4454_n3972# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X276 a_2260_1220# VB1 a_2002_1220# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X277 AVDD VB1 a_2712_1220# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X278 a_3744_n495# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X279 a_1486_n4589# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X280 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X281 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X282 a_2712_2589# VB1 VB2 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X283 VB1 VB1 a_3228_134# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X284 VB1 VB1 a_3228_n495# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X285 a_5228_134# VB1 a_4970_134# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X286 VB2 VB1 a_1486_n3972# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X287 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X288 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X289 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X290 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X291 a_3228_1220# VB1 AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X292 a_2002_134# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X293 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X294 a_4002_3476# VB1 a_3744_3476# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X295 a_4970_2589# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X296 a_2712_599# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X297 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X298 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X299 a_3744_3476# VB1 VB3 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X300 a_4970_599# VB1 VB1 AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X301 a_2260_n962# VB1 a_2002_n962# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X302 AVDD VB1 a_2712_n962# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X303 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X304 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X305 a_2260_n2468# VB1 a_2002_n2468# AVDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
.ends

