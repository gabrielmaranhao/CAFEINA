magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< pwell >>
rect -2484 2078 3567 2164
rect -2484 -1755 -2398 2078
rect 3481 -1755 3567 2078
rect -2484 -1841 3567 -1755
<< psubdiff >>
rect -2458 2104 -2273 2138
rect -2239 2104 -2205 2138
rect -2171 2104 -2137 2138
rect -2103 2104 -2069 2138
rect -2035 2104 -2001 2138
rect -1967 2104 -1933 2138
rect -1899 2104 -1865 2138
rect -1831 2104 -1797 2138
rect -1763 2104 -1729 2138
rect -1695 2104 -1661 2138
rect -1627 2104 -1593 2138
rect -1559 2104 -1525 2138
rect -1491 2104 -1457 2138
rect -1423 2104 -1389 2138
rect -1355 2104 -1321 2138
rect -1287 2104 -1253 2138
rect -1219 2104 -1185 2138
rect -1151 2104 -1117 2138
rect -1083 2104 -1049 2138
rect -1015 2104 -981 2138
rect -947 2104 -913 2138
rect -879 2104 -845 2138
rect -811 2104 -777 2138
rect -743 2104 -709 2138
rect -675 2104 -641 2138
rect -607 2104 -573 2138
rect -539 2104 -505 2138
rect -471 2104 -437 2138
rect -403 2104 -369 2138
rect -335 2104 -301 2138
rect -267 2104 -233 2138
rect -199 2104 -165 2138
rect -131 2104 -97 2138
rect -63 2104 -29 2138
rect 5 2104 39 2138
rect 73 2104 107 2138
rect 141 2104 175 2138
rect 209 2104 243 2138
rect 277 2104 311 2138
rect 345 2104 379 2138
rect 413 2104 447 2138
rect 481 2104 515 2138
rect 549 2104 583 2138
rect 617 2104 651 2138
rect 685 2104 719 2138
rect 753 2104 787 2138
rect 821 2104 855 2138
rect 889 2104 923 2138
rect 957 2104 991 2138
rect 1025 2104 1059 2138
rect 1093 2104 1127 2138
rect 1161 2104 1195 2138
rect 1229 2104 1263 2138
rect 1297 2104 1331 2138
rect 1365 2104 1399 2138
rect 1433 2104 1467 2138
rect 1501 2104 1535 2138
rect 1569 2104 1603 2138
rect 1637 2104 1671 2138
rect 1705 2104 1739 2138
rect 1773 2104 1807 2138
rect 1841 2104 1875 2138
rect 1909 2104 1943 2138
rect 1977 2104 2011 2138
rect 2045 2104 2079 2138
rect 2113 2104 2147 2138
rect 2181 2104 2215 2138
rect 2249 2104 2283 2138
rect 2317 2104 2351 2138
rect 2385 2104 2419 2138
rect 2453 2104 2487 2138
rect 2521 2104 2555 2138
rect 2589 2104 2623 2138
rect 2657 2104 2691 2138
rect 2725 2104 2759 2138
rect 2793 2104 2827 2138
rect 2861 2104 2895 2138
rect 2929 2104 2963 2138
rect 2997 2104 3031 2138
rect 3065 2104 3099 2138
rect 3133 2104 3167 2138
rect 3201 2104 3235 2138
rect 3269 2104 3303 2138
rect 3337 2104 3541 2138
rect -2458 1953 -2424 2104
rect -2458 1885 -2424 1919
rect -2458 1817 -2424 1851
rect -2458 1749 -2424 1783
rect -2458 1681 -2424 1715
rect -2458 1613 -2424 1647
rect -2458 1545 -2424 1579
rect -2458 1477 -2424 1511
rect -2458 1409 -2424 1443
rect -2458 1341 -2424 1375
rect -2458 1273 -2424 1307
rect -2458 1205 -2424 1239
rect -2458 1137 -2424 1171
rect -2458 1069 -2424 1103
rect -2458 1001 -2424 1035
rect -2458 933 -2424 967
rect -2458 865 -2424 899
rect -2458 797 -2424 831
rect -2458 729 -2424 763
rect -2458 661 -2424 695
rect -2458 593 -2424 627
rect -2458 525 -2424 559
rect -2458 457 -2424 491
rect -2458 389 -2424 423
rect -2458 321 -2424 355
rect -2458 253 -2424 287
rect -2458 185 -2424 219
rect -2458 117 -2424 151
rect -2458 49 -2424 83
rect -2458 -19 -2424 15
rect -2458 -87 -2424 -53
rect -2458 -155 -2424 -121
rect -2458 -223 -2424 -189
rect -2458 -291 -2424 -257
rect -2458 -359 -2424 -325
rect -2458 -427 -2424 -393
rect -2458 -495 -2424 -461
rect -2458 -563 -2424 -529
rect -2458 -631 -2424 -597
rect -2458 -699 -2424 -665
rect -2458 -767 -2424 -733
rect -2458 -835 -2424 -801
rect -2458 -903 -2424 -869
rect -2458 -971 -2424 -937
rect -2458 -1039 -2424 -1005
rect -2458 -1107 -2424 -1073
rect -2458 -1175 -2424 -1141
rect -2458 -1243 -2424 -1209
rect -2458 -1311 -2424 -1277
rect -2458 -1379 -2424 -1345
rect -2458 -1447 -2424 -1413
rect -2458 -1515 -2424 -1481
rect -2458 -1583 -2424 -1549
rect -2458 -1781 -2424 -1617
rect 3507 1953 3541 2104
rect 3507 1885 3541 1919
rect 3507 1817 3541 1851
rect 3507 1749 3541 1783
rect 3507 1681 3541 1715
rect 3507 1613 3541 1647
rect 3507 1545 3541 1579
rect 3507 1477 3541 1511
rect 3507 1409 3541 1443
rect 3507 1341 3541 1375
rect 3507 1273 3541 1307
rect 3507 1205 3541 1239
rect 3507 1137 3541 1171
rect 3507 1069 3541 1103
rect 3507 1001 3541 1035
rect 3507 933 3541 967
rect 3507 865 3541 899
rect 3507 797 3541 831
rect 3507 729 3541 763
rect 3507 661 3541 695
rect 3507 593 3541 627
rect 3507 525 3541 559
rect 3507 457 3541 491
rect 3507 389 3541 423
rect 3507 321 3541 355
rect 3507 253 3541 287
rect 3507 185 3541 219
rect 3507 117 3541 151
rect 3507 49 3541 83
rect 3507 -19 3541 15
rect 3507 -87 3541 -53
rect 3507 -155 3541 -121
rect 3507 -223 3541 -189
rect 3507 -291 3541 -257
rect 3507 -359 3541 -325
rect 3507 -427 3541 -393
rect 3507 -495 3541 -461
rect 3507 -563 3541 -529
rect 3507 -631 3541 -597
rect 3507 -699 3541 -665
rect 3507 -767 3541 -733
rect 3507 -835 3541 -801
rect 3507 -903 3541 -869
rect 3507 -971 3541 -937
rect 3507 -1039 3541 -1005
rect 3507 -1107 3541 -1073
rect 3507 -1175 3541 -1141
rect 3507 -1243 3541 -1209
rect 3507 -1781 3541 -1277
rect -2458 -1815 -2273 -1781
rect -2239 -1815 -2205 -1781
rect -2171 -1815 -2137 -1781
rect -2103 -1815 -2069 -1781
rect -2035 -1815 -2001 -1781
rect -1967 -1815 -1933 -1781
rect -1899 -1815 -1865 -1781
rect -1831 -1815 -1797 -1781
rect -1763 -1815 -1729 -1781
rect -1695 -1815 -1661 -1781
rect -1627 -1815 -1593 -1781
rect -1559 -1815 -1525 -1781
rect -1491 -1815 -1457 -1781
rect -1423 -1815 -1389 -1781
rect -1355 -1815 -1321 -1781
rect -1287 -1815 -1253 -1781
rect -1219 -1815 -1185 -1781
rect -1151 -1815 -1117 -1781
rect -1083 -1815 -1049 -1781
rect -1015 -1815 -981 -1781
rect -947 -1815 -913 -1781
rect -879 -1815 -845 -1781
rect -811 -1815 -777 -1781
rect -743 -1815 -709 -1781
rect -675 -1815 -641 -1781
rect -607 -1815 -573 -1781
rect -539 -1815 -505 -1781
rect -471 -1815 -437 -1781
rect -403 -1815 -369 -1781
rect -335 -1815 -301 -1781
rect -267 -1815 -233 -1781
rect -199 -1815 -165 -1781
rect -131 -1815 -97 -1781
rect -63 -1815 -29 -1781
rect 5 -1815 39 -1781
rect 73 -1815 107 -1781
rect 141 -1815 175 -1781
rect 209 -1815 243 -1781
rect 277 -1815 311 -1781
rect 345 -1815 379 -1781
rect 413 -1815 447 -1781
rect 481 -1815 515 -1781
rect 549 -1815 583 -1781
rect 617 -1815 651 -1781
rect 685 -1815 719 -1781
rect 753 -1815 787 -1781
rect 821 -1815 855 -1781
rect 889 -1815 923 -1781
rect 957 -1815 991 -1781
rect 1025 -1815 1059 -1781
rect 1093 -1815 1127 -1781
rect 1161 -1815 1195 -1781
rect 1229 -1815 1263 -1781
rect 1297 -1815 1331 -1781
rect 1365 -1815 1399 -1781
rect 1433 -1815 1467 -1781
rect 1501 -1815 1535 -1781
rect 1569 -1815 1603 -1781
rect 1637 -1815 1671 -1781
rect 1705 -1815 1739 -1781
rect 1773 -1815 1807 -1781
rect 1841 -1815 1875 -1781
rect 1909 -1815 1943 -1781
rect 1977 -1815 2011 -1781
rect 2045 -1815 2079 -1781
rect 2113 -1815 2147 -1781
rect 2181 -1815 2215 -1781
rect 2249 -1815 2283 -1781
rect 2317 -1815 2351 -1781
rect 2385 -1815 2419 -1781
rect 2453 -1815 2487 -1781
rect 2521 -1815 2555 -1781
rect 2589 -1815 2623 -1781
rect 2657 -1815 2691 -1781
rect 2725 -1815 2759 -1781
rect 2793 -1815 2827 -1781
rect 2861 -1815 2895 -1781
rect 2929 -1815 2963 -1781
rect 2997 -1815 3031 -1781
rect 3065 -1815 3099 -1781
rect 3133 -1815 3167 -1781
rect 3201 -1815 3235 -1781
rect 3269 -1815 3303 -1781
rect 3337 -1815 3541 -1781
<< psubdiffcont >>
rect -2273 2104 -2239 2138
rect -2205 2104 -2171 2138
rect -2137 2104 -2103 2138
rect -2069 2104 -2035 2138
rect -2001 2104 -1967 2138
rect -1933 2104 -1899 2138
rect -1865 2104 -1831 2138
rect -1797 2104 -1763 2138
rect -1729 2104 -1695 2138
rect -1661 2104 -1627 2138
rect -1593 2104 -1559 2138
rect -1525 2104 -1491 2138
rect -1457 2104 -1423 2138
rect -1389 2104 -1355 2138
rect -1321 2104 -1287 2138
rect -1253 2104 -1219 2138
rect -1185 2104 -1151 2138
rect -1117 2104 -1083 2138
rect -1049 2104 -1015 2138
rect -981 2104 -947 2138
rect -913 2104 -879 2138
rect -845 2104 -811 2138
rect -777 2104 -743 2138
rect -709 2104 -675 2138
rect -641 2104 -607 2138
rect -573 2104 -539 2138
rect -505 2104 -471 2138
rect -437 2104 -403 2138
rect -369 2104 -335 2138
rect -301 2104 -267 2138
rect -233 2104 -199 2138
rect -165 2104 -131 2138
rect -97 2104 -63 2138
rect -29 2104 5 2138
rect 39 2104 73 2138
rect 107 2104 141 2138
rect 175 2104 209 2138
rect 243 2104 277 2138
rect 311 2104 345 2138
rect 379 2104 413 2138
rect 447 2104 481 2138
rect 515 2104 549 2138
rect 583 2104 617 2138
rect 651 2104 685 2138
rect 719 2104 753 2138
rect 787 2104 821 2138
rect 855 2104 889 2138
rect 923 2104 957 2138
rect 991 2104 1025 2138
rect 1059 2104 1093 2138
rect 1127 2104 1161 2138
rect 1195 2104 1229 2138
rect 1263 2104 1297 2138
rect 1331 2104 1365 2138
rect 1399 2104 1433 2138
rect 1467 2104 1501 2138
rect 1535 2104 1569 2138
rect 1603 2104 1637 2138
rect 1671 2104 1705 2138
rect 1739 2104 1773 2138
rect 1807 2104 1841 2138
rect 1875 2104 1909 2138
rect 1943 2104 1977 2138
rect 2011 2104 2045 2138
rect 2079 2104 2113 2138
rect 2147 2104 2181 2138
rect 2215 2104 2249 2138
rect 2283 2104 2317 2138
rect 2351 2104 2385 2138
rect 2419 2104 2453 2138
rect 2487 2104 2521 2138
rect 2555 2104 2589 2138
rect 2623 2104 2657 2138
rect 2691 2104 2725 2138
rect 2759 2104 2793 2138
rect 2827 2104 2861 2138
rect 2895 2104 2929 2138
rect 2963 2104 2997 2138
rect 3031 2104 3065 2138
rect 3099 2104 3133 2138
rect 3167 2104 3201 2138
rect 3235 2104 3269 2138
rect 3303 2104 3337 2138
rect -2458 1919 -2424 1953
rect -2458 1851 -2424 1885
rect -2458 1783 -2424 1817
rect -2458 1715 -2424 1749
rect -2458 1647 -2424 1681
rect -2458 1579 -2424 1613
rect -2458 1511 -2424 1545
rect -2458 1443 -2424 1477
rect -2458 1375 -2424 1409
rect -2458 1307 -2424 1341
rect -2458 1239 -2424 1273
rect -2458 1171 -2424 1205
rect -2458 1103 -2424 1137
rect -2458 1035 -2424 1069
rect -2458 967 -2424 1001
rect -2458 899 -2424 933
rect -2458 831 -2424 865
rect -2458 763 -2424 797
rect -2458 695 -2424 729
rect -2458 627 -2424 661
rect -2458 559 -2424 593
rect -2458 491 -2424 525
rect -2458 423 -2424 457
rect -2458 355 -2424 389
rect -2458 287 -2424 321
rect -2458 219 -2424 253
rect -2458 151 -2424 185
rect -2458 83 -2424 117
rect -2458 15 -2424 49
rect -2458 -53 -2424 -19
rect -2458 -121 -2424 -87
rect -2458 -189 -2424 -155
rect -2458 -257 -2424 -223
rect -2458 -325 -2424 -291
rect -2458 -393 -2424 -359
rect -2458 -461 -2424 -427
rect -2458 -529 -2424 -495
rect -2458 -597 -2424 -563
rect -2458 -665 -2424 -631
rect -2458 -733 -2424 -699
rect -2458 -801 -2424 -767
rect -2458 -869 -2424 -835
rect -2458 -937 -2424 -903
rect -2458 -1005 -2424 -971
rect -2458 -1073 -2424 -1039
rect -2458 -1141 -2424 -1107
rect -2458 -1209 -2424 -1175
rect -2458 -1277 -2424 -1243
rect -2458 -1345 -2424 -1311
rect -2458 -1413 -2424 -1379
rect -2458 -1481 -2424 -1447
rect -2458 -1549 -2424 -1515
rect -2458 -1617 -2424 -1583
rect 3507 1919 3541 1953
rect 3507 1851 3541 1885
rect 3507 1783 3541 1817
rect 3507 1715 3541 1749
rect 3507 1647 3541 1681
rect 3507 1579 3541 1613
rect 3507 1511 3541 1545
rect 3507 1443 3541 1477
rect 3507 1375 3541 1409
rect 3507 1307 3541 1341
rect 3507 1239 3541 1273
rect 3507 1171 3541 1205
rect 3507 1103 3541 1137
rect 3507 1035 3541 1069
rect 3507 967 3541 1001
rect 3507 899 3541 933
rect 3507 831 3541 865
rect 3507 763 3541 797
rect 3507 695 3541 729
rect 3507 627 3541 661
rect 3507 559 3541 593
rect 3507 491 3541 525
rect 3507 423 3541 457
rect 3507 355 3541 389
rect 3507 287 3541 321
rect 3507 219 3541 253
rect 3507 151 3541 185
rect 3507 83 3541 117
rect 3507 15 3541 49
rect 3507 -53 3541 -19
rect 3507 -121 3541 -87
rect 3507 -189 3541 -155
rect 3507 -257 3541 -223
rect 3507 -325 3541 -291
rect 3507 -393 3541 -359
rect 3507 -461 3541 -427
rect 3507 -529 3541 -495
rect 3507 -597 3541 -563
rect 3507 -665 3541 -631
rect 3507 -733 3541 -699
rect 3507 -801 3541 -767
rect 3507 -869 3541 -835
rect 3507 -937 3541 -903
rect 3507 -1005 3541 -971
rect 3507 -1073 3541 -1039
rect 3507 -1141 3541 -1107
rect 3507 -1209 3541 -1175
rect 3507 -1277 3541 -1243
rect -2273 -1815 -2239 -1781
rect -2205 -1815 -2171 -1781
rect -2137 -1815 -2103 -1781
rect -2069 -1815 -2035 -1781
rect -2001 -1815 -1967 -1781
rect -1933 -1815 -1899 -1781
rect -1865 -1815 -1831 -1781
rect -1797 -1815 -1763 -1781
rect -1729 -1815 -1695 -1781
rect -1661 -1815 -1627 -1781
rect -1593 -1815 -1559 -1781
rect -1525 -1815 -1491 -1781
rect -1457 -1815 -1423 -1781
rect -1389 -1815 -1355 -1781
rect -1321 -1815 -1287 -1781
rect -1253 -1815 -1219 -1781
rect -1185 -1815 -1151 -1781
rect -1117 -1815 -1083 -1781
rect -1049 -1815 -1015 -1781
rect -981 -1815 -947 -1781
rect -913 -1815 -879 -1781
rect -845 -1815 -811 -1781
rect -777 -1815 -743 -1781
rect -709 -1815 -675 -1781
rect -641 -1815 -607 -1781
rect -573 -1815 -539 -1781
rect -505 -1815 -471 -1781
rect -437 -1815 -403 -1781
rect -369 -1815 -335 -1781
rect -301 -1815 -267 -1781
rect -233 -1815 -199 -1781
rect -165 -1815 -131 -1781
rect -97 -1815 -63 -1781
rect -29 -1815 5 -1781
rect 39 -1815 73 -1781
rect 107 -1815 141 -1781
rect 175 -1815 209 -1781
rect 243 -1815 277 -1781
rect 311 -1815 345 -1781
rect 379 -1815 413 -1781
rect 447 -1815 481 -1781
rect 515 -1815 549 -1781
rect 583 -1815 617 -1781
rect 651 -1815 685 -1781
rect 719 -1815 753 -1781
rect 787 -1815 821 -1781
rect 855 -1815 889 -1781
rect 923 -1815 957 -1781
rect 991 -1815 1025 -1781
rect 1059 -1815 1093 -1781
rect 1127 -1815 1161 -1781
rect 1195 -1815 1229 -1781
rect 1263 -1815 1297 -1781
rect 1331 -1815 1365 -1781
rect 1399 -1815 1433 -1781
rect 1467 -1815 1501 -1781
rect 1535 -1815 1569 -1781
rect 1603 -1815 1637 -1781
rect 1671 -1815 1705 -1781
rect 1739 -1815 1773 -1781
rect 1807 -1815 1841 -1781
rect 1875 -1815 1909 -1781
rect 1943 -1815 1977 -1781
rect 2011 -1815 2045 -1781
rect 2079 -1815 2113 -1781
rect 2147 -1815 2181 -1781
rect 2215 -1815 2249 -1781
rect 2283 -1815 2317 -1781
rect 2351 -1815 2385 -1781
rect 2419 -1815 2453 -1781
rect 2487 -1815 2521 -1781
rect 2555 -1815 2589 -1781
rect 2623 -1815 2657 -1781
rect 2691 -1815 2725 -1781
rect 2759 -1815 2793 -1781
rect 2827 -1815 2861 -1781
rect 2895 -1815 2929 -1781
rect 2963 -1815 2997 -1781
rect 3031 -1815 3065 -1781
rect 3099 -1815 3133 -1781
rect 3167 -1815 3201 -1781
rect 3235 -1815 3269 -1781
rect 3303 -1815 3337 -1781
<< locali >>
rect -2458 2104 -2293 2138
rect -2239 2104 -2221 2138
rect -2171 2104 -2149 2138
rect -2103 2104 -2077 2138
rect -2035 2104 -2005 2138
rect -1967 2104 -1933 2138
rect -1899 2104 -1865 2138
rect -1827 2104 -1797 2138
rect -1755 2104 -1729 2138
rect -1683 2104 -1661 2138
rect -1611 2104 -1593 2138
rect -1539 2104 -1525 2138
rect -1467 2104 -1457 2138
rect -1395 2104 -1389 2138
rect -1323 2104 -1321 2138
rect -1287 2104 -1285 2138
rect -1219 2104 -1213 2138
rect -1151 2104 -1141 2138
rect -1083 2104 -1069 2138
rect -1015 2104 -997 2138
rect -947 2104 -925 2138
rect -879 2104 -853 2138
rect -811 2104 -781 2138
rect -743 2104 -709 2138
rect -675 2104 -641 2138
rect -603 2104 -573 2138
rect -531 2104 -505 2138
rect -459 2104 -437 2138
rect -387 2104 -369 2138
rect -315 2104 -301 2138
rect -243 2104 -233 2138
rect -171 2104 -165 2138
rect -99 2104 -97 2138
rect -63 2104 -61 2138
rect 5 2104 11 2138
rect 73 2104 83 2138
rect 141 2104 155 2138
rect 209 2104 227 2138
rect 277 2104 299 2138
rect 345 2104 371 2138
rect 413 2104 443 2138
rect 481 2104 515 2138
rect 549 2104 583 2138
rect 621 2104 651 2138
rect 693 2104 719 2138
rect 765 2104 787 2138
rect 837 2104 855 2138
rect 909 2104 923 2138
rect 981 2104 991 2138
rect 1025 2104 1043 2138
rect 1093 2104 1115 2138
rect 1161 2104 1187 2138
rect 1229 2104 1259 2138
rect 1297 2104 1331 2138
rect 1365 2104 1399 2138
rect 1437 2104 1467 2138
rect 1509 2104 1535 2138
rect 1581 2104 1603 2138
rect 1653 2104 1671 2138
rect 1725 2104 1739 2138
rect 1797 2104 1807 2138
rect 1869 2104 1875 2138
rect 1941 2104 1943 2138
rect 1977 2104 1979 2138
rect 2045 2104 2051 2138
rect 2113 2104 2123 2138
rect 2181 2104 2195 2138
rect 2249 2104 2267 2138
rect 2317 2104 2339 2138
rect 2385 2104 2411 2138
rect 2453 2104 2483 2138
rect 2521 2104 2555 2138
rect 2589 2104 2623 2138
rect 2661 2104 2691 2138
rect 2733 2104 2759 2138
rect 2805 2104 2827 2138
rect 2877 2104 2895 2138
rect 2949 2104 2963 2138
rect 3021 2104 3031 2138
rect 3093 2104 3099 2138
rect 3165 2104 3167 2138
rect 3201 2104 3203 2138
rect 3269 2104 3275 2138
rect 3337 2104 3541 2138
rect -2458 1974 -2424 2104
rect -2458 1902 -2424 1919
rect -2458 1830 -2424 1851
rect -2458 1758 -2424 1783
rect -2458 1686 -2424 1715
rect -2458 1614 -2424 1647
rect -2458 1545 -2424 1579
rect -2458 1477 -2424 1508
rect -2458 1409 -2424 1436
rect -2458 1341 -2424 1364
rect -2458 1273 -2424 1292
rect -2458 1205 -2424 1220
rect -2458 1137 -2424 1148
rect -2458 1069 -2424 1076
rect -2458 1001 -2424 1004
rect -2458 966 -2424 967
rect -2458 894 -2424 899
rect -2458 822 -2424 831
rect -2458 750 -2424 763
rect -2458 678 -2424 695
rect -2458 606 -2424 627
rect -2458 534 -2424 559
rect -2458 462 -2424 491
rect -2458 390 -2424 423
rect -2458 321 -2424 355
rect -2458 253 -2424 284
rect -2458 185 -2424 212
rect -2458 117 -2424 140
rect -2458 49 -2424 68
rect -2458 -19 -2424 -4
rect -2458 -87 -2424 -76
rect -2458 -155 -2424 -148
rect -2458 -223 -2424 -220
rect -2458 -258 -2424 -257
rect -2458 -330 -2424 -325
rect -2458 -402 -2424 -393
rect -2458 -474 -2424 -461
rect -2458 -546 -2424 -529
rect -2458 -618 -2424 -597
rect -2458 -690 -2424 -665
rect -2458 -762 -2424 -733
rect -2458 -834 -2424 -801
rect -2458 -903 -2424 -869
rect -2458 -971 -2424 -940
rect -2458 -1039 -2424 -1012
rect -2458 -1107 -2424 -1084
rect -2458 -1175 -2424 -1156
rect -2458 -1243 -2424 -1228
rect -2458 -1311 -2424 -1300
rect -2458 -1379 -2424 -1372
rect -2458 -1447 -2424 -1444
rect -2458 -1482 -2424 -1481
rect -2458 -1554 -2424 -1549
rect -2458 -1626 -2424 -1617
rect -2458 -1781 -2424 -1660
rect 3507 1974 3541 2104
rect 3507 1902 3541 1919
rect 3507 1830 3541 1851
rect 3507 1758 3541 1783
rect 3507 1686 3541 1715
rect 3507 1614 3541 1647
rect 3507 1545 3541 1579
rect 3507 1477 3541 1508
rect 3507 1409 3541 1436
rect 3507 1341 3541 1364
rect 3507 1273 3541 1292
rect 3507 1205 3541 1220
rect 3507 1137 3541 1148
rect 3507 1069 3541 1076
rect 3507 1001 3541 1004
rect 3507 966 3541 967
rect 3507 894 3541 899
rect 3507 822 3541 831
rect 3507 750 3541 763
rect 3507 678 3541 695
rect 3507 606 3541 627
rect 3507 534 3541 559
rect 3507 462 3541 491
rect 3507 390 3541 423
rect 3507 321 3541 355
rect 3507 253 3541 284
rect 3507 185 3541 212
rect 3507 117 3541 140
rect 3507 49 3541 68
rect 3507 -19 3541 -4
rect 3507 -87 3541 -76
rect 3507 -155 3541 -148
rect 3507 -223 3541 -220
rect 3507 -258 3541 -257
rect 3507 -330 3541 -325
rect 3507 -402 3541 -393
rect 3507 -474 3541 -461
rect 3507 -546 3541 -529
rect 3507 -618 3541 -597
rect 3507 -690 3541 -665
rect 3507 -762 3541 -733
rect 3507 -834 3541 -801
rect 3507 -903 3541 -869
rect 3507 -971 3541 -940
rect 3507 -1039 3541 -1012
rect 3507 -1107 3541 -1084
rect 3507 -1175 3541 -1156
rect 3507 -1243 3541 -1228
rect 3507 -1338 3541 -1300
rect 3507 -1410 3541 -1372
rect 3507 -1482 3541 -1444
rect 3507 -1554 3541 -1516
rect 3507 -1626 3541 -1588
rect 3507 -1781 3541 -1660
rect -2458 -1815 -2293 -1781
rect -2239 -1815 -2221 -1781
rect -2171 -1815 -2149 -1781
rect -2103 -1815 -2077 -1781
rect -2035 -1815 -2005 -1781
rect -1967 -1815 -1933 -1781
rect -1899 -1815 -1865 -1781
rect -1827 -1815 -1797 -1781
rect -1755 -1815 -1729 -1781
rect -1683 -1815 -1661 -1781
rect -1611 -1815 -1593 -1781
rect -1539 -1815 -1525 -1781
rect -1467 -1815 -1457 -1781
rect -1395 -1815 -1389 -1781
rect -1323 -1815 -1321 -1781
rect -1287 -1815 -1285 -1781
rect -1219 -1815 -1213 -1781
rect -1151 -1815 -1141 -1781
rect -1083 -1815 -1069 -1781
rect -1015 -1815 -997 -1781
rect -947 -1815 -925 -1781
rect -879 -1815 -853 -1781
rect -811 -1815 -781 -1781
rect -743 -1815 -709 -1781
rect -675 -1815 -641 -1781
rect -603 -1815 -573 -1781
rect -531 -1815 -505 -1781
rect -459 -1815 -437 -1781
rect -387 -1815 -369 -1781
rect -315 -1815 -301 -1781
rect -243 -1815 -233 -1781
rect -171 -1815 -165 -1781
rect -99 -1815 -97 -1781
rect -63 -1815 -61 -1781
rect 5 -1815 11 -1781
rect 73 -1815 83 -1781
rect 141 -1815 155 -1781
rect 209 -1815 227 -1781
rect 277 -1815 299 -1781
rect 345 -1815 371 -1781
rect 413 -1815 443 -1781
rect 481 -1815 515 -1781
rect 549 -1815 583 -1781
rect 621 -1815 651 -1781
rect 693 -1815 719 -1781
rect 765 -1815 787 -1781
rect 837 -1815 855 -1781
rect 909 -1815 923 -1781
rect 981 -1815 991 -1781
rect 1025 -1815 1043 -1781
rect 1093 -1815 1115 -1781
rect 1161 -1815 1187 -1781
rect 1229 -1815 1259 -1781
rect 1297 -1815 1331 -1781
rect 1365 -1815 1399 -1781
rect 1437 -1815 1467 -1781
rect 1509 -1815 1535 -1781
rect 1581 -1815 1603 -1781
rect 1653 -1815 1671 -1781
rect 1725 -1815 1739 -1781
rect 1797 -1815 1807 -1781
rect 1869 -1815 1875 -1781
rect 1941 -1815 1943 -1781
rect 1977 -1815 1979 -1781
rect 2045 -1815 2051 -1781
rect 2113 -1815 2123 -1781
rect 2181 -1815 2195 -1781
rect 2249 -1815 2267 -1781
rect 2317 -1815 2339 -1781
rect 2385 -1815 2411 -1781
rect 2453 -1815 2483 -1781
rect 2521 -1815 2555 -1781
rect 2589 -1815 2623 -1781
rect 2661 -1815 2691 -1781
rect 2733 -1815 2759 -1781
rect 2805 -1815 2827 -1781
rect 2877 -1815 2895 -1781
rect 2949 -1815 2963 -1781
rect 3021 -1815 3031 -1781
rect 3093 -1815 3099 -1781
rect 3165 -1815 3167 -1781
rect 3201 -1815 3203 -1781
rect 3269 -1815 3275 -1781
rect 3337 -1815 3541 -1781
<< viali >>
rect -2293 2104 -2273 2138
rect -2273 2104 -2259 2138
rect -2221 2104 -2205 2138
rect -2205 2104 -2187 2138
rect -2149 2104 -2137 2138
rect -2137 2104 -2115 2138
rect -2077 2104 -2069 2138
rect -2069 2104 -2043 2138
rect -2005 2104 -2001 2138
rect -2001 2104 -1971 2138
rect -1933 2104 -1899 2138
rect -1861 2104 -1831 2138
rect -1831 2104 -1827 2138
rect -1789 2104 -1763 2138
rect -1763 2104 -1755 2138
rect -1717 2104 -1695 2138
rect -1695 2104 -1683 2138
rect -1645 2104 -1627 2138
rect -1627 2104 -1611 2138
rect -1573 2104 -1559 2138
rect -1559 2104 -1539 2138
rect -1501 2104 -1491 2138
rect -1491 2104 -1467 2138
rect -1429 2104 -1423 2138
rect -1423 2104 -1395 2138
rect -1357 2104 -1355 2138
rect -1355 2104 -1323 2138
rect -1285 2104 -1253 2138
rect -1253 2104 -1251 2138
rect -1213 2104 -1185 2138
rect -1185 2104 -1179 2138
rect -1141 2104 -1117 2138
rect -1117 2104 -1107 2138
rect -1069 2104 -1049 2138
rect -1049 2104 -1035 2138
rect -997 2104 -981 2138
rect -981 2104 -963 2138
rect -925 2104 -913 2138
rect -913 2104 -891 2138
rect -853 2104 -845 2138
rect -845 2104 -819 2138
rect -781 2104 -777 2138
rect -777 2104 -747 2138
rect -709 2104 -675 2138
rect -637 2104 -607 2138
rect -607 2104 -603 2138
rect -565 2104 -539 2138
rect -539 2104 -531 2138
rect -493 2104 -471 2138
rect -471 2104 -459 2138
rect -421 2104 -403 2138
rect -403 2104 -387 2138
rect -349 2104 -335 2138
rect -335 2104 -315 2138
rect -277 2104 -267 2138
rect -267 2104 -243 2138
rect -205 2104 -199 2138
rect -199 2104 -171 2138
rect -133 2104 -131 2138
rect -131 2104 -99 2138
rect -61 2104 -29 2138
rect -29 2104 -27 2138
rect 11 2104 39 2138
rect 39 2104 45 2138
rect 83 2104 107 2138
rect 107 2104 117 2138
rect 155 2104 175 2138
rect 175 2104 189 2138
rect 227 2104 243 2138
rect 243 2104 261 2138
rect 299 2104 311 2138
rect 311 2104 333 2138
rect 371 2104 379 2138
rect 379 2104 405 2138
rect 443 2104 447 2138
rect 447 2104 477 2138
rect 515 2104 549 2138
rect 587 2104 617 2138
rect 617 2104 621 2138
rect 659 2104 685 2138
rect 685 2104 693 2138
rect 731 2104 753 2138
rect 753 2104 765 2138
rect 803 2104 821 2138
rect 821 2104 837 2138
rect 875 2104 889 2138
rect 889 2104 909 2138
rect 947 2104 957 2138
rect 957 2104 981 2138
rect 1043 2104 1059 2138
rect 1059 2104 1077 2138
rect 1115 2104 1127 2138
rect 1127 2104 1149 2138
rect 1187 2104 1195 2138
rect 1195 2104 1221 2138
rect 1259 2104 1263 2138
rect 1263 2104 1293 2138
rect 1331 2104 1365 2138
rect 1403 2104 1433 2138
rect 1433 2104 1437 2138
rect 1475 2104 1501 2138
rect 1501 2104 1509 2138
rect 1547 2104 1569 2138
rect 1569 2104 1581 2138
rect 1619 2104 1637 2138
rect 1637 2104 1653 2138
rect 1691 2104 1705 2138
rect 1705 2104 1725 2138
rect 1763 2104 1773 2138
rect 1773 2104 1797 2138
rect 1835 2104 1841 2138
rect 1841 2104 1869 2138
rect 1907 2104 1909 2138
rect 1909 2104 1941 2138
rect 1979 2104 2011 2138
rect 2011 2104 2013 2138
rect 2051 2104 2079 2138
rect 2079 2104 2085 2138
rect 2123 2104 2147 2138
rect 2147 2104 2157 2138
rect 2195 2104 2215 2138
rect 2215 2104 2229 2138
rect 2267 2104 2283 2138
rect 2283 2104 2301 2138
rect 2339 2104 2351 2138
rect 2351 2104 2373 2138
rect 2411 2104 2419 2138
rect 2419 2104 2445 2138
rect 2483 2104 2487 2138
rect 2487 2104 2517 2138
rect 2555 2104 2589 2138
rect 2627 2104 2657 2138
rect 2657 2104 2661 2138
rect 2699 2104 2725 2138
rect 2725 2104 2733 2138
rect 2771 2104 2793 2138
rect 2793 2104 2805 2138
rect 2843 2104 2861 2138
rect 2861 2104 2877 2138
rect 2915 2104 2929 2138
rect 2929 2104 2949 2138
rect 2987 2104 2997 2138
rect 2997 2104 3021 2138
rect 3059 2104 3065 2138
rect 3065 2104 3093 2138
rect 3131 2104 3133 2138
rect 3133 2104 3165 2138
rect 3203 2104 3235 2138
rect 3235 2104 3237 2138
rect 3275 2104 3303 2138
rect 3303 2104 3309 2138
rect -2458 1953 -2424 1974
rect -2458 1940 -2424 1953
rect -2458 1885 -2424 1902
rect -2458 1868 -2424 1885
rect -2458 1817 -2424 1830
rect -2458 1796 -2424 1817
rect -2458 1749 -2424 1758
rect -2458 1724 -2424 1749
rect -2458 1681 -2424 1686
rect -2458 1652 -2424 1681
rect -2458 1613 -2424 1614
rect -2458 1580 -2424 1613
rect -2458 1511 -2424 1542
rect -2458 1508 -2424 1511
rect -2458 1443 -2424 1470
rect -2458 1436 -2424 1443
rect -2458 1375 -2424 1398
rect -2458 1364 -2424 1375
rect -2458 1307 -2424 1326
rect -2458 1292 -2424 1307
rect -2458 1239 -2424 1254
rect -2458 1220 -2424 1239
rect -2458 1171 -2424 1182
rect -2458 1148 -2424 1171
rect -2458 1103 -2424 1110
rect -2458 1076 -2424 1103
rect -2458 1035 -2424 1038
rect -2458 1004 -2424 1035
rect -2458 933 -2424 966
rect -2458 932 -2424 933
rect -2458 865 -2424 894
rect -2458 860 -2424 865
rect -2458 797 -2424 822
rect -2458 788 -2424 797
rect -2458 729 -2424 750
rect -2458 716 -2424 729
rect -2458 661 -2424 678
rect -2458 644 -2424 661
rect -2458 593 -2424 606
rect -2458 572 -2424 593
rect -2458 525 -2424 534
rect -2458 500 -2424 525
rect -2458 457 -2424 462
rect -2458 428 -2424 457
rect -2458 389 -2424 390
rect -2458 356 -2424 389
rect -2458 287 -2424 318
rect -2458 284 -2424 287
rect -2458 219 -2424 246
rect -2458 212 -2424 219
rect -2458 151 -2424 174
rect -2458 140 -2424 151
rect -2458 83 -2424 102
rect -2458 68 -2424 83
rect -2458 15 -2424 30
rect -2458 -4 -2424 15
rect -2458 -53 -2424 -42
rect -2458 -76 -2424 -53
rect -2458 -121 -2424 -114
rect -2458 -148 -2424 -121
rect -2458 -189 -2424 -186
rect -2458 -220 -2424 -189
rect -2458 -291 -2424 -258
rect -2458 -292 -2424 -291
rect -2458 -359 -2424 -330
rect -2458 -364 -2424 -359
rect -2458 -427 -2424 -402
rect -2458 -436 -2424 -427
rect -2458 -495 -2424 -474
rect -2458 -508 -2424 -495
rect -2458 -563 -2424 -546
rect -2458 -580 -2424 -563
rect -2458 -631 -2424 -618
rect -2458 -652 -2424 -631
rect -2458 -699 -2424 -690
rect -2458 -724 -2424 -699
rect -2458 -767 -2424 -762
rect -2458 -796 -2424 -767
rect -2458 -835 -2424 -834
rect -2458 -868 -2424 -835
rect -2458 -937 -2424 -906
rect -2458 -940 -2424 -937
rect -2458 -1005 -2424 -978
rect -2458 -1012 -2424 -1005
rect -2458 -1073 -2424 -1050
rect -2458 -1084 -2424 -1073
rect -2458 -1141 -2424 -1122
rect -2458 -1156 -2424 -1141
rect -2458 -1209 -2424 -1194
rect -2458 -1228 -2424 -1209
rect -2458 -1277 -2424 -1266
rect -2458 -1300 -2424 -1277
rect -2458 -1345 -2424 -1338
rect -2458 -1372 -2424 -1345
rect -2458 -1413 -2424 -1410
rect -2458 -1444 -2424 -1413
rect -2458 -1515 -2424 -1482
rect -2458 -1516 -2424 -1515
rect -2458 -1583 -2424 -1554
rect -2458 -1588 -2424 -1583
rect -2458 -1660 -2424 -1626
rect 3507 1953 3541 1974
rect 3507 1940 3541 1953
rect 3507 1885 3541 1902
rect 3507 1868 3541 1885
rect 3507 1817 3541 1830
rect 3507 1796 3541 1817
rect 3507 1749 3541 1758
rect 3507 1724 3541 1749
rect 3507 1681 3541 1686
rect 3507 1652 3541 1681
rect 3507 1613 3541 1614
rect 3507 1580 3541 1613
rect 3507 1511 3541 1542
rect 3507 1508 3541 1511
rect 3507 1443 3541 1470
rect 3507 1436 3541 1443
rect 3507 1375 3541 1398
rect 3507 1364 3541 1375
rect 3507 1307 3541 1326
rect 3507 1292 3541 1307
rect 3507 1239 3541 1254
rect 3507 1220 3541 1239
rect 3507 1171 3541 1182
rect 3507 1148 3541 1171
rect 3507 1103 3541 1110
rect 3507 1076 3541 1103
rect 3507 1035 3541 1038
rect 3507 1004 3541 1035
rect 3507 933 3541 966
rect 3507 932 3541 933
rect 3507 865 3541 894
rect 3507 860 3541 865
rect 3507 797 3541 822
rect 3507 788 3541 797
rect 3507 729 3541 750
rect 3507 716 3541 729
rect 3507 661 3541 678
rect 3507 644 3541 661
rect 3507 593 3541 606
rect 3507 572 3541 593
rect 3507 525 3541 534
rect 3507 500 3541 525
rect 3507 457 3541 462
rect 3507 428 3541 457
rect 3507 389 3541 390
rect 3507 356 3541 389
rect 3507 287 3541 318
rect 3507 284 3541 287
rect 3507 219 3541 246
rect 3507 212 3541 219
rect 3507 151 3541 174
rect 3507 140 3541 151
rect 3507 83 3541 102
rect 3507 68 3541 83
rect 3507 15 3541 30
rect 3507 -4 3541 15
rect 3507 -53 3541 -42
rect 3507 -76 3541 -53
rect 3507 -121 3541 -114
rect 3507 -148 3541 -121
rect 3507 -189 3541 -186
rect 3507 -220 3541 -189
rect 3507 -291 3541 -258
rect 3507 -292 3541 -291
rect 3507 -359 3541 -330
rect 3507 -364 3541 -359
rect 3507 -427 3541 -402
rect 3507 -436 3541 -427
rect 3507 -495 3541 -474
rect 3507 -508 3541 -495
rect 3507 -563 3541 -546
rect 3507 -580 3541 -563
rect 3507 -631 3541 -618
rect 3507 -652 3541 -631
rect 3507 -699 3541 -690
rect 3507 -724 3541 -699
rect 3507 -767 3541 -762
rect 3507 -796 3541 -767
rect 3507 -835 3541 -834
rect 3507 -868 3541 -835
rect 3507 -937 3541 -906
rect 3507 -940 3541 -937
rect 3507 -1005 3541 -978
rect 3507 -1012 3541 -1005
rect 3507 -1073 3541 -1050
rect 3507 -1084 3541 -1073
rect 3507 -1141 3541 -1122
rect 3507 -1156 3541 -1141
rect 3507 -1209 3541 -1194
rect 3507 -1228 3541 -1209
rect 3507 -1277 3541 -1266
rect 3507 -1300 3541 -1277
rect 3507 -1372 3541 -1338
rect 3507 -1444 3541 -1410
rect 3507 -1516 3541 -1482
rect 3507 -1588 3541 -1554
rect 3507 -1660 3541 -1626
rect -2293 -1815 -2273 -1781
rect -2273 -1815 -2259 -1781
rect -2221 -1815 -2205 -1781
rect -2205 -1815 -2187 -1781
rect -2149 -1815 -2137 -1781
rect -2137 -1815 -2115 -1781
rect -2077 -1815 -2069 -1781
rect -2069 -1815 -2043 -1781
rect -2005 -1815 -2001 -1781
rect -2001 -1815 -1971 -1781
rect -1933 -1815 -1899 -1781
rect -1861 -1815 -1831 -1781
rect -1831 -1815 -1827 -1781
rect -1789 -1815 -1763 -1781
rect -1763 -1815 -1755 -1781
rect -1717 -1815 -1695 -1781
rect -1695 -1815 -1683 -1781
rect -1645 -1815 -1627 -1781
rect -1627 -1815 -1611 -1781
rect -1573 -1815 -1559 -1781
rect -1559 -1815 -1539 -1781
rect -1501 -1815 -1491 -1781
rect -1491 -1815 -1467 -1781
rect -1429 -1815 -1423 -1781
rect -1423 -1815 -1395 -1781
rect -1357 -1815 -1355 -1781
rect -1355 -1815 -1323 -1781
rect -1285 -1815 -1253 -1781
rect -1253 -1815 -1251 -1781
rect -1213 -1815 -1185 -1781
rect -1185 -1815 -1179 -1781
rect -1141 -1815 -1117 -1781
rect -1117 -1815 -1107 -1781
rect -1069 -1815 -1049 -1781
rect -1049 -1815 -1035 -1781
rect -997 -1815 -981 -1781
rect -981 -1815 -963 -1781
rect -925 -1815 -913 -1781
rect -913 -1815 -891 -1781
rect -853 -1815 -845 -1781
rect -845 -1815 -819 -1781
rect -781 -1815 -777 -1781
rect -777 -1815 -747 -1781
rect -709 -1815 -675 -1781
rect -637 -1815 -607 -1781
rect -607 -1815 -603 -1781
rect -565 -1815 -539 -1781
rect -539 -1815 -531 -1781
rect -493 -1815 -471 -1781
rect -471 -1815 -459 -1781
rect -421 -1815 -403 -1781
rect -403 -1815 -387 -1781
rect -349 -1815 -335 -1781
rect -335 -1815 -315 -1781
rect -277 -1815 -267 -1781
rect -267 -1815 -243 -1781
rect -205 -1815 -199 -1781
rect -199 -1815 -171 -1781
rect -133 -1815 -131 -1781
rect -131 -1815 -99 -1781
rect -61 -1815 -29 -1781
rect -29 -1815 -27 -1781
rect 11 -1815 39 -1781
rect 39 -1815 45 -1781
rect 83 -1815 107 -1781
rect 107 -1815 117 -1781
rect 155 -1815 175 -1781
rect 175 -1815 189 -1781
rect 227 -1815 243 -1781
rect 243 -1815 261 -1781
rect 299 -1815 311 -1781
rect 311 -1815 333 -1781
rect 371 -1815 379 -1781
rect 379 -1815 405 -1781
rect 443 -1815 447 -1781
rect 447 -1815 477 -1781
rect 515 -1815 549 -1781
rect 587 -1815 617 -1781
rect 617 -1815 621 -1781
rect 659 -1815 685 -1781
rect 685 -1815 693 -1781
rect 731 -1815 753 -1781
rect 753 -1815 765 -1781
rect 803 -1815 821 -1781
rect 821 -1815 837 -1781
rect 875 -1815 889 -1781
rect 889 -1815 909 -1781
rect 947 -1815 957 -1781
rect 957 -1815 981 -1781
rect 1043 -1815 1059 -1781
rect 1059 -1815 1077 -1781
rect 1115 -1815 1127 -1781
rect 1127 -1815 1149 -1781
rect 1187 -1815 1195 -1781
rect 1195 -1815 1221 -1781
rect 1259 -1815 1263 -1781
rect 1263 -1815 1293 -1781
rect 1331 -1815 1365 -1781
rect 1403 -1815 1433 -1781
rect 1433 -1815 1437 -1781
rect 1475 -1815 1501 -1781
rect 1501 -1815 1509 -1781
rect 1547 -1815 1569 -1781
rect 1569 -1815 1581 -1781
rect 1619 -1815 1637 -1781
rect 1637 -1815 1653 -1781
rect 1691 -1815 1705 -1781
rect 1705 -1815 1725 -1781
rect 1763 -1815 1773 -1781
rect 1773 -1815 1797 -1781
rect 1835 -1815 1841 -1781
rect 1841 -1815 1869 -1781
rect 1907 -1815 1909 -1781
rect 1909 -1815 1941 -1781
rect 1979 -1815 2011 -1781
rect 2011 -1815 2013 -1781
rect 2051 -1815 2079 -1781
rect 2079 -1815 2085 -1781
rect 2123 -1815 2147 -1781
rect 2147 -1815 2157 -1781
rect 2195 -1815 2215 -1781
rect 2215 -1815 2229 -1781
rect 2267 -1815 2283 -1781
rect 2283 -1815 2301 -1781
rect 2339 -1815 2351 -1781
rect 2351 -1815 2373 -1781
rect 2411 -1815 2419 -1781
rect 2419 -1815 2445 -1781
rect 2483 -1815 2487 -1781
rect 2487 -1815 2517 -1781
rect 2555 -1815 2589 -1781
rect 2627 -1815 2657 -1781
rect 2657 -1815 2661 -1781
rect 2699 -1815 2725 -1781
rect 2725 -1815 2733 -1781
rect 2771 -1815 2793 -1781
rect 2793 -1815 2805 -1781
rect 2843 -1815 2861 -1781
rect 2861 -1815 2877 -1781
rect 2915 -1815 2929 -1781
rect 2929 -1815 2949 -1781
rect 2987 -1815 2997 -1781
rect 2997 -1815 3021 -1781
rect 3059 -1815 3065 -1781
rect 3065 -1815 3093 -1781
rect 3131 -1815 3133 -1781
rect 3133 -1815 3165 -1781
rect 3203 -1815 3235 -1781
rect 3235 -1815 3237 -1781
rect 3275 -1815 3303 -1781
rect 3303 -1815 3309 -1781
<< metal1 >>
rect -2476 2138 3566 2163
rect -2476 2104 -2293 2138
rect -2259 2104 -2221 2138
rect -2187 2104 -2149 2138
rect -2115 2104 -2077 2138
rect -2043 2104 -2005 2138
rect -1971 2104 -1933 2138
rect -1899 2104 -1861 2138
rect -1827 2104 -1789 2138
rect -1755 2104 -1717 2138
rect -1683 2104 -1645 2138
rect -1611 2104 -1573 2138
rect -1539 2104 -1501 2138
rect -1467 2104 -1429 2138
rect -1395 2104 -1357 2138
rect -1323 2104 -1285 2138
rect -1251 2104 -1213 2138
rect -1179 2104 -1141 2138
rect -1107 2104 -1069 2138
rect -1035 2104 -997 2138
rect -963 2104 -925 2138
rect -891 2104 -853 2138
rect -819 2104 -781 2138
rect -747 2104 -709 2138
rect -675 2104 -637 2138
rect -603 2104 -565 2138
rect -531 2104 -493 2138
rect -459 2104 -421 2138
rect -387 2104 -349 2138
rect -315 2104 -277 2138
rect -243 2104 -205 2138
rect -171 2104 -133 2138
rect -99 2104 -61 2138
rect -27 2104 11 2138
rect 45 2104 83 2138
rect 117 2104 155 2138
rect 189 2104 227 2138
rect 261 2104 299 2138
rect 333 2104 371 2138
rect 405 2104 443 2138
rect 477 2104 515 2138
rect 549 2104 587 2138
rect 621 2104 659 2138
rect 693 2104 731 2138
rect 765 2104 803 2138
rect 837 2104 875 2138
rect 909 2104 947 2138
rect 981 2104 1043 2138
rect 1077 2104 1115 2138
rect 1149 2104 1187 2138
rect 1221 2104 1259 2138
rect 1293 2104 1331 2138
rect 1365 2104 1403 2138
rect 1437 2104 1475 2138
rect 1509 2104 1547 2138
rect 1581 2104 1619 2138
rect 1653 2104 1691 2138
rect 1725 2104 1763 2138
rect 1797 2104 1835 2138
rect 1869 2104 1907 2138
rect 1941 2104 1979 2138
rect 2013 2104 2051 2138
rect 2085 2104 2123 2138
rect 2157 2104 2195 2138
rect 2229 2104 2267 2138
rect 2301 2104 2339 2138
rect 2373 2104 2411 2138
rect 2445 2104 2483 2138
rect 2517 2104 2555 2138
rect 2589 2104 2627 2138
rect 2661 2104 2699 2138
rect 2733 2104 2771 2138
rect 2805 2104 2843 2138
rect 2877 2104 2915 2138
rect 2949 2104 2987 2138
rect 3021 2104 3059 2138
rect 3093 2104 3131 2138
rect 3165 2104 3203 2138
rect 3237 2104 3275 2138
rect 3309 2104 3566 2138
rect -2476 1974 3566 2104
rect -2476 1940 -2458 1974
rect -2424 1940 3507 1974
rect 3541 1940 3566 1974
rect -2476 1902 3566 1940
rect -2476 1868 -2458 1902
rect -2424 1868 3507 1902
rect 3541 1868 3566 1902
rect -2476 1830 3566 1868
rect -2476 1796 -2458 1830
rect -2424 1796 3507 1830
rect 3541 1796 3566 1830
rect -2476 1758 3566 1796
rect -2476 1724 -2458 1758
rect -2424 1746 3507 1758
rect -2424 1724 -1727 1746
rect -2476 1686 -1727 1724
rect -2476 1652 -2458 1686
rect -2424 1652 -1727 1686
rect -2476 1614 -1727 1652
rect -2476 1580 -2458 1614
rect -2424 1580 -1727 1614
rect -2476 1542 -1727 1580
rect -2476 1508 -2458 1542
rect -2424 1508 -1727 1542
rect -2476 1470 -1727 1508
rect -2476 1436 -2458 1470
rect -2424 1436 -1727 1470
rect -1512 1500 -1316 1510
rect -1512 1448 -1503 1500
rect -1451 1448 -1439 1500
rect -1387 1448 -1375 1500
rect -1323 1448 -1316 1500
rect -1512 1440 -1316 1448
rect -2476 1398 -1727 1436
rect -2476 1364 -2458 1398
rect -2424 1364 -1727 1398
rect -2476 1326 -1727 1364
rect -2476 1292 -2458 1326
rect -2424 1292 -1727 1326
rect -2476 1254 -1727 1292
rect -1436 1289 -1390 1440
rect -778 1403 -678 1746
rect -141 1640 55 1650
rect -141 1588 -134 1640
rect -82 1588 -70 1640
rect -18 1588 -6 1640
rect 46 1588 55 1640
rect -141 1580 55 1588
rect -2476 1220 -2458 1254
rect -2424 1220 -1727 1254
rect -2476 1182 -1727 1220
rect -920 1203 -537 1403
rect -67 1289 -21 1580
rect 200 1500 396 1510
rect 200 1448 207 1500
rect 259 1448 271 1500
rect 323 1448 335 1500
rect 387 1448 396 1500
rect 200 1440 396 1448
rect 270 1289 316 1440
rect 929 1403 1029 1746
rect 2635 1724 3507 1746
rect 3541 1724 3566 1758
rect 2635 1686 3566 1724
rect 2635 1652 3507 1686
rect 3541 1652 3566 1686
rect 1559 1640 1755 1650
rect 1559 1588 1568 1640
rect 1620 1588 1632 1640
rect 1684 1588 1696 1640
rect 1748 1588 1755 1640
rect 1559 1580 1755 1588
rect 2635 1614 3566 1652
rect 2635 1580 3507 1614
rect 3541 1580 3566 1614
rect 786 1203 1170 1403
rect 1640 1289 1686 1580
rect 2635 1542 3566 1580
rect 1903 1500 2099 1510
rect 1903 1448 1912 1500
rect 1964 1448 1976 1500
rect 2028 1448 2040 1500
rect 2092 1448 2099 1500
rect 1903 1440 2099 1448
rect 2635 1508 3507 1542
rect 3541 1508 3566 1542
rect 2635 1470 3566 1508
rect 1977 1289 2023 1440
rect 2635 1436 3507 1470
rect 3541 1436 3566 1470
rect 2635 1403 3566 1436
rect 2493 1398 3566 1403
rect 2493 1364 3507 1398
rect 3541 1364 3566 1398
rect 2493 1326 3566 1364
rect 2493 1292 3507 1326
rect 3541 1292 3566 1326
rect 2493 1254 3566 1292
rect 2493 1220 3507 1254
rect 3541 1220 3566 1254
rect 2493 1203 3566 1220
rect -2476 1148 -2458 1182
rect -2424 1148 -1727 1182
rect -2476 1110 -1727 1148
rect -2476 1076 -2458 1110
rect -2424 1076 -1727 1110
rect -2476 1038 -1727 1076
rect -1436 1101 -930 1171
rect -1436 1049 -1360 1101
rect -1308 1049 -1296 1101
rect -1244 1049 -1232 1101
rect -1180 1049 -1139 1101
rect -1087 1049 -1075 1101
rect -1023 1049 -1011 1101
rect -959 1049 -930 1101
rect -1436 1041 -930 1049
rect -2476 1004 -2458 1038
rect -2424 1004 -1727 1038
rect -2476 966 -1727 1004
rect -2476 932 -2458 966
rect -2424 932 -1727 966
rect -2476 894 -1727 932
rect -2476 860 -2458 894
rect -2424 860 -1727 894
rect -2476 822 -1727 860
rect -2476 788 -2458 822
rect -2424 788 -1727 822
rect -2476 750 -1727 788
rect -2476 716 -2458 750
rect -2424 716 -1727 750
rect -2476 678 -1727 716
rect -2476 644 -2458 678
rect -2424 644 -1727 678
rect -2476 606 -1727 644
rect -2476 572 -2458 606
rect -2424 572 -1727 606
rect -2476 534 -1727 572
rect -2476 500 -2458 534
rect -2424 500 -1727 534
rect -2476 462 -1727 500
rect -2476 428 -2458 462
rect -2424 428 -1727 462
rect -1436 800 -930 810
rect -1436 748 -1360 800
rect -1308 748 -1296 800
rect -1244 748 -1232 800
rect -1180 748 -1139 800
rect -1087 748 -1075 800
rect -1023 748 -1011 800
rect -959 748 -930 800
rect -1436 530 -930 748
rect -1436 453 -1390 530
rect -778 498 -678 1203
rect -527 951 -21 1171
rect 270 1101 776 1171
rect 270 1049 351 1101
rect 403 1049 415 1101
rect 467 1049 479 1101
rect 531 1049 572 1101
rect 624 1049 636 1101
rect 688 1049 700 1101
rect 752 1049 776 1101
rect 270 1041 776 1049
rect -527 899 -501 951
rect -449 899 -437 951
rect -385 899 -373 951
rect -321 899 -280 951
rect -228 899 -216 951
rect -164 899 -152 951
rect -100 899 -21 951
rect -527 891 -21 899
rect 270 800 776 810
rect 270 748 351 800
rect 403 748 415 800
rect 467 748 479 800
rect 531 748 572 800
rect 624 748 636 800
rect 688 748 700 800
rect 752 748 776 800
rect -527 650 -21 660
rect -527 598 -501 650
rect -449 598 -437 650
rect -385 598 -373 650
rect -321 598 -280 650
rect -228 598 -216 650
rect -164 598 -152 650
rect -100 598 -21 650
rect -527 530 -21 598
rect -2476 390 -1727 428
rect -2476 356 -2458 390
rect -2424 356 -1727 390
rect -2476 318 -1727 356
rect -2476 284 -2458 318
rect -2424 284 -1727 318
rect -920 298 -537 498
rect -67 453 -21 530
rect 270 530 776 748
rect 270 453 316 530
rect 929 498 1029 1203
rect 2635 1182 3566 1203
rect 1180 951 1686 1171
rect 1977 1101 2483 1171
rect 1977 1049 2056 1101
rect 2108 1049 2120 1101
rect 2172 1049 2184 1101
rect 2236 1049 2277 1101
rect 2329 1049 2341 1101
rect 2393 1049 2405 1101
rect 2457 1049 2483 1101
rect 1977 1041 2483 1049
rect 2635 1148 3507 1182
rect 3541 1148 3566 1182
rect 2635 1110 3566 1148
rect 2635 1076 3507 1110
rect 3541 1076 3566 1110
rect 1180 899 1206 951
rect 1258 899 1270 951
rect 1322 899 1334 951
rect 1386 899 1427 951
rect 1479 899 1491 951
rect 1543 899 1555 951
rect 1607 899 1686 951
rect 1180 891 1686 899
rect 2635 1038 3566 1076
rect 2635 1004 3507 1038
rect 3541 1004 3566 1038
rect 2635 966 3566 1004
rect 2635 932 3507 966
rect 3541 932 3566 966
rect 2635 894 3566 932
rect 2635 860 3507 894
rect 3541 860 3566 894
rect 2635 822 3566 860
rect 1977 800 2483 810
rect 1977 748 2056 800
rect 2108 748 2120 800
rect 2172 748 2184 800
rect 2236 748 2277 800
rect 2329 748 2341 800
rect 2393 748 2405 800
rect 2457 748 2483 800
rect 1180 650 1686 660
rect 1180 598 1206 650
rect 1258 598 1270 650
rect 1322 598 1334 650
rect 1386 598 1427 650
rect 1479 598 1491 650
rect 1543 598 1555 650
rect 1607 598 1686 650
rect 1180 530 1686 598
rect 786 298 1170 498
rect 1640 453 1686 530
rect 1977 530 2483 748
rect 2635 788 3507 822
rect 3541 788 3566 822
rect 2635 750 3566 788
rect 2635 716 3507 750
rect 3541 716 3566 750
rect 2635 678 3566 716
rect 2635 644 3507 678
rect 3541 644 3566 678
rect 2635 606 3566 644
rect 2635 572 3507 606
rect 3541 572 3566 606
rect 2635 534 3566 572
rect 1977 453 2023 530
rect 2635 500 3507 534
rect 3541 500 3566 534
rect 2635 498 3566 500
rect 2493 462 3566 498
rect 2493 428 3507 462
rect 3541 428 3566 462
rect 2493 390 3566 428
rect 2493 356 3507 390
rect 3541 356 3566 390
rect 2493 318 3566 356
rect 2493 298 3507 318
rect -2476 246 -1727 284
rect -2476 212 -2458 246
rect -2424 212 -1727 246
rect -2476 174 -1727 212
rect -2476 140 -2458 174
rect -2424 140 -1727 174
rect -2476 102 -1727 140
rect -2476 68 -2458 102
rect -2424 68 -1727 102
rect -2476 30 -1727 68
rect -2476 -4 -2458 30
rect -2424 -4 -1727 30
rect -778 26 -678 298
rect 195 251 391 261
rect 195 199 204 251
rect 256 199 268 251
rect 320 199 332 251
rect 384 199 391 251
rect 195 191 391 199
rect -146 122 50 132
rect -146 70 -137 122
rect -85 70 -73 122
rect -21 70 -9 122
rect 43 70 50 122
rect -146 62 50 70
rect -2476 -42 -1727 -4
rect -2476 -76 -2458 -42
rect -2424 -76 -1727 -42
rect -2476 -114 -1727 -76
rect -2476 -148 -2458 -114
rect -2424 -148 -1727 -114
rect -2476 -186 -1727 -148
rect -2476 -220 -2458 -186
rect -2424 -220 -1727 -186
rect -2476 -258 -1727 -220
rect -2476 -292 -2458 -258
rect -2424 -292 -1727 -258
rect -2476 -330 -1727 -292
rect -2476 -364 -2458 -330
rect -2424 -364 -1727 -330
rect -2476 -402 -1727 -364
rect -2476 -436 -2458 -402
rect -2424 -436 -1727 -402
rect -2476 -474 -1727 -436
rect -2476 -508 -2458 -474
rect -2424 -508 -1727 -474
rect -1436 -206 -1390 -136
rect -920 -174 -537 26
rect -67 -105 -21 62
rect 270 -105 316 191
rect 929 26 1029 298
rect 2635 284 3507 298
rect 3541 284 3566 318
rect 2635 246 3566 284
rect 2635 212 3507 246
rect 3541 212 3566 246
rect 2635 174 3566 212
rect 2635 140 3507 174
rect 3541 140 3566 174
rect 1559 122 1755 132
rect 1559 70 1568 122
rect 1620 70 1632 122
rect 1684 70 1696 122
rect 1748 70 1755 122
rect 1559 62 1755 70
rect 2635 102 3566 140
rect 2635 68 3507 102
rect 3541 68 3566 102
rect -1436 -427 -930 -206
rect -1436 -479 -1354 -427
rect -1302 -479 -1290 -427
rect -1238 -479 -1226 -427
rect -1174 -479 -1133 -427
rect -1081 -479 -1069 -427
rect -1017 -479 -1005 -427
rect -953 -479 -930 -427
rect -1436 -487 -930 -479
rect -2476 -546 -1727 -508
rect -2476 -580 -2458 -546
rect -2424 -580 -1727 -546
rect -2476 -618 -1727 -580
rect -2476 -652 -2458 -618
rect -2424 -652 -1727 -618
rect -2476 -690 -1727 -652
rect -2476 -724 -2458 -690
rect -2424 -724 -1727 -690
rect -2476 -762 -1727 -724
rect -2476 -796 -2458 -762
rect -2424 -796 -1727 -762
rect -2476 -834 -1727 -796
rect -2476 -868 -2458 -834
rect -2424 -868 -1727 -834
rect -1436 -728 -930 -718
rect -1436 -780 -1354 -728
rect -1302 -780 -1290 -728
rect -1238 -780 -1226 -728
rect -1174 -780 -1133 -728
rect -1081 -780 -1069 -728
rect -1017 -780 -1005 -728
rect -953 -780 -930 -728
rect -1436 -848 -930 -780
rect -2476 -906 -1727 -868
rect -778 -880 -678 -174
rect -67 -206 -21 -136
rect -527 -276 -21 -206
rect -527 -328 -501 -276
rect -449 -328 -437 -276
rect -385 -328 -373 -276
rect -321 -328 -280 -276
rect -228 -328 -216 -276
rect -164 -328 -152 -276
rect -100 -328 -21 -276
rect -527 -336 -21 -328
rect 270 -206 316 -136
rect 786 -174 1170 26
rect 1640 -105 1686 62
rect 2635 30 3566 68
rect 2635 26 3507 30
rect 2493 -4 3507 26
rect 3541 -4 3566 30
rect 2493 -42 3566 -4
rect 2493 -76 3507 -42
rect 3541 -76 3566 -42
rect 2493 -114 3566 -76
rect 270 -427 776 -206
rect 270 -479 349 -427
rect 401 -479 413 -427
rect 465 -479 477 -427
rect 529 -479 570 -427
rect 622 -479 634 -427
rect 686 -479 698 -427
rect 750 -479 776 -427
rect 270 -487 776 -479
rect -527 -577 -21 -567
rect -527 -629 -501 -577
rect -449 -629 -437 -577
rect -385 -629 -373 -577
rect -321 -629 -280 -577
rect -228 -629 -216 -577
rect -164 -629 -152 -577
rect -100 -629 -21 -577
rect -527 -848 -21 -629
rect 270 -728 776 -718
rect 270 -780 349 -728
rect 401 -780 413 -728
rect 465 -780 477 -728
rect 529 -780 570 -728
rect 622 -780 634 -728
rect 686 -780 698 -728
rect 750 -780 776 -728
rect 270 -848 776 -780
rect 929 -880 1029 -174
rect 1640 -206 1686 -136
rect 1180 -276 1686 -206
rect 1180 -328 1206 -276
rect 1258 -328 1270 -276
rect 1322 -328 1334 -276
rect 1386 -328 1427 -276
rect 1479 -328 1491 -276
rect 1543 -328 1555 -276
rect 1607 -328 1686 -276
rect 1180 -336 1686 -328
rect 1977 -206 2023 -136
rect 2493 -148 3507 -114
rect 3541 -148 3566 -114
rect 2493 -174 3566 -148
rect 2635 -186 3566 -174
rect 1977 -427 2483 -206
rect 1977 -479 2056 -427
rect 2108 -479 2120 -427
rect 2172 -479 2184 -427
rect 2236 -479 2277 -427
rect 2329 -479 2341 -427
rect 2393 -479 2405 -427
rect 2457 -479 2483 -427
rect 1977 -487 2483 -479
rect 2635 -220 3507 -186
rect 3541 -220 3566 -186
rect 2635 -258 3566 -220
rect 2635 -292 3507 -258
rect 3541 -292 3566 -258
rect 2635 -330 3566 -292
rect 2635 -364 3507 -330
rect 3541 -364 3566 -330
rect 2635 -402 3566 -364
rect 2635 -436 3507 -402
rect 3541 -436 3566 -402
rect 2635 -474 3566 -436
rect 2635 -508 3507 -474
rect 3541 -508 3566 -474
rect 2635 -546 3566 -508
rect 1180 -577 1686 -567
rect 1180 -629 1206 -577
rect 1258 -629 1270 -577
rect 1322 -629 1334 -577
rect 1386 -629 1427 -577
rect 1479 -629 1491 -577
rect 1543 -629 1555 -577
rect 1607 -629 1686 -577
rect 1180 -848 1686 -629
rect 2635 -580 3507 -546
rect 3541 -580 3566 -546
rect 2635 -618 3566 -580
rect 2635 -652 3507 -618
rect 3541 -652 3566 -618
rect 2635 -690 3566 -652
rect 1977 -728 2483 -718
rect 1977 -780 2056 -728
rect 2108 -780 2120 -728
rect 2172 -780 2184 -728
rect 2236 -780 2277 -728
rect 2329 -780 2341 -728
rect 2393 -780 2405 -728
rect 2457 -780 2483 -728
rect 1977 -848 2483 -780
rect 2635 -724 3507 -690
rect 3541 -724 3566 -690
rect 2635 -762 3566 -724
rect 2635 -796 3507 -762
rect 3541 -796 3566 -762
rect 2635 -834 3566 -796
rect 2635 -868 3507 -834
rect 3541 -868 3566 -834
rect 2635 -880 3566 -868
rect -2476 -940 -2458 -906
rect -2424 -940 -1727 -906
rect -2476 -978 -1727 -940
rect -2476 -1012 -2458 -978
rect -2424 -1012 -1727 -978
rect -2476 -1050 -1727 -1012
rect -2476 -1084 -2458 -1050
rect -2424 -1084 -1727 -1050
rect -2476 -1122 -1727 -1084
rect -1436 -1116 -1390 -946
rect -920 -1080 -537 -880
rect -2476 -1156 -2458 -1122
rect -2424 -1156 -1727 -1122
rect -2476 -1194 -1727 -1156
rect -1512 -1126 -1316 -1116
rect -1512 -1178 -1503 -1126
rect -1451 -1178 -1439 -1126
rect -1387 -1178 -1375 -1126
rect -1323 -1178 -1316 -1126
rect -1512 -1186 -1316 -1178
rect -2476 -1228 -2458 -1194
rect -2424 -1228 -1727 -1194
rect -2476 -1266 -1727 -1228
rect -2476 -1300 -2458 -1266
rect -2424 -1300 -1727 -1266
rect -2476 -1338 -1727 -1300
rect -2476 -1372 -2458 -1338
rect -2424 -1372 -1727 -1338
rect -2476 -1410 -1727 -1372
rect -2476 -1444 -2458 -1410
rect -2424 -1422 -1727 -1410
rect -778 -1422 -678 -1080
rect -67 -1256 -21 -946
rect 270 -1116 316 -946
rect 786 -1080 1170 -880
rect 2493 -906 3566 -880
rect 2493 -940 3507 -906
rect 3541 -940 3566 -906
rect 200 -1126 396 -1116
rect 200 -1178 207 -1126
rect 259 -1178 271 -1126
rect 323 -1178 335 -1126
rect 387 -1178 396 -1126
rect 200 -1186 396 -1178
rect -141 -1266 55 -1256
rect -141 -1318 -134 -1266
rect -82 -1318 -70 -1266
rect -18 -1318 -6 -1266
rect 46 -1318 55 -1266
rect -141 -1326 55 -1318
rect 929 -1422 1029 -1080
rect 1640 -1256 1686 -946
rect 1977 -1116 2023 -946
rect 2493 -978 3566 -940
rect 2493 -1012 3507 -978
rect 3541 -1012 3566 -978
rect 2493 -1050 3566 -1012
rect 2493 -1080 3507 -1050
rect 2635 -1084 3507 -1080
rect 3541 -1084 3566 -1050
rect 1903 -1126 2099 -1116
rect 1903 -1178 1912 -1126
rect 1964 -1178 1976 -1126
rect 2028 -1178 2040 -1126
rect 2092 -1178 2099 -1126
rect 1903 -1186 2099 -1178
rect 2635 -1122 3566 -1084
rect 2635 -1156 3507 -1122
rect 3541 -1156 3566 -1122
rect 2635 -1194 3566 -1156
rect 2635 -1228 3507 -1194
rect 3541 -1228 3566 -1194
rect 1559 -1266 1755 -1256
rect 1559 -1318 1568 -1266
rect 1620 -1318 1632 -1266
rect 1684 -1318 1696 -1266
rect 1748 -1318 1755 -1266
rect 1559 -1326 1755 -1318
rect 2635 -1266 3566 -1228
rect 2635 -1300 3507 -1266
rect 3541 -1300 3566 -1266
rect 2635 -1338 3566 -1300
rect 2635 -1372 3507 -1338
rect 3541 -1372 3566 -1338
rect 2635 -1410 3566 -1372
rect 2635 -1422 3507 -1410
rect -2424 -1444 3507 -1422
rect 3541 -1444 3566 -1410
rect -2476 -1482 3566 -1444
rect -2476 -1516 -2458 -1482
rect -2424 -1516 3507 -1482
rect 3541 -1516 3566 -1482
rect -2476 -1554 3566 -1516
rect -2476 -1588 -2458 -1554
rect -2424 -1588 3507 -1554
rect 3541 -1588 3566 -1554
rect -2476 -1626 3566 -1588
rect -2476 -1660 -2458 -1626
rect -2424 -1660 3507 -1626
rect 3541 -1660 3566 -1626
rect -2476 -1781 3566 -1660
rect -2476 -1815 -2293 -1781
rect -2259 -1815 -2221 -1781
rect -2187 -1815 -2149 -1781
rect -2115 -1815 -2077 -1781
rect -2043 -1815 -2005 -1781
rect -1971 -1815 -1933 -1781
rect -1899 -1815 -1861 -1781
rect -1827 -1815 -1789 -1781
rect -1755 -1815 -1717 -1781
rect -1683 -1815 -1645 -1781
rect -1611 -1815 -1573 -1781
rect -1539 -1815 -1501 -1781
rect -1467 -1815 -1429 -1781
rect -1395 -1815 -1357 -1781
rect -1323 -1815 -1285 -1781
rect -1251 -1815 -1213 -1781
rect -1179 -1815 -1141 -1781
rect -1107 -1815 -1069 -1781
rect -1035 -1815 -997 -1781
rect -963 -1815 -925 -1781
rect -891 -1815 -853 -1781
rect -819 -1815 -781 -1781
rect -747 -1815 -709 -1781
rect -675 -1815 -637 -1781
rect -603 -1815 -565 -1781
rect -531 -1815 -493 -1781
rect -459 -1815 -421 -1781
rect -387 -1815 -349 -1781
rect -315 -1815 -277 -1781
rect -243 -1815 -205 -1781
rect -171 -1815 -133 -1781
rect -99 -1815 -61 -1781
rect -27 -1815 11 -1781
rect 45 -1815 83 -1781
rect 117 -1815 155 -1781
rect 189 -1815 227 -1781
rect 261 -1815 299 -1781
rect 333 -1815 371 -1781
rect 405 -1815 443 -1781
rect 477 -1815 515 -1781
rect 549 -1815 587 -1781
rect 621 -1815 659 -1781
rect 693 -1815 731 -1781
rect 765 -1815 803 -1781
rect 837 -1815 875 -1781
rect 909 -1815 947 -1781
rect 981 -1815 1043 -1781
rect 1077 -1815 1115 -1781
rect 1149 -1815 1187 -1781
rect 1221 -1815 1259 -1781
rect 1293 -1815 1331 -1781
rect 1365 -1815 1403 -1781
rect 1437 -1815 1475 -1781
rect 1509 -1815 1547 -1781
rect 1581 -1815 1619 -1781
rect 1653 -1815 1691 -1781
rect 1725 -1815 1763 -1781
rect 1797 -1815 1835 -1781
rect 1869 -1815 1907 -1781
rect 1941 -1815 1979 -1781
rect 2013 -1815 2051 -1781
rect 2085 -1815 2123 -1781
rect 2157 -1815 2195 -1781
rect 2229 -1815 2267 -1781
rect 2301 -1815 2339 -1781
rect 2373 -1815 2411 -1781
rect 2445 -1815 2483 -1781
rect 2517 -1815 2555 -1781
rect 2589 -1815 2627 -1781
rect 2661 -1815 2699 -1781
rect 2733 -1815 2771 -1781
rect 2805 -1815 2843 -1781
rect 2877 -1815 2915 -1781
rect 2949 -1815 2987 -1781
rect 3021 -1815 3059 -1781
rect 3093 -1815 3131 -1781
rect 3165 -1815 3203 -1781
rect 3237 -1815 3275 -1781
rect 3309 -1815 3566 -1781
rect -2476 -1840 3566 -1815
<< via1 >>
rect -1503 1448 -1451 1500
rect -1439 1448 -1387 1500
rect -1375 1448 -1323 1500
rect -134 1588 -82 1640
rect -70 1588 -18 1640
rect -6 1588 46 1640
rect 207 1448 259 1500
rect 271 1448 323 1500
rect 335 1448 387 1500
rect 1568 1588 1620 1640
rect 1632 1588 1684 1640
rect 1696 1588 1748 1640
rect 1912 1448 1964 1500
rect 1976 1448 2028 1500
rect 2040 1448 2092 1500
rect -1360 1049 -1308 1101
rect -1296 1049 -1244 1101
rect -1232 1049 -1180 1101
rect -1139 1049 -1087 1101
rect -1075 1049 -1023 1101
rect -1011 1049 -959 1101
rect -1360 748 -1308 800
rect -1296 748 -1244 800
rect -1232 748 -1180 800
rect -1139 748 -1087 800
rect -1075 748 -1023 800
rect -1011 748 -959 800
rect 351 1049 403 1101
rect 415 1049 467 1101
rect 479 1049 531 1101
rect 572 1049 624 1101
rect 636 1049 688 1101
rect 700 1049 752 1101
rect -501 899 -449 951
rect -437 899 -385 951
rect -373 899 -321 951
rect -280 899 -228 951
rect -216 899 -164 951
rect -152 899 -100 951
rect 351 748 403 800
rect 415 748 467 800
rect 479 748 531 800
rect 572 748 624 800
rect 636 748 688 800
rect 700 748 752 800
rect -501 598 -449 650
rect -437 598 -385 650
rect -373 598 -321 650
rect -280 598 -228 650
rect -216 598 -164 650
rect -152 598 -100 650
rect 2056 1049 2108 1101
rect 2120 1049 2172 1101
rect 2184 1049 2236 1101
rect 2277 1049 2329 1101
rect 2341 1049 2393 1101
rect 2405 1049 2457 1101
rect 1206 899 1258 951
rect 1270 899 1322 951
rect 1334 899 1386 951
rect 1427 899 1479 951
rect 1491 899 1543 951
rect 1555 899 1607 951
rect 2056 748 2108 800
rect 2120 748 2172 800
rect 2184 748 2236 800
rect 2277 748 2329 800
rect 2341 748 2393 800
rect 2405 748 2457 800
rect 1206 598 1258 650
rect 1270 598 1322 650
rect 1334 598 1386 650
rect 1427 598 1479 650
rect 1491 598 1543 650
rect 1555 598 1607 650
rect 204 199 256 251
rect 268 199 320 251
rect 332 199 384 251
rect -137 70 -85 122
rect -73 70 -21 122
rect -9 70 43 122
rect 1568 70 1620 122
rect 1632 70 1684 122
rect 1696 70 1748 122
rect -1354 -479 -1302 -427
rect -1290 -479 -1238 -427
rect -1226 -479 -1174 -427
rect -1133 -479 -1081 -427
rect -1069 -479 -1017 -427
rect -1005 -479 -953 -427
rect -1354 -780 -1302 -728
rect -1290 -780 -1238 -728
rect -1226 -780 -1174 -728
rect -1133 -780 -1081 -728
rect -1069 -780 -1017 -728
rect -1005 -780 -953 -728
rect -501 -328 -449 -276
rect -437 -328 -385 -276
rect -373 -328 -321 -276
rect -280 -328 -228 -276
rect -216 -328 -164 -276
rect -152 -328 -100 -276
rect 349 -479 401 -427
rect 413 -479 465 -427
rect 477 -479 529 -427
rect 570 -479 622 -427
rect 634 -479 686 -427
rect 698 -479 750 -427
rect -501 -629 -449 -577
rect -437 -629 -385 -577
rect -373 -629 -321 -577
rect -280 -629 -228 -577
rect -216 -629 -164 -577
rect -152 -629 -100 -577
rect 349 -780 401 -728
rect 413 -780 465 -728
rect 477 -780 529 -728
rect 570 -780 622 -728
rect 634 -780 686 -728
rect 698 -780 750 -728
rect 1206 -328 1258 -276
rect 1270 -328 1322 -276
rect 1334 -328 1386 -276
rect 1427 -328 1479 -276
rect 1491 -328 1543 -276
rect 1555 -328 1607 -276
rect 2056 -479 2108 -427
rect 2120 -479 2172 -427
rect 2184 -479 2236 -427
rect 2277 -479 2329 -427
rect 2341 -479 2393 -427
rect 2405 -479 2457 -427
rect 1206 -629 1258 -577
rect 1270 -629 1322 -577
rect 1334 -629 1386 -577
rect 1427 -629 1479 -577
rect 1491 -629 1543 -577
rect 1555 -629 1607 -577
rect 2056 -780 2108 -728
rect 2120 -780 2172 -728
rect 2184 -780 2236 -728
rect 2277 -780 2329 -728
rect 2341 -780 2393 -728
rect 2405 -780 2457 -728
rect -1503 -1178 -1451 -1126
rect -1439 -1178 -1387 -1126
rect -1375 -1178 -1323 -1126
rect 207 -1178 259 -1126
rect 271 -1178 323 -1126
rect 335 -1178 387 -1126
rect -134 -1318 -82 -1266
rect -70 -1318 -18 -1266
rect -6 -1318 46 -1266
rect 1912 -1178 1964 -1126
rect 1976 -1178 2028 -1126
rect 2040 -1178 2092 -1126
rect 1568 -1318 1620 -1266
rect 1632 -1318 1684 -1266
rect 1696 -1318 1748 -1266
<< metal2 >>
rect 1715 1658 2015 1680
rect 1715 1650 1755 1658
rect -1380 1640 1755 1650
rect -1380 1588 -134 1640
rect -82 1588 -70 1640
rect -18 1588 -6 1640
rect 46 1588 1568 1640
rect 1620 1588 1632 1640
rect 1684 1588 1696 1640
rect 1748 1602 1755 1640
rect 1811 1602 1835 1658
rect 1891 1602 1915 1658
rect 1971 1650 2015 1658
rect 1971 1602 2483 1650
rect 1748 1588 2483 1602
rect -1380 1580 2483 1588
rect -60 1518 240 1540
rect -60 1510 -20 1518
rect -1512 1500 -20 1510
rect -1512 1448 -1503 1500
rect -1451 1448 -1439 1500
rect -1387 1448 -1375 1500
rect -1323 1462 -20 1500
rect 36 1462 60 1518
rect 116 1462 140 1518
rect 196 1510 240 1518
rect 196 1500 2483 1510
rect 196 1462 207 1500
rect -1323 1448 207 1462
rect 259 1448 271 1500
rect 323 1448 335 1500
rect 387 1448 1912 1500
rect 1964 1448 1976 1500
rect 2028 1448 2040 1500
rect 2092 1448 2483 1500
rect -1512 1440 2483 1448
rect -1380 1101 2483 1111
rect -1380 1049 -1360 1101
rect -1308 1049 -1296 1101
rect -1244 1049 -1232 1101
rect -1180 1049 -1139 1101
rect -1087 1049 -1075 1101
rect -1023 1049 -1011 1101
rect -959 1089 351 1101
rect -959 1049 -838 1089
rect -1380 1041 -838 1049
rect -878 1033 -838 1041
rect -782 1033 -758 1089
rect -702 1033 -678 1089
rect -622 1049 351 1089
rect 403 1049 415 1101
rect 467 1049 479 1101
rect 531 1049 572 1101
rect 624 1049 636 1101
rect 688 1049 700 1101
rect 752 1049 2056 1101
rect 2108 1049 2120 1101
rect 2172 1049 2184 1101
rect 2236 1049 2277 1101
rect 2329 1049 2341 1101
rect 2393 1049 2405 1101
rect 2457 1049 2483 1101
rect -622 1041 2483 1049
rect -622 1033 -578 1041
rect -878 1011 -578 1033
rect -1380 951 2483 961
rect -1380 899 -501 951
rect -449 899 -437 951
rect -385 899 -373 951
rect -321 899 -280 951
rect -228 899 -216 951
rect -164 899 -152 951
rect -100 939 1206 951
rect -100 899 865 939
rect -1380 891 865 899
rect 825 883 865 891
rect 921 883 945 939
rect 1001 883 1025 939
rect 1081 899 1206 939
rect 1258 899 1270 951
rect 1322 899 1334 951
rect 1386 899 1427 951
rect 1479 899 1491 951
rect 1543 899 1555 951
rect 1607 899 2483 951
rect 1081 891 2483 899
rect 1081 883 1125 891
rect 825 861 1125 883
rect -878 818 -578 840
rect -878 810 -838 818
rect -1380 800 -838 810
rect -1380 748 -1360 800
rect -1308 748 -1296 800
rect -1244 748 -1232 800
rect -1180 748 -1139 800
rect -1087 748 -1075 800
rect -1023 748 -1011 800
rect -959 762 -838 800
rect -782 762 -758 818
rect -702 762 -678 818
rect -622 810 -578 818
rect -622 800 2483 810
rect -622 762 351 800
rect -959 748 351 762
rect 403 748 415 800
rect 467 748 479 800
rect 531 748 572 800
rect 624 748 636 800
rect 688 748 700 800
rect 752 748 2056 800
rect 2108 748 2120 800
rect 2172 748 2184 800
rect 2236 748 2277 800
rect 2329 748 2341 800
rect 2393 748 2405 800
rect 2457 748 2483 800
rect -1380 740 2483 748
rect 825 668 1125 690
rect 825 660 865 668
rect -1380 650 865 660
rect -1380 598 -501 650
rect -449 598 -437 650
rect -385 598 -373 650
rect -321 598 -280 650
rect -228 598 -216 650
rect -164 598 -152 650
rect -100 612 865 650
rect 921 612 945 668
rect 1001 612 1025 668
rect 1081 660 1125 668
rect 1081 650 2483 660
rect 1081 612 1206 650
rect -100 598 1206 612
rect 1258 598 1270 650
rect 1322 598 1334 650
rect 1386 598 1427 650
rect 1479 598 1491 650
rect 1543 598 1555 650
rect 1607 598 2483 650
rect -1380 590 2483 598
rect -1380 251 2483 261
rect -1380 199 204 251
rect 256 199 268 251
rect 320 199 332 251
rect 384 199 2483 251
rect -1380 191 2483 199
rect -1380 122 2483 132
rect -1380 70 -137 122
rect -85 70 -73 122
rect -21 70 -9 122
rect 43 70 1568 122
rect 1620 70 1632 122
rect 1684 70 1696 122
rect 1748 70 2483 122
rect -1380 62 2483 70
rect -1380 -276 2483 -266
rect -1380 -288 -501 -276
rect -1380 -336 -838 -288
rect -878 -344 -838 -336
rect -782 -344 -758 -288
rect -702 -344 -678 -288
rect -622 -328 -501 -288
rect -449 -328 -437 -276
rect -385 -328 -373 -276
rect -321 -328 -280 -276
rect -228 -328 -216 -276
rect -164 -328 -152 -276
rect -100 -328 1206 -276
rect 1258 -328 1270 -276
rect 1322 -328 1334 -276
rect 1386 -328 1427 -276
rect 1479 -328 1491 -276
rect 1543 -328 1555 -276
rect 1607 -328 2483 -276
rect -622 -336 2483 -328
rect -622 -344 -578 -336
rect -878 -366 -578 -344
rect -1380 -427 2483 -417
rect -1380 -479 -1354 -427
rect -1302 -479 -1290 -427
rect -1238 -479 -1226 -427
rect -1174 -479 -1133 -427
rect -1081 -479 -1069 -427
rect -1017 -479 -1005 -427
rect -953 -479 349 -427
rect 401 -479 413 -427
rect 465 -479 477 -427
rect 529 -479 570 -427
rect 622 -479 634 -427
rect 686 -479 698 -427
rect 750 -439 2056 -427
rect 750 -479 865 -439
rect -1380 -487 865 -479
rect 825 -495 865 -487
rect 921 -495 945 -439
rect 1001 -495 1025 -439
rect 1081 -479 2056 -439
rect 2108 -479 2120 -427
rect 2172 -479 2184 -427
rect 2236 -479 2277 -427
rect 2329 -479 2341 -427
rect 2393 -479 2405 -427
rect 2457 -479 2483 -427
rect 1081 -487 2483 -479
rect 1081 -495 1125 -487
rect 825 -517 1125 -495
rect -878 -559 -578 -537
rect -878 -567 -838 -559
rect -1380 -615 -838 -567
rect -782 -615 -758 -559
rect -702 -615 -678 -559
rect -622 -567 -578 -559
rect -622 -577 2483 -567
rect -622 -615 -501 -577
rect -1380 -629 -501 -615
rect -449 -629 -437 -577
rect -385 -629 -373 -577
rect -321 -629 -280 -577
rect -228 -629 -216 -577
rect -164 -629 -152 -577
rect -100 -629 1206 -577
rect 1258 -629 1270 -577
rect 1322 -629 1334 -577
rect 1386 -629 1427 -577
rect 1479 -629 1491 -577
rect 1543 -629 1555 -577
rect 1607 -629 2483 -577
rect -1380 -637 2483 -629
rect 825 -710 1125 -688
rect 825 -718 865 -710
rect -1380 -728 865 -718
rect -1380 -780 -1354 -728
rect -1302 -780 -1290 -728
rect -1238 -780 -1226 -728
rect -1174 -780 -1133 -728
rect -1081 -780 -1069 -728
rect -1017 -780 -1005 -728
rect -953 -780 349 -728
rect 401 -780 413 -728
rect 465 -780 477 -728
rect 529 -780 570 -728
rect 622 -780 634 -728
rect 686 -780 698 -728
rect 750 -766 865 -728
rect 921 -766 945 -710
rect 1001 -766 1025 -710
rect 1081 -718 1125 -710
rect 1081 -728 2483 -718
rect 1081 -766 2056 -728
rect 750 -780 2056 -766
rect 2108 -780 2120 -728
rect 2172 -780 2184 -728
rect 2236 -780 2277 -728
rect 2329 -780 2341 -728
rect 2393 -780 2405 -728
rect 2457 -780 2483 -728
rect -1380 -788 2483 -780
rect -1512 -1126 2483 -1116
rect -1512 -1178 -1503 -1126
rect -1451 -1178 -1439 -1126
rect -1387 -1178 -1375 -1126
rect -1323 -1178 207 -1126
rect 259 -1178 271 -1126
rect 323 -1178 335 -1126
rect 387 -1138 1912 -1126
rect 1964 -1138 1976 -1126
rect 387 -1178 1755 -1138
rect -1512 -1186 1755 -1178
rect 1715 -1194 1755 -1186
rect 1811 -1194 1835 -1138
rect 1891 -1178 1912 -1138
rect 1971 -1178 1976 -1138
rect 2028 -1178 2040 -1126
rect 2092 -1178 2483 -1126
rect 1891 -1194 1915 -1178
rect 1971 -1186 2483 -1178
rect 1971 -1194 2015 -1186
rect 1715 -1216 2015 -1194
rect -1380 -1266 2483 -1256
rect -1380 -1318 -134 -1266
rect -82 -1318 -70 -1266
rect -18 -1278 -6 -1266
rect 46 -1278 1568 -1266
rect 46 -1318 60 -1278
rect -1380 -1326 -20 -1318
rect -60 -1334 -20 -1326
rect 36 -1334 60 -1318
rect 116 -1334 140 -1278
rect 196 -1318 1568 -1278
rect 1620 -1318 1632 -1266
rect 1684 -1318 1696 -1266
rect 1748 -1318 2483 -1266
rect 196 -1326 2483 -1318
rect 196 -1334 240 -1326
rect -60 -1356 240 -1334
<< via2 >>
rect 1755 1602 1811 1658
rect 1835 1602 1891 1658
rect 1915 1602 1971 1658
rect -20 1462 36 1518
rect 60 1462 116 1518
rect 140 1462 196 1518
rect -838 1033 -782 1089
rect -758 1033 -702 1089
rect -678 1033 -622 1089
rect 865 883 921 939
rect 945 883 1001 939
rect 1025 883 1081 939
rect -838 762 -782 818
rect -758 762 -702 818
rect -678 762 -622 818
rect 865 612 921 668
rect 945 612 1001 668
rect 1025 612 1081 668
rect -838 -344 -782 -288
rect -758 -344 -702 -288
rect -678 -344 -622 -288
rect 865 -495 921 -439
rect 945 -495 1001 -439
rect 1025 -495 1081 -439
rect -838 -615 -782 -559
rect -758 -615 -702 -559
rect -678 -615 -622 -559
rect 865 -766 921 -710
rect 945 -766 1001 -710
rect 1025 -766 1081 -710
rect 1755 -1194 1811 -1138
rect 1835 -1194 1891 -1138
rect 1915 -1178 1964 -1138
rect 1964 -1178 1971 -1138
rect 1915 -1194 1971 -1178
rect -20 -1318 -18 -1278
rect -18 -1318 -6 -1278
rect -6 -1318 36 -1278
rect -20 -1334 36 -1318
rect 60 -1334 116 -1278
rect 140 -1334 196 -1278
<< metal3 >>
rect 1715 1658 2015 1680
rect 1715 1602 1755 1658
rect 1811 1602 1835 1658
rect 1891 1602 1915 1658
rect 1971 1602 2015 1658
rect -60 1518 240 1540
rect -60 1462 -20 1518
rect 36 1462 60 1518
rect 116 1462 140 1518
rect 196 1462 240 1518
rect -878 1089 -578 1111
rect -878 1033 -838 1089
rect -782 1033 -758 1089
rect -702 1033 -678 1089
rect -622 1033 -578 1089
rect -878 818 -578 1033
rect -878 762 -838 818
rect -782 762 -758 818
rect -702 762 -678 818
rect -622 762 -578 818
rect -878 -288 -578 762
rect -878 -344 -838 -288
rect -782 -344 -758 -288
rect -702 -344 -678 -288
rect -622 -344 -578 -288
rect -878 -559 -578 -344
rect -878 -615 -838 -559
rect -782 -615 -758 -559
rect -702 -615 -678 -559
rect -622 -615 -578 -559
rect -878 -637 -578 -615
rect -60 -1278 240 1462
rect 825 939 1125 961
rect 825 883 865 939
rect 921 883 945 939
rect 1001 883 1025 939
rect 1081 883 1125 939
rect 825 668 1125 883
rect 825 612 865 668
rect 921 612 945 668
rect 1001 612 1025 668
rect 1081 612 1125 668
rect 825 -439 1125 612
rect 825 -495 865 -439
rect 921 -495 945 -439
rect 1001 -495 1025 -439
rect 1081 -495 1125 -439
rect 825 -710 1125 -495
rect 825 -766 865 -710
rect 921 -766 945 -710
rect 1001 -766 1025 -710
rect 1081 -766 1125 -710
rect 825 -788 1125 -766
rect 1715 -1138 2015 1602
rect 1715 -1194 1755 -1138
rect 1811 -1194 1835 -1138
rect 1891 -1194 1915 -1138
rect 1971 -1194 2015 -1138
rect 1715 -1216 2015 -1194
rect -60 -1334 -20 -1278
rect 36 -1334 60 -1278
rect 116 -1334 140 -1278
rect 196 -1334 240 -1278
rect -60 -1356 240 -1334
use nfet_2series  nfet_2series_0
timestamp 1698888477
transform 1 0 -4443 0 1 390
box 2121 -118 2747 196
use nfet_2series  nfet_2series_1
timestamp 1698888477
transform 1 0 -1030 0 1 390
box 2121 -118 2747 196
use nfet_2series  nfet_2series_2
timestamp 1698888477
transform 1 0 -4443 0 -1 -1514
box 2121 -118 2747 196
use nfet_2series  nfet_2series_3
timestamp 1698888477
transform 1 0 -1885 0 -1 -1514
box 2121 -118 2747 196
use nfet_2series  nfet_2series_4
timestamp 1698888477
transform 1 0 -2739 0 -1 -1514
box 2121 -118 2747 196
use nfet_2series  nfet_2series_5
timestamp 1698888477
transform 1 0 -1032 0 -1 -1514
box 2121 -118 2747 196
use nfet_2series  nfet_2series_6
timestamp 1698888477
transform 1 0 -1890 0 1 1838
box 2121 -118 2747 196
use nfet_2series  nfet_2series_7
timestamp 1698888477
transform 1 0 -179 0 -1 -1514
box 2121 -118 2747 196
use nfet_2series  nfet_2series_8
timestamp 1698888477
transform 1 0 677 0 -1 -1514
box 2121 -118 2747 196
use nfet_2series  nfet_2series_9
timestamp 1698888477
transform 1 0 -1037 0 1 1838
box 2121 -118 2747 196
use nfet_2series  nfet_2series_10
timestamp 1698888477
transform 1 0 -184 0 1 1838
box 2121 -118 2747 196
use nfet_2series  nfet_2series_11
timestamp 1698888477
transform 1 0 -3589 0 -1 1311
box 2121 -118 2747 196
use nfet_2series  nfet_2series_12
timestamp 1698888477
transform 1 0 677 0 1 1838
box 2121 -118 2747 196
use nfet_2series  nfet_2series_13
timestamp 1698888477
transform 1 0 -2743 0 1 1838
box 2121 -118 2747 196
use nfet_2series  nfet_2series_14
timestamp 1698888477
transform 1 0 -3597 0 1 1838
box 2121 -118 2747 196
use nfet_2series  nfet_2series_15
timestamp 1698888477
transform 1 0 -177 0 -1 1311
box 2121 -118 2747 196
use nfet_2series  nfet_2series_16
timestamp 1698888477
transform 1 0 -177 0 1 390
box 2121 -118 2747 196
use nfet_2series  nfet_2series_17
timestamp 1698888477
transform 1 0 677 0 -1 1311
box 2121 -118 2747 196
use nfet_2series  nfet_2series_18
timestamp 1698888477
transform 1 0 -2736 0 1 390
box 2121 -118 2747 196
use nfet_2series  nfet_2series_19
timestamp 1698888477
transform 1 0 677 0 1 390
box 2121 -118 2747 196
use nfet_2series  nfet_2series_20
timestamp 1698888477
transform 1 0 -3589 0 1 390
box 2121 -118 2747 196
use nfet_2series  nfet_2series_21
timestamp 1698888477
transform 1 0 -3592 0 -1 -1514
box 2121 -118 2747 196
use nfet_2series  nfet_2series_22
timestamp 1698888477
transform 1 0 -1883 0 1 390
box 2121 -118 2747 196
use nfet_2series  nfet_2series_23
timestamp 1698888477
transform 1 0 -3589 0 -1 -66
box 2121 -118 2747 196
use nfet_2series  nfet_2series_24
timestamp 1698888477
transform 1 0 -3589 0 1 -988
box 2121 -118 2747 196
use nfet_2series  nfet_2series_25
timestamp 1698888477
transform 1 0 677 0 1 -988
box 2121 -118 2747 196
use nfet_2series  nfet_2series_26
timestamp 1698888477
transform 1 0 677 0 -1 -66
box 2121 -118 2747 196
use nfet_2series  nfet_2series_27
timestamp 1698888477
transform 1 0 -177 0 1 -988
box 2121 -118 2747 196
use nfet_2series  nfet_2series_28
timestamp 1698888477
transform 1 0 -177 0 -1 -66
box 2121 -118 2747 196
use nfet_2series  nfet_2series_29
timestamp 1698888477
transform 1 0 -1030 0 -1 -66
box 2121 -118 2747 196
use nfet_2series  nfet_2series_30
timestamp 1698888477
transform 1 0 -2736 0 -1 -66
box 2121 -118 2747 196
use nfet_2series  nfet_2series_31
timestamp 1698888477
transform 1 0 -1883 0 -1 -66
box 2121 -118 2747 196
use nfet_2series  nfet_2series_32
timestamp 1698888477
transform 1 0 -4443 0 -1 -66
box 2121 -118 2747 196
use nfet_2series  nfet_2series_33
timestamp 1698888477
transform 1 0 -4443 0 1 -988
box 2121 -118 2747 196
use nfet_2series  nfet_2series_34
timestamp 1698888477
transform 1 0 -1883 0 1 -988
box 2121 -118 2747 196
use nfet_2series  nfet_2series_35
timestamp 1698888477
transform 1 0 -2736 0 1 -988
box 2121 -118 2747 196
use nfet_2series  nfet_2series_36
timestamp 1698888477
transform 1 0 -1030 0 1 -988
box 2121 -118 2747 196
use nfet_2series  nfet_2series_37
timestamp 1698888477
transform 1 0 -4443 0 -1 1311
box 2121 -118 2747 196
use nfet_2series  nfet_2series_38
timestamp 1698888477
transform 1 0 -1030 0 -1 1311
box 2121 -118 2747 196
use nfet_2series  nfet_2series_39
timestamp 1698888477
transform 1 0 -2736 0 -1 1311
box 2121 -118 2747 196
use nfet_2series  nfet_2series_40
timestamp 1698888477
transform 1 0 -1883 0 -1 1311
box 2121 -118 2747 196
use nfet_2series  nfet_2series_41
timestamp 1698888477
transform 1 0 -4443 0 1 1838
box 2121 -118 2747 196
<< labels >>
flabel metal3 s -820 490 -640 600 2 FreeSans 3126 0 0 0 IREF
port 1 nsew
flabel metal3 s 20 120 150 230 2 FreeSans 3126 0 0 0 VB1
port 2 nsew
flabel metal3 s 890 110 1040 210 2 FreeSans 3126 0 0 0 VB2
port 3 nsew
flabel metal3 s 1780 90 1930 210 2 FreeSans 3126 0 0 0 VB4
port 4 nsew
flabel metal1 s 2822 -1607 3377 1617 2 FreeSans 3126 0 0 0 AVSS
port 5 nsew
<< end >>
