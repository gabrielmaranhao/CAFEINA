magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< nwell >>
rect 290 -5592 6219 6020
<< pmoshvt >>
rect 576 5589 776 5789
rect 834 5589 1034 5789
rect 1286 5589 1486 5789
rect 1544 5589 1744 5789
rect 1802 5589 2002 5789
rect 2060 5589 2260 5789
rect 2512 5589 2712 5789
rect 2770 5589 2970 5789
rect 3028 5589 3228 5789
rect 3286 5589 3486 5789
rect 3544 5589 3744 5789
rect 3802 5589 4002 5789
rect 4254 5589 4454 5789
rect 4512 5589 4712 5789
rect 4770 5589 4970 5789
rect 5028 5589 5228 5789
rect 5479 5589 5679 5789
rect 5737 5589 5937 5789
rect 576 4980 776 5180
rect 834 4980 1034 5180
rect 5479 4980 5679 5180
rect 5737 4980 5937 5180
rect 576 4085 776 4285
rect 834 4085 1034 4285
rect 5479 4085 5679 4285
rect 5737 4085 5937 4285
rect 576 3476 776 3676
rect 834 3476 1034 3676
rect 5479 3476 5679 3676
rect 5737 3476 5937 3676
rect 576 2578 776 2778
rect 834 2578 1034 2778
rect 5479 2578 5679 2778
rect 5737 2578 5937 2778
rect 576 1969 776 2169
rect 834 1969 1034 2169
rect 5479 1969 5679 2169
rect 5737 1969 5937 2169
rect 576 1209 776 1409
rect 834 1209 1034 1409
rect 5479 1209 5679 1409
rect 5737 1209 5937 1409
rect 576 600 776 800
rect 834 600 1034 800
rect 5479 600 5679 800
rect 5737 600 5937 800
rect 576 114 776 314
rect 834 114 1034 314
rect 5479 114 5679 314
rect 5737 114 5937 314
rect 576 -495 776 -295
rect 834 -495 1034 -295
rect 5479 -495 5679 -295
rect 5737 -495 5937 -295
rect 576 -972 776 -772
rect 834 -972 1034 -772
rect 5479 -972 5679 -772
rect 5737 -972 5937 -772
rect 576 -1581 776 -1381
rect 834 -1581 1034 -1381
rect 5479 -1581 5679 -1381
rect 5737 -1581 5937 -1381
rect 576 -2476 776 -2276
rect 834 -2476 1034 -2276
rect 5479 -2476 5679 -2276
rect 5737 -2476 5937 -2276
rect 576 -3085 776 -2885
rect 834 -3085 1034 -2885
rect 5479 -3085 5679 -2885
rect 5737 -3085 5937 -2885
rect 576 -3980 776 -3780
rect 834 -3980 1034 -3780
rect 5479 -3980 5679 -3780
rect 5737 -3980 5937 -3780
rect 576 -4589 776 -4389
rect 834 -4589 1034 -4389
rect 5479 -4589 5679 -4389
rect 5737 -4589 5937 -4389
rect 576 -5336 776 -5136
rect 834 -5336 1034 -5136
rect 1286 -5336 1486 -5136
rect 1544 -5336 1744 -5136
rect 1802 -5336 2002 -5136
rect 2060 -5336 2260 -5136
rect 2512 -5336 2712 -5136
rect 2770 -5336 2970 -5136
rect 3028 -5336 3228 -5136
rect 3286 -5336 3486 -5136
rect 3544 -5336 3744 -5136
rect 3802 -5336 4002 -5136
rect 4254 -5336 4454 -5136
rect 4512 -5336 4712 -5136
rect 4770 -5336 4970 -5136
rect 5028 -5336 5228 -5136
rect 5479 -5336 5679 -5136
rect 5737 -5336 5937 -5136
<< pdiff >>
rect 518 5774 576 5789
rect 518 5740 530 5774
rect 564 5740 576 5774
rect 518 5706 576 5740
rect 518 5672 530 5706
rect 564 5672 576 5706
rect 518 5638 576 5672
rect 518 5604 530 5638
rect 564 5604 576 5638
rect 518 5589 576 5604
rect 776 5774 834 5789
rect 776 5740 788 5774
rect 822 5740 834 5774
rect 776 5706 834 5740
rect 776 5672 788 5706
rect 822 5672 834 5706
rect 776 5638 834 5672
rect 776 5604 788 5638
rect 822 5604 834 5638
rect 776 5589 834 5604
rect 1034 5774 1092 5789
rect 1034 5740 1046 5774
rect 1080 5740 1092 5774
rect 1034 5706 1092 5740
rect 1034 5672 1046 5706
rect 1080 5672 1092 5706
rect 1034 5638 1092 5672
rect 1034 5604 1046 5638
rect 1080 5604 1092 5638
rect 1034 5589 1092 5604
rect 1228 5774 1286 5789
rect 1228 5740 1240 5774
rect 1274 5740 1286 5774
rect 1228 5706 1286 5740
rect 1228 5672 1240 5706
rect 1274 5672 1286 5706
rect 1228 5638 1286 5672
rect 1228 5604 1240 5638
rect 1274 5604 1286 5638
rect 1228 5589 1286 5604
rect 1486 5774 1544 5789
rect 1486 5740 1498 5774
rect 1532 5740 1544 5774
rect 1486 5706 1544 5740
rect 1486 5672 1498 5706
rect 1532 5672 1544 5706
rect 1486 5638 1544 5672
rect 1486 5604 1498 5638
rect 1532 5604 1544 5638
rect 1486 5589 1544 5604
rect 1744 5774 1802 5789
rect 1744 5740 1756 5774
rect 1790 5740 1802 5774
rect 1744 5706 1802 5740
rect 1744 5672 1756 5706
rect 1790 5672 1802 5706
rect 1744 5638 1802 5672
rect 1744 5604 1756 5638
rect 1790 5604 1802 5638
rect 1744 5589 1802 5604
rect 2002 5774 2060 5789
rect 2002 5740 2014 5774
rect 2048 5740 2060 5774
rect 2002 5706 2060 5740
rect 2002 5672 2014 5706
rect 2048 5672 2060 5706
rect 2002 5638 2060 5672
rect 2002 5604 2014 5638
rect 2048 5604 2060 5638
rect 2002 5589 2060 5604
rect 2260 5774 2318 5789
rect 2260 5740 2272 5774
rect 2306 5740 2318 5774
rect 2260 5706 2318 5740
rect 2260 5672 2272 5706
rect 2306 5672 2318 5706
rect 2260 5638 2318 5672
rect 2260 5604 2272 5638
rect 2306 5604 2318 5638
rect 2260 5589 2318 5604
rect 2454 5774 2512 5789
rect 2454 5740 2466 5774
rect 2500 5740 2512 5774
rect 2454 5706 2512 5740
rect 2454 5672 2466 5706
rect 2500 5672 2512 5706
rect 2454 5638 2512 5672
rect 2454 5604 2466 5638
rect 2500 5604 2512 5638
rect 2454 5589 2512 5604
rect 2712 5774 2770 5789
rect 2712 5740 2724 5774
rect 2758 5740 2770 5774
rect 2712 5706 2770 5740
rect 2712 5672 2724 5706
rect 2758 5672 2770 5706
rect 2712 5638 2770 5672
rect 2712 5604 2724 5638
rect 2758 5604 2770 5638
rect 2712 5589 2770 5604
rect 2970 5774 3028 5789
rect 2970 5740 2982 5774
rect 3016 5740 3028 5774
rect 2970 5706 3028 5740
rect 2970 5672 2982 5706
rect 3016 5672 3028 5706
rect 2970 5638 3028 5672
rect 2970 5604 2982 5638
rect 3016 5604 3028 5638
rect 2970 5589 3028 5604
rect 3228 5774 3286 5789
rect 3228 5740 3240 5774
rect 3274 5740 3286 5774
rect 3228 5706 3286 5740
rect 3228 5672 3240 5706
rect 3274 5672 3286 5706
rect 3228 5638 3286 5672
rect 3228 5604 3240 5638
rect 3274 5604 3286 5638
rect 3228 5589 3286 5604
rect 3486 5774 3544 5789
rect 3486 5740 3498 5774
rect 3532 5740 3544 5774
rect 3486 5706 3544 5740
rect 3486 5672 3498 5706
rect 3532 5672 3544 5706
rect 3486 5638 3544 5672
rect 3486 5604 3498 5638
rect 3532 5604 3544 5638
rect 3486 5589 3544 5604
rect 3744 5774 3802 5789
rect 3744 5740 3756 5774
rect 3790 5740 3802 5774
rect 3744 5706 3802 5740
rect 3744 5672 3756 5706
rect 3790 5672 3802 5706
rect 3744 5638 3802 5672
rect 3744 5604 3756 5638
rect 3790 5604 3802 5638
rect 3744 5589 3802 5604
rect 4002 5774 4060 5789
rect 4002 5740 4014 5774
rect 4048 5740 4060 5774
rect 4002 5706 4060 5740
rect 4002 5672 4014 5706
rect 4048 5672 4060 5706
rect 4002 5638 4060 5672
rect 4002 5604 4014 5638
rect 4048 5604 4060 5638
rect 4002 5589 4060 5604
rect 4196 5774 4254 5789
rect 4196 5740 4208 5774
rect 4242 5740 4254 5774
rect 4196 5706 4254 5740
rect 4196 5672 4208 5706
rect 4242 5672 4254 5706
rect 4196 5638 4254 5672
rect 4196 5604 4208 5638
rect 4242 5604 4254 5638
rect 4196 5589 4254 5604
rect 4454 5774 4512 5789
rect 4454 5740 4466 5774
rect 4500 5740 4512 5774
rect 4454 5706 4512 5740
rect 4454 5672 4466 5706
rect 4500 5672 4512 5706
rect 4454 5638 4512 5672
rect 4454 5604 4466 5638
rect 4500 5604 4512 5638
rect 4454 5589 4512 5604
rect 4712 5774 4770 5789
rect 4712 5740 4724 5774
rect 4758 5740 4770 5774
rect 4712 5706 4770 5740
rect 4712 5672 4724 5706
rect 4758 5672 4770 5706
rect 4712 5638 4770 5672
rect 4712 5604 4724 5638
rect 4758 5604 4770 5638
rect 4712 5589 4770 5604
rect 4970 5774 5028 5789
rect 4970 5740 4982 5774
rect 5016 5740 5028 5774
rect 4970 5706 5028 5740
rect 4970 5672 4982 5706
rect 5016 5672 5028 5706
rect 4970 5638 5028 5672
rect 4970 5604 4982 5638
rect 5016 5604 5028 5638
rect 4970 5589 5028 5604
rect 5228 5774 5286 5789
rect 5228 5740 5240 5774
rect 5274 5740 5286 5774
rect 5228 5706 5286 5740
rect 5228 5672 5240 5706
rect 5274 5672 5286 5706
rect 5228 5638 5286 5672
rect 5228 5604 5240 5638
rect 5274 5604 5286 5638
rect 5228 5589 5286 5604
rect 5421 5774 5479 5789
rect 5421 5740 5433 5774
rect 5467 5740 5479 5774
rect 5421 5706 5479 5740
rect 5421 5672 5433 5706
rect 5467 5672 5479 5706
rect 5421 5638 5479 5672
rect 5421 5604 5433 5638
rect 5467 5604 5479 5638
rect 5421 5589 5479 5604
rect 5679 5774 5737 5789
rect 5679 5740 5691 5774
rect 5725 5740 5737 5774
rect 5679 5706 5737 5740
rect 5679 5672 5691 5706
rect 5725 5672 5737 5706
rect 5679 5638 5737 5672
rect 5679 5604 5691 5638
rect 5725 5604 5737 5638
rect 5679 5589 5737 5604
rect 5937 5774 5995 5789
rect 5937 5740 5949 5774
rect 5983 5740 5995 5774
rect 5937 5706 5995 5740
rect 5937 5672 5949 5706
rect 5983 5672 5995 5706
rect 5937 5638 5995 5672
rect 5937 5604 5949 5638
rect 5983 5604 5995 5638
rect 5937 5589 5995 5604
rect 518 5165 576 5180
rect 518 5131 530 5165
rect 564 5131 576 5165
rect 518 5097 576 5131
rect 518 5063 530 5097
rect 564 5063 576 5097
rect 518 5029 576 5063
rect 518 4995 530 5029
rect 564 4995 576 5029
rect 518 4980 576 4995
rect 776 5165 834 5180
rect 776 5131 788 5165
rect 822 5131 834 5165
rect 776 5097 834 5131
rect 776 5063 788 5097
rect 822 5063 834 5097
rect 776 5029 834 5063
rect 776 4995 788 5029
rect 822 4995 834 5029
rect 776 4980 834 4995
rect 1034 5165 1092 5180
rect 1034 5131 1046 5165
rect 1080 5131 1092 5165
rect 1034 5097 1092 5131
rect 1034 5063 1046 5097
rect 1080 5063 1092 5097
rect 1034 5029 1092 5063
rect 1034 4995 1046 5029
rect 1080 4995 1092 5029
rect 1034 4980 1092 4995
rect 5421 5165 5479 5180
rect 5421 5131 5433 5165
rect 5467 5131 5479 5165
rect 5421 5097 5479 5131
rect 5421 5063 5433 5097
rect 5467 5063 5479 5097
rect 5421 5029 5479 5063
rect 5421 4995 5433 5029
rect 5467 4995 5479 5029
rect 5421 4980 5479 4995
rect 5679 5165 5737 5180
rect 5679 5131 5691 5165
rect 5725 5131 5737 5165
rect 5679 5097 5737 5131
rect 5679 5063 5691 5097
rect 5725 5063 5737 5097
rect 5679 5029 5737 5063
rect 5679 4995 5691 5029
rect 5725 4995 5737 5029
rect 5679 4980 5737 4995
rect 5937 5165 5995 5180
rect 5937 5131 5949 5165
rect 5983 5131 5995 5165
rect 5937 5097 5995 5131
rect 5937 5063 5949 5097
rect 5983 5063 5995 5097
rect 5937 5029 5995 5063
rect 5937 4995 5949 5029
rect 5983 4995 5995 5029
rect 5937 4980 5995 4995
rect 518 4270 576 4285
rect 518 4236 530 4270
rect 564 4236 576 4270
rect 518 4202 576 4236
rect 518 4168 530 4202
rect 564 4168 576 4202
rect 518 4134 576 4168
rect 518 4100 530 4134
rect 564 4100 576 4134
rect 518 4085 576 4100
rect 776 4270 834 4285
rect 776 4236 788 4270
rect 822 4236 834 4270
rect 776 4202 834 4236
rect 776 4168 788 4202
rect 822 4168 834 4202
rect 776 4134 834 4168
rect 776 4100 788 4134
rect 822 4100 834 4134
rect 776 4085 834 4100
rect 1034 4270 1092 4285
rect 1034 4236 1046 4270
rect 1080 4236 1092 4270
rect 1034 4202 1092 4236
rect 1034 4168 1046 4202
rect 1080 4168 1092 4202
rect 1034 4134 1092 4168
rect 1034 4100 1046 4134
rect 1080 4100 1092 4134
rect 1034 4085 1092 4100
rect 5421 4270 5479 4285
rect 5421 4236 5433 4270
rect 5467 4236 5479 4270
rect 5421 4202 5479 4236
rect 5421 4168 5433 4202
rect 5467 4168 5479 4202
rect 5421 4134 5479 4168
rect 5421 4100 5433 4134
rect 5467 4100 5479 4134
rect 5421 4085 5479 4100
rect 5679 4270 5737 4285
rect 5679 4236 5691 4270
rect 5725 4236 5737 4270
rect 5679 4202 5737 4236
rect 5679 4168 5691 4202
rect 5725 4168 5737 4202
rect 5679 4134 5737 4168
rect 5679 4100 5691 4134
rect 5725 4100 5737 4134
rect 5679 4085 5737 4100
rect 5937 4270 5995 4285
rect 5937 4236 5949 4270
rect 5983 4236 5995 4270
rect 5937 4202 5995 4236
rect 5937 4168 5949 4202
rect 5983 4168 5995 4202
rect 5937 4134 5995 4168
rect 5937 4100 5949 4134
rect 5983 4100 5995 4134
rect 5937 4085 5995 4100
rect 518 3661 576 3676
rect 518 3627 530 3661
rect 564 3627 576 3661
rect 518 3593 576 3627
rect 518 3559 530 3593
rect 564 3559 576 3593
rect 518 3525 576 3559
rect 518 3491 530 3525
rect 564 3491 576 3525
rect 518 3476 576 3491
rect 776 3661 834 3676
rect 776 3627 788 3661
rect 822 3627 834 3661
rect 776 3593 834 3627
rect 776 3559 788 3593
rect 822 3559 834 3593
rect 776 3525 834 3559
rect 776 3491 788 3525
rect 822 3491 834 3525
rect 776 3476 834 3491
rect 1034 3661 1092 3676
rect 1034 3627 1046 3661
rect 1080 3627 1092 3661
rect 1034 3593 1092 3627
rect 1034 3559 1046 3593
rect 1080 3559 1092 3593
rect 1034 3525 1092 3559
rect 1034 3491 1046 3525
rect 1080 3491 1092 3525
rect 1034 3476 1092 3491
rect 5421 3661 5479 3676
rect 5421 3627 5433 3661
rect 5467 3627 5479 3661
rect 5421 3593 5479 3627
rect 5421 3559 5433 3593
rect 5467 3559 5479 3593
rect 5421 3525 5479 3559
rect 5421 3491 5433 3525
rect 5467 3491 5479 3525
rect 5421 3476 5479 3491
rect 5679 3661 5737 3676
rect 5679 3627 5691 3661
rect 5725 3627 5737 3661
rect 5679 3593 5737 3627
rect 5679 3559 5691 3593
rect 5725 3559 5737 3593
rect 5679 3525 5737 3559
rect 5679 3491 5691 3525
rect 5725 3491 5737 3525
rect 5679 3476 5737 3491
rect 5937 3661 5995 3676
rect 5937 3627 5949 3661
rect 5983 3627 5995 3661
rect 5937 3593 5995 3627
rect 5937 3559 5949 3593
rect 5983 3559 5995 3593
rect 5937 3525 5995 3559
rect 5937 3491 5949 3525
rect 5983 3491 5995 3525
rect 5937 3476 5995 3491
rect 518 2763 576 2778
rect 518 2729 530 2763
rect 564 2729 576 2763
rect 518 2695 576 2729
rect 518 2661 530 2695
rect 564 2661 576 2695
rect 518 2627 576 2661
rect 518 2593 530 2627
rect 564 2593 576 2627
rect 518 2578 576 2593
rect 776 2763 834 2778
rect 776 2729 788 2763
rect 822 2729 834 2763
rect 776 2695 834 2729
rect 776 2661 788 2695
rect 822 2661 834 2695
rect 776 2627 834 2661
rect 776 2593 788 2627
rect 822 2593 834 2627
rect 776 2578 834 2593
rect 1034 2763 1092 2778
rect 1034 2729 1046 2763
rect 1080 2729 1092 2763
rect 1034 2695 1092 2729
rect 1034 2661 1046 2695
rect 1080 2661 1092 2695
rect 1034 2627 1092 2661
rect 1034 2593 1046 2627
rect 1080 2593 1092 2627
rect 1034 2578 1092 2593
rect 5421 2763 5479 2778
rect 5421 2729 5433 2763
rect 5467 2729 5479 2763
rect 5421 2695 5479 2729
rect 5421 2661 5433 2695
rect 5467 2661 5479 2695
rect 5421 2627 5479 2661
rect 5421 2593 5433 2627
rect 5467 2593 5479 2627
rect 5421 2578 5479 2593
rect 5679 2763 5737 2778
rect 5679 2729 5691 2763
rect 5725 2729 5737 2763
rect 5679 2695 5737 2729
rect 5679 2661 5691 2695
rect 5725 2661 5737 2695
rect 5679 2627 5737 2661
rect 5679 2593 5691 2627
rect 5725 2593 5737 2627
rect 5679 2578 5737 2593
rect 5937 2763 5995 2778
rect 5937 2729 5949 2763
rect 5983 2729 5995 2763
rect 5937 2695 5995 2729
rect 5937 2661 5949 2695
rect 5983 2661 5995 2695
rect 5937 2627 5995 2661
rect 5937 2593 5949 2627
rect 5983 2593 5995 2627
rect 5937 2578 5995 2593
rect 518 2154 576 2169
rect 518 2120 530 2154
rect 564 2120 576 2154
rect 518 2086 576 2120
rect 518 2052 530 2086
rect 564 2052 576 2086
rect 518 2018 576 2052
rect 518 1984 530 2018
rect 564 1984 576 2018
rect 518 1969 576 1984
rect 776 2154 834 2169
rect 776 2120 788 2154
rect 822 2120 834 2154
rect 776 2086 834 2120
rect 776 2052 788 2086
rect 822 2052 834 2086
rect 776 2018 834 2052
rect 776 1984 788 2018
rect 822 1984 834 2018
rect 776 1969 834 1984
rect 1034 2154 1092 2169
rect 1034 2120 1046 2154
rect 1080 2120 1092 2154
rect 1034 2086 1092 2120
rect 1034 2052 1046 2086
rect 1080 2052 1092 2086
rect 1034 2018 1092 2052
rect 1034 1984 1046 2018
rect 1080 1984 1092 2018
rect 1034 1969 1092 1984
rect 5421 2154 5479 2169
rect 5421 2120 5433 2154
rect 5467 2120 5479 2154
rect 5421 2086 5479 2120
rect 5421 2052 5433 2086
rect 5467 2052 5479 2086
rect 5421 2018 5479 2052
rect 5421 1984 5433 2018
rect 5467 1984 5479 2018
rect 5421 1969 5479 1984
rect 5679 2154 5737 2169
rect 5679 2120 5691 2154
rect 5725 2120 5737 2154
rect 5679 2086 5737 2120
rect 5679 2052 5691 2086
rect 5725 2052 5737 2086
rect 5679 2018 5737 2052
rect 5679 1984 5691 2018
rect 5725 1984 5737 2018
rect 5679 1969 5737 1984
rect 5937 2154 5995 2169
rect 5937 2120 5949 2154
rect 5983 2120 5995 2154
rect 5937 2086 5995 2120
rect 5937 2052 5949 2086
rect 5983 2052 5995 2086
rect 5937 2018 5995 2052
rect 5937 1984 5949 2018
rect 5983 1984 5995 2018
rect 5937 1969 5995 1984
rect 518 1394 576 1409
rect 518 1360 530 1394
rect 564 1360 576 1394
rect 518 1326 576 1360
rect 518 1292 530 1326
rect 564 1292 576 1326
rect 518 1258 576 1292
rect 518 1224 530 1258
rect 564 1224 576 1258
rect 518 1209 576 1224
rect 776 1394 834 1409
rect 776 1360 788 1394
rect 822 1360 834 1394
rect 776 1326 834 1360
rect 776 1292 788 1326
rect 822 1292 834 1326
rect 776 1258 834 1292
rect 776 1224 788 1258
rect 822 1224 834 1258
rect 776 1209 834 1224
rect 1034 1394 1092 1409
rect 1034 1360 1046 1394
rect 1080 1360 1092 1394
rect 1034 1326 1092 1360
rect 1034 1292 1046 1326
rect 1080 1292 1092 1326
rect 1034 1258 1092 1292
rect 1034 1224 1046 1258
rect 1080 1224 1092 1258
rect 1034 1209 1092 1224
rect 5421 1394 5479 1409
rect 5421 1360 5433 1394
rect 5467 1360 5479 1394
rect 5421 1326 5479 1360
rect 5421 1292 5433 1326
rect 5467 1292 5479 1326
rect 5421 1258 5479 1292
rect 5421 1224 5433 1258
rect 5467 1224 5479 1258
rect 5421 1209 5479 1224
rect 5679 1394 5737 1409
rect 5679 1360 5691 1394
rect 5725 1360 5737 1394
rect 5679 1326 5737 1360
rect 5679 1292 5691 1326
rect 5725 1292 5737 1326
rect 5679 1258 5737 1292
rect 5679 1224 5691 1258
rect 5725 1224 5737 1258
rect 5679 1209 5737 1224
rect 5937 1394 5995 1409
rect 5937 1360 5949 1394
rect 5983 1360 5995 1394
rect 5937 1326 5995 1360
rect 5937 1292 5949 1326
rect 5983 1292 5995 1326
rect 5937 1258 5995 1292
rect 5937 1224 5949 1258
rect 5983 1224 5995 1258
rect 5937 1209 5995 1224
rect 518 785 576 800
rect 518 751 530 785
rect 564 751 576 785
rect 518 717 576 751
rect 518 683 530 717
rect 564 683 576 717
rect 518 649 576 683
rect 518 615 530 649
rect 564 615 576 649
rect 518 600 576 615
rect 776 785 834 800
rect 776 751 788 785
rect 822 751 834 785
rect 776 717 834 751
rect 776 683 788 717
rect 822 683 834 717
rect 776 649 834 683
rect 776 615 788 649
rect 822 615 834 649
rect 776 600 834 615
rect 1034 785 1092 800
rect 1034 751 1046 785
rect 1080 751 1092 785
rect 1034 717 1092 751
rect 1034 683 1046 717
rect 1080 683 1092 717
rect 1034 649 1092 683
rect 1034 615 1046 649
rect 1080 615 1092 649
rect 1034 600 1092 615
rect 5421 785 5479 800
rect 5421 751 5433 785
rect 5467 751 5479 785
rect 5421 717 5479 751
rect 5421 683 5433 717
rect 5467 683 5479 717
rect 5421 649 5479 683
rect 5421 615 5433 649
rect 5467 615 5479 649
rect 5421 600 5479 615
rect 5679 785 5737 800
rect 5679 751 5691 785
rect 5725 751 5737 785
rect 5679 717 5737 751
rect 5679 683 5691 717
rect 5725 683 5737 717
rect 5679 649 5737 683
rect 5679 615 5691 649
rect 5725 615 5737 649
rect 5679 600 5737 615
rect 5937 785 5995 800
rect 5937 751 5949 785
rect 5983 751 5995 785
rect 5937 717 5995 751
rect 5937 683 5949 717
rect 5983 683 5995 717
rect 5937 649 5995 683
rect 5937 615 5949 649
rect 5983 615 5995 649
rect 5937 600 5995 615
rect 518 299 576 314
rect 518 265 530 299
rect 564 265 576 299
rect 518 231 576 265
rect 518 197 530 231
rect 564 197 576 231
rect 518 163 576 197
rect 518 129 530 163
rect 564 129 576 163
rect 518 114 576 129
rect 776 299 834 314
rect 776 265 788 299
rect 822 265 834 299
rect 776 231 834 265
rect 776 197 788 231
rect 822 197 834 231
rect 776 163 834 197
rect 776 129 788 163
rect 822 129 834 163
rect 776 114 834 129
rect 1034 299 1092 314
rect 1034 265 1046 299
rect 1080 265 1092 299
rect 1034 231 1092 265
rect 1034 197 1046 231
rect 1080 197 1092 231
rect 1034 163 1092 197
rect 1034 129 1046 163
rect 1080 129 1092 163
rect 1034 114 1092 129
rect 5421 299 5479 314
rect 5421 265 5433 299
rect 5467 265 5479 299
rect 5421 231 5479 265
rect 5421 197 5433 231
rect 5467 197 5479 231
rect 5421 163 5479 197
rect 5421 129 5433 163
rect 5467 129 5479 163
rect 5421 114 5479 129
rect 5679 299 5737 314
rect 5679 265 5691 299
rect 5725 265 5737 299
rect 5679 231 5737 265
rect 5679 197 5691 231
rect 5725 197 5737 231
rect 5679 163 5737 197
rect 5679 129 5691 163
rect 5725 129 5737 163
rect 5679 114 5737 129
rect 5937 299 5995 314
rect 5937 265 5949 299
rect 5983 265 5995 299
rect 5937 231 5995 265
rect 5937 197 5949 231
rect 5983 197 5995 231
rect 5937 163 5995 197
rect 5937 129 5949 163
rect 5983 129 5995 163
rect 5937 114 5995 129
rect 518 -310 576 -295
rect 518 -344 530 -310
rect 564 -344 576 -310
rect 518 -378 576 -344
rect 518 -412 530 -378
rect 564 -412 576 -378
rect 518 -446 576 -412
rect 518 -480 530 -446
rect 564 -480 576 -446
rect 518 -495 576 -480
rect 776 -310 834 -295
rect 776 -344 788 -310
rect 822 -344 834 -310
rect 776 -378 834 -344
rect 776 -412 788 -378
rect 822 -412 834 -378
rect 776 -446 834 -412
rect 776 -480 788 -446
rect 822 -480 834 -446
rect 776 -495 834 -480
rect 1034 -310 1092 -295
rect 1034 -344 1046 -310
rect 1080 -344 1092 -310
rect 1034 -378 1092 -344
rect 1034 -412 1046 -378
rect 1080 -412 1092 -378
rect 1034 -446 1092 -412
rect 1034 -480 1046 -446
rect 1080 -480 1092 -446
rect 1034 -495 1092 -480
rect 5421 -310 5479 -295
rect 5421 -344 5433 -310
rect 5467 -344 5479 -310
rect 5421 -378 5479 -344
rect 5421 -412 5433 -378
rect 5467 -412 5479 -378
rect 5421 -446 5479 -412
rect 5421 -480 5433 -446
rect 5467 -480 5479 -446
rect 5421 -495 5479 -480
rect 5679 -310 5737 -295
rect 5679 -344 5691 -310
rect 5725 -344 5737 -310
rect 5679 -378 5737 -344
rect 5679 -412 5691 -378
rect 5725 -412 5737 -378
rect 5679 -446 5737 -412
rect 5679 -480 5691 -446
rect 5725 -480 5737 -446
rect 5679 -495 5737 -480
rect 5937 -310 5995 -295
rect 5937 -344 5949 -310
rect 5983 -344 5995 -310
rect 5937 -378 5995 -344
rect 5937 -412 5949 -378
rect 5983 -412 5995 -378
rect 5937 -446 5995 -412
rect 5937 -480 5949 -446
rect 5983 -480 5995 -446
rect 5937 -495 5995 -480
rect 518 -787 576 -772
rect 518 -821 530 -787
rect 564 -821 576 -787
rect 518 -855 576 -821
rect 518 -889 530 -855
rect 564 -889 576 -855
rect 518 -923 576 -889
rect 518 -957 530 -923
rect 564 -957 576 -923
rect 518 -972 576 -957
rect 776 -787 834 -772
rect 776 -821 788 -787
rect 822 -821 834 -787
rect 776 -855 834 -821
rect 776 -889 788 -855
rect 822 -889 834 -855
rect 776 -923 834 -889
rect 776 -957 788 -923
rect 822 -957 834 -923
rect 776 -972 834 -957
rect 1034 -787 1092 -772
rect 1034 -821 1046 -787
rect 1080 -821 1092 -787
rect 1034 -855 1092 -821
rect 1034 -889 1046 -855
rect 1080 -889 1092 -855
rect 1034 -923 1092 -889
rect 1034 -957 1046 -923
rect 1080 -957 1092 -923
rect 1034 -972 1092 -957
rect 5421 -787 5479 -772
rect 5421 -821 5433 -787
rect 5467 -821 5479 -787
rect 5421 -855 5479 -821
rect 5421 -889 5433 -855
rect 5467 -889 5479 -855
rect 5421 -923 5479 -889
rect 5421 -957 5433 -923
rect 5467 -957 5479 -923
rect 5421 -972 5479 -957
rect 5679 -787 5737 -772
rect 5679 -821 5691 -787
rect 5725 -821 5737 -787
rect 5679 -855 5737 -821
rect 5679 -889 5691 -855
rect 5725 -889 5737 -855
rect 5679 -923 5737 -889
rect 5679 -957 5691 -923
rect 5725 -957 5737 -923
rect 5679 -972 5737 -957
rect 5937 -787 5995 -772
rect 5937 -821 5949 -787
rect 5983 -821 5995 -787
rect 5937 -855 5995 -821
rect 5937 -889 5949 -855
rect 5983 -889 5995 -855
rect 5937 -923 5995 -889
rect 5937 -957 5949 -923
rect 5983 -957 5995 -923
rect 5937 -972 5995 -957
rect 518 -1396 576 -1381
rect 518 -1430 530 -1396
rect 564 -1430 576 -1396
rect 518 -1464 576 -1430
rect 518 -1498 530 -1464
rect 564 -1498 576 -1464
rect 518 -1532 576 -1498
rect 518 -1566 530 -1532
rect 564 -1566 576 -1532
rect 518 -1581 576 -1566
rect 776 -1396 834 -1381
rect 776 -1430 788 -1396
rect 822 -1430 834 -1396
rect 776 -1464 834 -1430
rect 776 -1498 788 -1464
rect 822 -1498 834 -1464
rect 776 -1532 834 -1498
rect 776 -1566 788 -1532
rect 822 -1566 834 -1532
rect 776 -1581 834 -1566
rect 1034 -1396 1092 -1381
rect 1034 -1430 1046 -1396
rect 1080 -1430 1092 -1396
rect 1034 -1464 1092 -1430
rect 1034 -1498 1046 -1464
rect 1080 -1498 1092 -1464
rect 1034 -1532 1092 -1498
rect 1034 -1566 1046 -1532
rect 1080 -1566 1092 -1532
rect 1034 -1581 1092 -1566
rect 5421 -1396 5479 -1381
rect 5421 -1430 5433 -1396
rect 5467 -1430 5479 -1396
rect 5421 -1464 5479 -1430
rect 5421 -1498 5433 -1464
rect 5467 -1498 5479 -1464
rect 5421 -1532 5479 -1498
rect 5421 -1566 5433 -1532
rect 5467 -1566 5479 -1532
rect 5421 -1581 5479 -1566
rect 5679 -1396 5737 -1381
rect 5679 -1430 5691 -1396
rect 5725 -1430 5737 -1396
rect 5679 -1464 5737 -1430
rect 5679 -1498 5691 -1464
rect 5725 -1498 5737 -1464
rect 5679 -1532 5737 -1498
rect 5679 -1566 5691 -1532
rect 5725 -1566 5737 -1532
rect 5679 -1581 5737 -1566
rect 5937 -1396 5995 -1381
rect 5937 -1430 5949 -1396
rect 5983 -1430 5995 -1396
rect 5937 -1464 5995 -1430
rect 5937 -1498 5949 -1464
rect 5983 -1498 5995 -1464
rect 5937 -1532 5995 -1498
rect 5937 -1566 5949 -1532
rect 5983 -1566 5995 -1532
rect 5937 -1581 5995 -1566
rect 518 -2291 576 -2276
rect 518 -2325 530 -2291
rect 564 -2325 576 -2291
rect 518 -2359 576 -2325
rect 518 -2393 530 -2359
rect 564 -2393 576 -2359
rect 518 -2427 576 -2393
rect 518 -2461 530 -2427
rect 564 -2461 576 -2427
rect 518 -2476 576 -2461
rect 776 -2291 834 -2276
rect 776 -2325 788 -2291
rect 822 -2325 834 -2291
rect 776 -2359 834 -2325
rect 776 -2393 788 -2359
rect 822 -2393 834 -2359
rect 776 -2427 834 -2393
rect 776 -2461 788 -2427
rect 822 -2461 834 -2427
rect 776 -2476 834 -2461
rect 1034 -2291 1092 -2276
rect 1034 -2325 1046 -2291
rect 1080 -2325 1092 -2291
rect 1034 -2359 1092 -2325
rect 1034 -2393 1046 -2359
rect 1080 -2393 1092 -2359
rect 1034 -2427 1092 -2393
rect 1034 -2461 1046 -2427
rect 1080 -2461 1092 -2427
rect 1034 -2476 1092 -2461
rect 5421 -2291 5479 -2276
rect 5421 -2325 5433 -2291
rect 5467 -2325 5479 -2291
rect 5421 -2359 5479 -2325
rect 5421 -2393 5433 -2359
rect 5467 -2393 5479 -2359
rect 5421 -2427 5479 -2393
rect 5421 -2461 5433 -2427
rect 5467 -2461 5479 -2427
rect 5421 -2476 5479 -2461
rect 5679 -2291 5737 -2276
rect 5679 -2325 5691 -2291
rect 5725 -2325 5737 -2291
rect 5679 -2359 5737 -2325
rect 5679 -2393 5691 -2359
rect 5725 -2393 5737 -2359
rect 5679 -2427 5737 -2393
rect 5679 -2461 5691 -2427
rect 5725 -2461 5737 -2427
rect 5679 -2476 5737 -2461
rect 5937 -2291 5995 -2276
rect 5937 -2325 5949 -2291
rect 5983 -2325 5995 -2291
rect 5937 -2359 5995 -2325
rect 5937 -2393 5949 -2359
rect 5983 -2393 5995 -2359
rect 5937 -2427 5995 -2393
rect 5937 -2461 5949 -2427
rect 5983 -2461 5995 -2427
rect 5937 -2476 5995 -2461
rect 518 -2900 576 -2885
rect 518 -2934 530 -2900
rect 564 -2934 576 -2900
rect 518 -2968 576 -2934
rect 518 -3002 530 -2968
rect 564 -3002 576 -2968
rect 518 -3036 576 -3002
rect 518 -3070 530 -3036
rect 564 -3070 576 -3036
rect 518 -3085 576 -3070
rect 776 -2900 834 -2885
rect 776 -2934 788 -2900
rect 822 -2934 834 -2900
rect 776 -2968 834 -2934
rect 776 -3002 788 -2968
rect 822 -3002 834 -2968
rect 776 -3036 834 -3002
rect 776 -3070 788 -3036
rect 822 -3070 834 -3036
rect 776 -3085 834 -3070
rect 1034 -2900 1092 -2885
rect 1034 -2934 1046 -2900
rect 1080 -2934 1092 -2900
rect 1034 -2968 1092 -2934
rect 1034 -3002 1046 -2968
rect 1080 -3002 1092 -2968
rect 1034 -3036 1092 -3002
rect 1034 -3070 1046 -3036
rect 1080 -3070 1092 -3036
rect 1034 -3085 1092 -3070
rect 5421 -2900 5479 -2885
rect 5421 -2934 5433 -2900
rect 5467 -2934 5479 -2900
rect 5421 -2968 5479 -2934
rect 5421 -3002 5433 -2968
rect 5467 -3002 5479 -2968
rect 5421 -3036 5479 -3002
rect 5421 -3070 5433 -3036
rect 5467 -3070 5479 -3036
rect 5421 -3085 5479 -3070
rect 5679 -2900 5737 -2885
rect 5679 -2934 5691 -2900
rect 5725 -2934 5737 -2900
rect 5679 -2968 5737 -2934
rect 5679 -3002 5691 -2968
rect 5725 -3002 5737 -2968
rect 5679 -3036 5737 -3002
rect 5679 -3070 5691 -3036
rect 5725 -3070 5737 -3036
rect 5679 -3085 5737 -3070
rect 5937 -2900 5995 -2885
rect 5937 -2934 5949 -2900
rect 5983 -2934 5995 -2900
rect 5937 -2968 5995 -2934
rect 5937 -3002 5949 -2968
rect 5983 -3002 5995 -2968
rect 5937 -3036 5995 -3002
rect 5937 -3070 5949 -3036
rect 5983 -3070 5995 -3036
rect 5937 -3085 5995 -3070
rect 518 -3795 576 -3780
rect 518 -3829 530 -3795
rect 564 -3829 576 -3795
rect 518 -3863 576 -3829
rect 518 -3897 530 -3863
rect 564 -3897 576 -3863
rect 518 -3931 576 -3897
rect 518 -3965 530 -3931
rect 564 -3965 576 -3931
rect 518 -3980 576 -3965
rect 776 -3795 834 -3780
rect 776 -3829 788 -3795
rect 822 -3829 834 -3795
rect 776 -3863 834 -3829
rect 776 -3897 788 -3863
rect 822 -3897 834 -3863
rect 776 -3931 834 -3897
rect 776 -3965 788 -3931
rect 822 -3965 834 -3931
rect 776 -3980 834 -3965
rect 1034 -3795 1092 -3780
rect 1034 -3829 1046 -3795
rect 1080 -3829 1092 -3795
rect 1034 -3863 1092 -3829
rect 1034 -3897 1046 -3863
rect 1080 -3897 1092 -3863
rect 1034 -3931 1092 -3897
rect 1034 -3965 1046 -3931
rect 1080 -3965 1092 -3931
rect 1034 -3980 1092 -3965
rect 5421 -3795 5479 -3780
rect 5421 -3829 5433 -3795
rect 5467 -3829 5479 -3795
rect 5421 -3863 5479 -3829
rect 5421 -3897 5433 -3863
rect 5467 -3897 5479 -3863
rect 5421 -3931 5479 -3897
rect 5421 -3965 5433 -3931
rect 5467 -3965 5479 -3931
rect 5421 -3980 5479 -3965
rect 5679 -3795 5737 -3780
rect 5679 -3829 5691 -3795
rect 5725 -3829 5737 -3795
rect 5679 -3863 5737 -3829
rect 5679 -3897 5691 -3863
rect 5725 -3897 5737 -3863
rect 5679 -3931 5737 -3897
rect 5679 -3965 5691 -3931
rect 5725 -3965 5737 -3931
rect 5679 -3980 5737 -3965
rect 5937 -3795 5995 -3780
rect 5937 -3829 5949 -3795
rect 5983 -3829 5995 -3795
rect 5937 -3863 5995 -3829
rect 5937 -3897 5949 -3863
rect 5983 -3897 5995 -3863
rect 5937 -3931 5995 -3897
rect 5937 -3965 5949 -3931
rect 5983 -3965 5995 -3931
rect 5937 -3980 5995 -3965
rect 518 -4404 576 -4389
rect 518 -4438 530 -4404
rect 564 -4438 576 -4404
rect 518 -4472 576 -4438
rect 518 -4506 530 -4472
rect 564 -4506 576 -4472
rect 518 -4540 576 -4506
rect 518 -4574 530 -4540
rect 564 -4574 576 -4540
rect 518 -4589 576 -4574
rect 776 -4404 834 -4389
rect 776 -4438 788 -4404
rect 822 -4438 834 -4404
rect 776 -4472 834 -4438
rect 776 -4506 788 -4472
rect 822 -4506 834 -4472
rect 776 -4540 834 -4506
rect 776 -4574 788 -4540
rect 822 -4574 834 -4540
rect 776 -4589 834 -4574
rect 1034 -4404 1092 -4389
rect 1034 -4438 1046 -4404
rect 1080 -4438 1092 -4404
rect 1034 -4472 1092 -4438
rect 1034 -4506 1046 -4472
rect 1080 -4506 1092 -4472
rect 1034 -4540 1092 -4506
rect 1034 -4574 1046 -4540
rect 1080 -4574 1092 -4540
rect 1034 -4589 1092 -4574
rect 5421 -4404 5479 -4389
rect 5421 -4438 5433 -4404
rect 5467 -4438 5479 -4404
rect 5421 -4472 5479 -4438
rect 5421 -4506 5433 -4472
rect 5467 -4506 5479 -4472
rect 5421 -4540 5479 -4506
rect 5421 -4574 5433 -4540
rect 5467 -4574 5479 -4540
rect 5421 -4589 5479 -4574
rect 5679 -4404 5737 -4389
rect 5679 -4438 5691 -4404
rect 5725 -4438 5737 -4404
rect 5679 -4472 5737 -4438
rect 5679 -4506 5691 -4472
rect 5725 -4506 5737 -4472
rect 5679 -4540 5737 -4506
rect 5679 -4574 5691 -4540
rect 5725 -4574 5737 -4540
rect 5679 -4589 5737 -4574
rect 5937 -4404 5995 -4389
rect 5937 -4438 5949 -4404
rect 5983 -4438 5995 -4404
rect 5937 -4472 5995 -4438
rect 5937 -4506 5949 -4472
rect 5983 -4506 5995 -4472
rect 5937 -4540 5995 -4506
rect 5937 -4574 5949 -4540
rect 5983 -4574 5995 -4540
rect 5937 -4589 5995 -4574
rect 518 -5151 576 -5136
rect 518 -5185 530 -5151
rect 564 -5185 576 -5151
rect 518 -5219 576 -5185
rect 518 -5253 530 -5219
rect 564 -5253 576 -5219
rect 518 -5287 576 -5253
rect 518 -5321 530 -5287
rect 564 -5321 576 -5287
rect 518 -5336 576 -5321
rect 776 -5151 834 -5136
rect 776 -5185 788 -5151
rect 822 -5185 834 -5151
rect 776 -5219 834 -5185
rect 776 -5253 788 -5219
rect 822 -5253 834 -5219
rect 776 -5287 834 -5253
rect 776 -5321 788 -5287
rect 822 -5321 834 -5287
rect 776 -5336 834 -5321
rect 1034 -5151 1092 -5136
rect 1034 -5185 1046 -5151
rect 1080 -5185 1092 -5151
rect 1034 -5219 1092 -5185
rect 1034 -5253 1046 -5219
rect 1080 -5253 1092 -5219
rect 1034 -5287 1092 -5253
rect 1034 -5321 1046 -5287
rect 1080 -5321 1092 -5287
rect 1034 -5336 1092 -5321
rect 1228 -5151 1286 -5136
rect 1228 -5185 1240 -5151
rect 1274 -5185 1286 -5151
rect 1228 -5219 1286 -5185
rect 1228 -5253 1240 -5219
rect 1274 -5253 1286 -5219
rect 1228 -5287 1286 -5253
rect 1228 -5321 1240 -5287
rect 1274 -5321 1286 -5287
rect 1228 -5336 1286 -5321
rect 1486 -5151 1544 -5136
rect 1486 -5185 1498 -5151
rect 1532 -5185 1544 -5151
rect 1486 -5219 1544 -5185
rect 1486 -5253 1498 -5219
rect 1532 -5253 1544 -5219
rect 1486 -5287 1544 -5253
rect 1486 -5321 1498 -5287
rect 1532 -5321 1544 -5287
rect 1486 -5336 1544 -5321
rect 1744 -5151 1802 -5136
rect 1744 -5185 1756 -5151
rect 1790 -5185 1802 -5151
rect 1744 -5219 1802 -5185
rect 1744 -5253 1756 -5219
rect 1790 -5253 1802 -5219
rect 1744 -5287 1802 -5253
rect 1744 -5321 1756 -5287
rect 1790 -5321 1802 -5287
rect 1744 -5336 1802 -5321
rect 2002 -5151 2060 -5136
rect 2002 -5185 2014 -5151
rect 2048 -5185 2060 -5151
rect 2002 -5219 2060 -5185
rect 2002 -5253 2014 -5219
rect 2048 -5253 2060 -5219
rect 2002 -5287 2060 -5253
rect 2002 -5321 2014 -5287
rect 2048 -5321 2060 -5287
rect 2002 -5336 2060 -5321
rect 2260 -5151 2318 -5136
rect 2260 -5185 2272 -5151
rect 2306 -5185 2318 -5151
rect 2260 -5219 2318 -5185
rect 2260 -5253 2272 -5219
rect 2306 -5253 2318 -5219
rect 2260 -5287 2318 -5253
rect 2260 -5321 2272 -5287
rect 2306 -5321 2318 -5287
rect 2260 -5336 2318 -5321
rect 2454 -5151 2512 -5136
rect 2454 -5185 2466 -5151
rect 2500 -5185 2512 -5151
rect 2454 -5219 2512 -5185
rect 2454 -5253 2466 -5219
rect 2500 -5253 2512 -5219
rect 2454 -5287 2512 -5253
rect 2454 -5321 2466 -5287
rect 2500 -5321 2512 -5287
rect 2454 -5336 2512 -5321
rect 2712 -5151 2770 -5136
rect 2712 -5185 2724 -5151
rect 2758 -5185 2770 -5151
rect 2712 -5219 2770 -5185
rect 2712 -5253 2724 -5219
rect 2758 -5253 2770 -5219
rect 2712 -5287 2770 -5253
rect 2712 -5321 2724 -5287
rect 2758 -5321 2770 -5287
rect 2712 -5336 2770 -5321
rect 2970 -5151 3028 -5136
rect 2970 -5185 2982 -5151
rect 3016 -5185 3028 -5151
rect 2970 -5219 3028 -5185
rect 2970 -5253 2982 -5219
rect 3016 -5253 3028 -5219
rect 2970 -5287 3028 -5253
rect 2970 -5321 2982 -5287
rect 3016 -5321 3028 -5287
rect 2970 -5336 3028 -5321
rect 3228 -5151 3286 -5136
rect 3228 -5185 3240 -5151
rect 3274 -5185 3286 -5151
rect 3228 -5219 3286 -5185
rect 3228 -5253 3240 -5219
rect 3274 -5253 3286 -5219
rect 3228 -5287 3286 -5253
rect 3228 -5321 3240 -5287
rect 3274 -5321 3286 -5287
rect 3228 -5336 3286 -5321
rect 3486 -5151 3544 -5136
rect 3486 -5185 3498 -5151
rect 3532 -5185 3544 -5151
rect 3486 -5219 3544 -5185
rect 3486 -5253 3498 -5219
rect 3532 -5253 3544 -5219
rect 3486 -5287 3544 -5253
rect 3486 -5321 3498 -5287
rect 3532 -5321 3544 -5287
rect 3486 -5336 3544 -5321
rect 3744 -5151 3802 -5136
rect 3744 -5185 3756 -5151
rect 3790 -5185 3802 -5151
rect 3744 -5219 3802 -5185
rect 3744 -5253 3756 -5219
rect 3790 -5253 3802 -5219
rect 3744 -5287 3802 -5253
rect 3744 -5321 3756 -5287
rect 3790 -5321 3802 -5287
rect 3744 -5336 3802 -5321
rect 4002 -5151 4060 -5136
rect 4002 -5185 4014 -5151
rect 4048 -5185 4060 -5151
rect 4002 -5219 4060 -5185
rect 4002 -5253 4014 -5219
rect 4048 -5253 4060 -5219
rect 4002 -5287 4060 -5253
rect 4002 -5321 4014 -5287
rect 4048 -5321 4060 -5287
rect 4002 -5336 4060 -5321
rect 4196 -5151 4254 -5136
rect 4196 -5185 4208 -5151
rect 4242 -5185 4254 -5151
rect 4196 -5219 4254 -5185
rect 4196 -5253 4208 -5219
rect 4242 -5253 4254 -5219
rect 4196 -5287 4254 -5253
rect 4196 -5321 4208 -5287
rect 4242 -5321 4254 -5287
rect 4196 -5336 4254 -5321
rect 4454 -5151 4512 -5136
rect 4454 -5185 4466 -5151
rect 4500 -5185 4512 -5151
rect 4454 -5219 4512 -5185
rect 4454 -5253 4466 -5219
rect 4500 -5253 4512 -5219
rect 4454 -5287 4512 -5253
rect 4454 -5321 4466 -5287
rect 4500 -5321 4512 -5287
rect 4454 -5336 4512 -5321
rect 4712 -5151 4770 -5136
rect 4712 -5185 4724 -5151
rect 4758 -5185 4770 -5151
rect 4712 -5219 4770 -5185
rect 4712 -5253 4724 -5219
rect 4758 -5253 4770 -5219
rect 4712 -5287 4770 -5253
rect 4712 -5321 4724 -5287
rect 4758 -5321 4770 -5287
rect 4712 -5336 4770 -5321
rect 4970 -5151 5028 -5136
rect 4970 -5185 4982 -5151
rect 5016 -5185 5028 -5151
rect 4970 -5219 5028 -5185
rect 4970 -5253 4982 -5219
rect 5016 -5253 5028 -5219
rect 4970 -5287 5028 -5253
rect 4970 -5321 4982 -5287
rect 5016 -5321 5028 -5287
rect 4970 -5336 5028 -5321
rect 5228 -5151 5286 -5136
rect 5228 -5185 5240 -5151
rect 5274 -5185 5286 -5151
rect 5228 -5219 5286 -5185
rect 5228 -5253 5240 -5219
rect 5274 -5253 5286 -5219
rect 5228 -5287 5286 -5253
rect 5228 -5321 5240 -5287
rect 5274 -5321 5286 -5287
rect 5228 -5336 5286 -5321
rect 5421 -5151 5479 -5136
rect 5421 -5185 5433 -5151
rect 5467 -5185 5479 -5151
rect 5421 -5219 5479 -5185
rect 5421 -5253 5433 -5219
rect 5467 -5253 5479 -5219
rect 5421 -5287 5479 -5253
rect 5421 -5321 5433 -5287
rect 5467 -5321 5479 -5287
rect 5421 -5336 5479 -5321
rect 5679 -5151 5737 -5136
rect 5679 -5185 5691 -5151
rect 5725 -5185 5737 -5151
rect 5679 -5219 5737 -5185
rect 5679 -5253 5691 -5219
rect 5725 -5253 5737 -5219
rect 5679 -5287 5737 -5253
rect 5679 -5321 5691 -5287
rect 5725 -5321 5737 -5287
rect 5679 -5336 5737 -5321
rect 5937 -5151 5995 -5136
rect 5937 -5185 5949 -5151
rect 5983 -5185 5995 -5151
rect 5937 -5219 5995 -5185
rect 5937 -5253 5949 -5219
rect 5983 -5253 5995 -5219
rect 5937 -5287 5995 -5253
rect 5937 -5321 5949 -5287
rect 5983 -5321 5995 -5287
rect 5937 -5336 5995 -5321
<< pdiffc >>
rect 530 5740 564 5774
rect 530 5672 564 5706
rect 530 5604 564 5638
rect 788 5740 822 5774
rect 788 5672 822 5706
rect 788 5604 822 5638
rect 1046 5740 1080 5774
rect 1046 5672 1080 5706
rect 1046 5604 1080 5638
rect 1240 5740 1274 5774
rect 1240 5672 1274 5706
rect 1240 5604 1274 5638
rect 1498 5740 1532 5774
rect 1498 5672 1532 5706
rect 1498 5604 1532 5638
rect 1756 5740 1790 5774
rect 1756 5672 1790 5706
rect 1756 5604 1790 5638
rect 2014 5740 2048 5774
rect 2014 5672 2048 5706
rect 2014 5604 2048 5638
rect 2272 5740 2306 5774
rect 2272 5672 2306 5706
rect 2272 5604 2306 5638
rect 2466 5740 2500 5774
rect 2466 5672 2500 5706
rect 2466 5604 2500 5638
rect 2724 5740 2758 5774
rect 2724 5672 2758 5706
rect 2724 5604 2758 5638
rect 2982 5740 3016 5774
rect 2982 5672 3016 5706
rect 2982 5604 3016 5638
rect 3240 5740 3274 5774
rect 3240 5672 3274 5706
rect 3240 5604 3274 5638
rect 3498 5740 3532 5774
rect 3498 5672 3532 5706
rect 3498 5604 3532 5638
rect 3756 5740 3790 5774
rect 3756 5672 3790 5706
rect 3756 5604 3790 5638
rect 4014 5740 4048 5774
rect 4014 5672 4048 5706
rect 4014 5604 4048 5638
rect 4208 5740 4242 5774
rect 4208 5672 4242 5706
rect 4208 5604 4242 5638
rect 4466 5740 4500 5774
rect 4466 5672 4500 5706
rect 4466 5604 4500 5638
rect 4724 5740 4758 5774
rect 4724 5672 4758 5706
rect 4724 5604 4758 5638
rect 4982 5740 5016 5774
rect 4982 5672 5016 5706
rect 4982 5604 5016 5638
rect 5240 5740 5274 5774
rect 5240 5672 5274 5706
rect 5240 5604 5274 5638
rect 5433 5740 5467 5774
rect 5433 5672 5467 5706
rect 5433 5604 5467 5638
rect 5691 5740 5725 5774
rect 5691 5672 5725 5706
rect 5691 5604 5725 5638
rect 5949 5740 5983 5774
rect 5949 5672 5983 5706
rect 5949 5604 5983 5638
rect 530 5131 564 5165
rect 530 5063 564 5097
rect 530 4995 564 5029
rect 788 5131 822 5165
rect 788 5063 822 5097
rect 788 4995 822 5029
rect 1046 5131 1080 5165
rect 1046 5063 1080 5097
rect 1046 4995 1080 5029
rect 5433 5131 5467 5165
rect 5433 5063 5467 5097
rect 5433 4995 5467 5029
rect 5691 5131 5725 5165
rect 5691 5063 5725 5097
rect 5691 4995 5725 5029
rect 5949 5131 5983 5165
rect 5949 5063 5983 5097
rect 5949 4995 5983 5029
rect 530 4236 564 4270
rect 530 4168 564 4202
rect 530 4100 564 4134
rect 788 4236 822 4270
rect 788 4168 822 4202
rect 788 4100 822 4134
rect 1046 4236 1080 4270
rect 1046 4168 1080 4202
rect 1046 4100 1080 4134
rect 5433 4236 5467 4270
rect 5433 4168 5467 4202
rect 5433 4100 5467 4134
rect 5691 4236 5725 4270
rect 5691 4168 5725 4202
rect 5691 4100 5725 4134
rect 5949 4236 5983 4270
rect 5949 4168 5983 4202
rect 5949 4100 5983 4134
rect 530 3627 564 3661
rect 530 3559 564 3593
rect 530 3491 564 3525
rect 788 3627 822 3661
rect 788 3559 822 3593
rect 788 3491 822 3525
rect 1046 3627 1080 3661
rect 1046 3559 1080 3593
rect 1046 3491 1080 3525
rect 5433 3627 5467 3661
rect 5433 3559 5467 3593
rect 5433 3491 5467 3525
rect 5691 3627 5725 3661
rect 5691 3559 5725 3593
rect 5691 3491 5725 3525
rect 5949 3627 5983 3661
rect 5949 3559 5983 3593
rect 5949 3491 5983 3525
rect 530 2729 564 2763
rect 530 2661 564 2695
rect 530 2593 564 2627
rect 788 2729 822 2763
rect 788 2661 822 2695
rect 788 2593 822 2627
rect 1046 2729 1080 2763
rect 1046 2661 1080 2695
rect 1046 2593 1080 2627
rect 5433 2729 5467 2763
rect 5433 2661 5467 2695
rect 5433 2593 5467 2627
rect 5691 2729 5725 2763
rect 5691 2661 5725 2695
rect 5691 2593 5725 2627
rect 5949 2729 5983 2763
rect 5949 2661 5983 2695
rect 5949 2593 5983 2627
rect 530 2120 564 2154
rect 530 2052 564 2086
rect 530 1984 564 2018
rect 788 2120 822 2154
rect 788 2052 822 2086
rect 788 1984 822 2018
rect 1046 2120 1080 2154
rect 1046 2052 1080 2086
rect 1046 1984 1080 2018
rect 5433 2120 5467 2154
rect 5433 2052 5467 2086
rect 5433 1984 5467 2018
rect 5691 2120 5725 2154
rect 5691 2052 5725 2086
rect 5691 1984 5725 2018
rect 5949 2120 5983 2154
rect 5949 2052 5983 2086
rect 5949 1984 5983 2018
rect 530 1360 564 1394
rect 530 1292 564 1326
rect 530 1224 564 1258
rect 788 1360 822 1394
rect 788 1292 822 1326
rect 788 1224 822 1258
rect 1046 1360 1080 1394
rect 1046 1292 1080 1326
rect 1046 1224 1080 1258
rect 5433 1360 5467 1394
rect 5433 1292 5467 1326
rect 5433 1224 5467 1258
rect 5691 1360 5725 1394
rect 5691 1292 5725 1326
rect 5691 1224 5725 1258
rect 5949 1360 5983 1394
rect 5949 1292 5983 1326
rect 5949 1224 5983 1258
rect 530 751 564 785
rect 530 683 564 717
rect 530 615 564 649
rect 788 751 822 785
rect 788 683 822 717
rect 788 615 822 649
rect 1046 751 1080 785
rect 1046 683 1080 717
rect 1046 615 1080 649
rect 5433 751 5467 785
rect 5433 683 5467 717
rect 5433 615 5467 649
rect 5691 751 5725 785
rect 5691 683 5725 717
rect 5691 615 5725 649
rect 5949 751 5983 785
rect 5949 683 5983 717
rect 5949 615 5983 649
rect 530 265 564 299
rect 530 197 564 231
rect 530 129 564 163
rect 788 265 822 299
rect 788 197 822 231
rect 788 129 822 163
rect 1046 265 1080 299
rect 1046 197 1080 231
rect 1046 129 1080 163
rect 5433 265 5467 299
rect 5433 197 5467 231
rect 5433 129 5467 163
rect 5691 265 5725 299
rect 5691 197 5725 231
rect 5691 129 5725 163
rect 5949 265 5983 299
rect 5949 197 5983 231
rect 5949 129 5983 163
rect 530 -344 564 -310
rect 530 -412 564 -378
rect 530 -480 564 -446
rect 788 -344 822 -310
rect 788 -412 822 -378
rect 788 -480 822 -446
rect 1046 -344 1080 -310
rect 1046 -412 1080 -378
rect 1046 -480 1080 -446
rect 5433 -344 5467 -310
rect 5433 -412 5467 -378
rect 5433 -480 5467 -446
rect 5691 -344 5725 -310
rect 5691 -412 5725 -378
rect 5691 -480 5725 -446
rect 5949 -344 5983 -310
rect 5949 -412 5983 -378
rect 5949 -480 5983 -446
rect 530 -821 564 -787
rect 530 -889 564 -855
rect 530 -957 564 -923
rect 788 -821 822 -787
rect 788 -889 822 -855
rect 788 -957 822 -923
rect 1046 -821 1080 -787
rect 1046 -889 1080 -855
rect 1046 -957 1080 -923
rect 5433 -821 5467 -787
rect 5433 -889 5467 -855
rect 5433 -957 5467 -923
rect 5691 -821 5725 -787
rect 5691 -889 5725 -855
rect 5691 -957 5725 -923
rect 5949 -821 5983 -787
rect 5949 -889 5983 -855
rect 5949 -957 5983 -923
rect 530 -1430 564 -1396
rect 530 -1498 564 -1464
rect 530 -1566 564 -1532
rect 788 -1430 822 -1396
rect 788 -1498 822 -1464
rect 788 -1566 822 -1532
rect 1046 -1430 1080 -1396
rect 1046 -1498 1080 -1464
rect 1046 -1566 1080 -1532
rect 5433 -1430 5467 -1396
rect 5433 -1498 5467 -1464
rect 5433 -1566 5467 -1532
rect 5691 -1430 5725 -1396
rect 5691 -1498 5725 -1464
rect 5691 -1566 5725 -1532
rect 5949 -1430 5983 -1396
rect 5949 -1498 5983 -1464
rect 5949 -1566 5983 -1532
rect 530 -2325 564 -2291
rect 530 -2393 564 -2359
rect 530 -2461 564 -2427
rect 788 -2325 822 -2291
rect 788 -2393 822 -2359
rect 788 -2461 822 -2427
rect 1046 -2325 1080 -2291
rect 1046 -2393 1080 -2359
rect 1046 -2461 1080 -2427
rect 5433 -2325 5467 -2291
rect 5433 -2393 5467 -2359
rect 5433 -2461 5467 -2427
rect 5691 -2325 5725 -2291
rect 5691 -2393 5725 -2359
rect 5691 -2461 5725 -2427
rect 5949 -2325 5983 -2291
rect 5949 -2393 5983 -2359
rect 5949 -2461 5983 -2427
rect 530 -2934 564 -2900
rect 530 -3002 564 -2968
rect 530 -3070 564 -3036
rect 788 -2934 822 -2900
rect 788 -3002 822 -2968
rect 788 -3070 822 -3036
rect 1046 -2934 1080 -2900
rect 1046 -3002 1080 -2968
rect 1046 -3070 1080 -3036
rect 5433 -2934 5467 -2900
rect 5433 -3002 5467 -2968
rect 5433 -3070 5467 -3036
rect 5691 -2934 5725 -2900
rect 5691 -3002 5725 -2968
rect 5691 -3070 5725 -3036
rect 5949 -2934 5983 -2900
rect 5949 -3002 5983 -2968
rect 5949 -3070 5983 -3036
rect 530 -3829 564 -3795
rect 530 -3897 564 -3863
rect 530 -3965 564 -3931
rect 788 -3829 822 -3795
rect 788 -3897 822 -3863
rect 788 -3965 822 -3931
rect 1046 -3829 1080 -3795
rect 1046 -3897 1080 -3863
rect 1046 -3965 1080 -3931
rect 5433 -3829 5467 -3795
rect 5433 -3897 5467 -3863
rect 5433 -3965 5467 -3931
rect 5691 -3829 5725 -3795
rect 5691 -3897 5725 -3863
rect 5691 -3965 5725 -3931
rect 5949 -3829 5983 -3795
rect 5949 -3897 5983 -3863
rect 5949 -3965 5983 -3931
rect 530 -4438 564 -4404
rect 530 -4506 564 -4472
rect 530 -4574 564 -4540
rect 788 -4438 822 -4404
rect 788 -4506 822 -4472
rect 788 -4574 822 -4540
rect 1046 -4438 1080 -4404
rect 1046 -4506 1080 -4472
rect 1046 -4574 1080 -4540
rect 5433 -4438 5467 -4404
rect 5433 -4506 5467 -4472
rect 5433 -4574 5467 -4540
rect 5691 -4438 5725 -4404
rect 5691 -4506 5725 -4472
rect 5691 -4574 5725 -4540
rect 5949 -4438 5983 -4404
rect 5949 -4506 5983 -4472
rect 5949 -4574 5983 -4540
rect 530 -5185 564 -5151
rect 530 -5253 564 -5219
rect 530 -5321 564 -5287
rect 788 -5185 822 -5151
rect 788 -5253 822 -5219
rect 788 -5321 822 -5287
rect 1046 -5185 1080 -5151
rect 1046 -5253 1080 -5219
rect 1046 -5321 1080 -5287
rect 1240 -5185 1274 -5151
rect 1240 -5253 1274 -5219
rect 1240 -5321 1274 -5287
rect 1498 -5185 1532 -5151
rect 1498 -5253 1532 -5219
rect 1498 -5321 1532 -5287
rect 1756 -5185 1790 -5151
rect 1756 -5253 1790 -5219
rect 1756 -5321 1790 -5287
rect 2014 -5185 2048 -5151
rect 2014 -5253 2048 -5219
rect 2014 -5321 2048 -5287
rect 2272 -5185 2306 -5151
rect 2272 -5253 2306 -5219
rect 2272 -5321 2306 -5287
rect 2466 -5185 2500 -5151
rect 2466 -5253 2500 -5219
rect 2466 -5321 2500 -5287
rect 2724 -5185 2758 -5151
rect 2724 -5253 2758 -5219
rect 2724 -5321 2758 -5287
rect 2982 -5185 3016 -5151
rect 2982 -5253 3016 -5219
rect 2982 -5321 3016 -5287
rect 3240 -5185 3274 -5151
rect 3240 -5253 3274 -5219
rect 3240 -5321 3274 -5287
rect 3498 -5185 3532 -5151
rect 3498 -5253 3532 -5219
rect 3498 -5321 3532 -5287
rect 3756 -5185 3790 -5151
rect 3756 -5253 3790 -5219
rect 3756 -5321 3790 -5287
rect 4014 -5185 4048 -5151
rect 4014 -5253 4048 -5219
rect 4014 -5321 4048 -5287
rect 4208 -5185 4242 -5151
rect 4208 -5253 4242 -5219
rect 4208 -5321 4242 -5287
rect 4466 -5185 4500 -5151
rect 4466 -5253 4500 -5219
rect 4466 -5321 4500 -5287
rect 4724 -5185 4758 -5151
rect 4724 -5253 4758 -5219
rect 4724 -5321 4758 -5287
rect 4982 -5185 5016 -5151
rect 4982 -5253 5016 -5219
rect 4982 -5321 5016 -5287
rect 5240 -5185 5274 -5151
rect 5240 -5253 5274 -5219
rect 5240 -5321 5274 -5287
rect 5433 -5185 5467 -5151
rect 5433 -5253 5467 -5219
rect 5433 -5321 5467 -5287
rect 5691 -5185 5725 -5151
rect 5691 -5253 5725 -5219
rect 5691 -5321 5725 -5287
rect 5949 -5185 5983 -5151
rect 5949 -5253 5983 -5219
rect 5949 -5321 5983 -5287
<< nsubdiff >>
rect 340 5922 461 5956
rect 495 5922 529 5956
rect 563 5922 597 5956
rect 631 5922 665 5956
rect 699 5922 733 5956
rect 767 5922 801 5956
rect 835 5922 869 5956
rect 903 5922 937 5956
rect 971 5922 1005 5956
rect 1039 5922 1073 5956
rect 1107 5922 1141 5956
rect 1175 5922 1209 5956
rect 1243 5922 1277 5956
rect 1311 5922 1345 5956
rect 1379 5922 1413 5956
rect 1447 5922 1481 5956
rect 1515 5922 1549 5956
rect 1583 5922 1617 5956
rect 1651 5922 1685 5956
rect 1719 5922 1753 5956
rect 1787 5922 1821 5956
rect 1855 5922 1889 5956
rect 1923 5922 1957 5956
rect 1991 5922 2025 5956
rect 2059 5922 2093 5956
rect 2127 5922 2161 5956
rect 2195 5922 2229 5956
rect 2263 5922 2297 5956
rect 2331 5922 2365 5956
rect 2399 5922 2433 5956
rect 2467 5922 2501 5956
rect 2535 5922 2569 5956
rect 2603 5922 2637 5956
rect 2671 5922 2705 5956
rect 2739 5922 2773 5956
rect 2807 5922 2841 5956
rect 2875 5922 2909 5956
rect 2943 5922 2977 5956
rect 3011 5922 3045 5956
rect 3079 5922 3113 5956
rect 3147 5922 3181 5956
rect 3215 5922 3249 5956
rect 3283 5922 3317 5956
rect 3351 5922 3385 5956
rect 3419 5922 3453 5956
rect 3487 5922 3521 5956
rect 3555 5922 3589 5956
rect 3623 5922 3657 5956
rect 3691 5922 3725 5956
rect 3759 5922 3793 5956
rect 3827 5922 3861 5956
rect 3895 5922 3929 5956
rect 3963 5922 3997 5956
rect 4031 5922 4065 5956
rect 4099 5922 4133 5956
rect 4167 5922 4201 5956
rect 4235 5922 4269 5956
rect 4303 5922 4337 5956
rect 4371 5922 4405 5956
rect 4439 5922 4473 5956
rect 4507 5922 4541 5956
rect 4575 5922 4609 5956
rect 4643 5922 4677 5956
rect 4711 5922 4745 5956
rect 4779 5922 4813 5956
rect 4847 5922 4881 5956
rect 4915 5922 4949 5956
rect 4983 5922 5017 5956
rect 5051 5922 5085 5956
rect 5119 5922 5153 5956
rect 5187 5922 5221 5956
rect 5255 5922 5289 5956
rect 5323 5922 5357 5956
rect 5391 5922 5425 5956
rect 5459 5922 5493 5956
rect 5527 5922 5561 5956
rect 5595 5922 5629 5956
rect 5663 5922 5697 5956
rect 5731 5922 5765 5956
rect 5799 5922 5833 5956
rect 5867 5922 5901 5956
rect 5935 5922 5969 5956
rect 6003 5922 6166 5956
rect 340 5795 374 5922
rect 6132 5795 6166 5922
rect 340 5727 374 5761
rect 340 5659 374 5693
rect 340 5591 374 5625
rect 6132 5727 6166 5761
rect 6132 5659 6166 5693
rect 6132 5591 6166 5625
rect 340 5523 374 5557
rect 6132 5523 6166 5557
rect 340 5455 374 5489
rect 340 5387 374 5421
rect 340 5319 374 5353
rect 340 5251 374 5285
rect 6132 5455 6166 5489
rect 6132 5387 6166 5421
rect 6132 5319 6166 5353
rect 340 5183 374 5217
rect 6132 5251 6166 5285
rect 6132 5183 6166 5217
rect 340 5115 374 5149
rect 340 5047 374 5081
rect 340 4979 374 5013
rect 6132 5115 6166 5149
rect 6132 5047 6166 5081
rect 6132 4979 6166 5013
rect 340 4911 374 4945
rect 340 4843 374 4877
rect 340 4775 374 4809
rect 340 4707 374 4741
rect 340 4639 374 4673
rect 340 4571 374 4605
rect 340 4503 374 4537
rect 340 4435 374 4469
rect 340 4367 374 4401
rect 340 4299 374 4333
rect 6132 4911 6166 4945
rect 6132 4843 6166 4877
rect 6132 4775 6166 4809
rect 6132 4707 6166 4741
rect 6132 4639 6166 4673
rect 6132 4571 6166 4605
rect 6132 4503 6166 4537
rect 6132 4435 6166 4469
rect 6132 4367 6166 4401
rect 6132 4299 6166 4333
rect 340 4231 374 4265
rect 340 4163 374 4197
rect 340 4095 374 4129
rect 6132 4231 6166 4265
rect 6132 4163 6166 4197
rect 6132 4095 6166 4129
rect 340 4027 374 4061
rect 340 3959 374 3993
rect 6132 4027 6166 4061
rect 340 3891 374 3925
rect 340 3823 374 3857
rect 340 3755 374 3789
rect 6132 3959 6166 3993
rect 6132 3891 6166 3925
rect 6132 3823 6166 3857
rect 340 3687 374 3721
rect 6132 3755 6166 3789
rect 6132 3687 6166 3721
rect 340 3619 374 3653
rect 340 3551 374 3585
rect 340 3483 374 3517
rect 6132 3619 6166 3653
rect 6132 3551 6166 3585
rect 6132 3483 6166 3517
rect 340 3415 374 3449
rect 340 3347 374 3381
rect 340 3279 374 3313
rect 340 3211 374 3245
rect 340 3143 374 3177
rect 340 3075 374 3109
rect 340 3007 374 3041
rect 340 2939 374 2973
rect 340 2871 374 2905
rect 340 2803 374 2837
rect 6132 3415 6166 3449
rect 6132 3347 6166 3381
rect 6132 3279 6166 3313
rect 6132 3211 6166 3245
rect 6132 3143 6166 3177
rect 6132 3075 6166 3109
rect 6132 3007 6166 3041
rect 6132 2939 6166 2973
rect 6132 2871 6166 2905
rect 6132 2803 6166 2837
rect 340 2735 374 2769
rect 340 2667 374 2701
rect 340 2599 374 2633
rect 6132 2735 6166 2769
rect 6132 2667 6166 2701
rect 6132 2599 6166 2633
rect 340 2531 374 2565
rect 340 2463 374 2497
rect 6132 2531 6166 2565
rect 340 2395 374 2429
rect 340 2327 374 2361
rect 340 2259 374 2293
rect 6132 2463 6166 2497
rect 6132 2395 6166 2429
rect 6132 2327 6166 2361
rect 340 2191 374 2225
rect 6132 2259 6166 2293
rect 6132 2191 6166 2225
rect 340 2123 374 2157
rect 340 1882 374 2089
rect 6132 2123 6166 2157
rect 340 1814 374 1848
rect 340 1746 374 1780
rect 340 1678 374 1712
rect 340 1610 374 1644
rect 340 1570 374 1576
rect 6132 1882 6166 2089
rect 6132 1814 6166 1848
rect 6132 1746 6166 1780
rect 6132 1678 6166 1712
rect 6132 1610 6166 1644
rect 6132 1570 6166 1576
rect 340 1542 6166 1570
rect 374 1536 6132 1542
rect 340 1474 374 1508
rect 340 1406 374 1440
rect 6132 1474 6166 1508
rect 340 1338 374 1372
rect 340 1270 374 1304
rect 340 1202 374 1236
rect 6132 1406 6166 1440
rect 6132 1338 6166 1372
rect 6132 1270 6166 1304
rect 340 1134 374 1168
rect 6132 1202 6166 1236
rect 6132 1134 6166 1168
rect 340 1066 374 1100
rect 340 998 374 1032
rect 340 930 374 964
rect 6132 1066 6166 1100
rect 6132 998 6166 1032
rect 6132 930 6166 964
rect 340 862 374 896
rect 340 794 374 828
rect 6132 862 6166 896
rect 340 726 374 760
rect 340 658 374 692
rect 340 590 374 624
rect 6132 794 6166 828
rect 6132 726 6166 760
rect 6132 658 6166 692
rect 6132 590 6166 624
rect 340 522 374 556
rect 340 454 374 488
rect 340 386 374 420
rect 340 318 374 352
rect 6132 522 6166 556
rect 6132 454 6166 488
rect 6132 386 6166 420
rect 6132 318 6166 352
rect 340 250 374 284
rect 340 182 374 216
rect 340 114 374 148
rect 6132 250 6166 284
rect 6132 182 6166 216
rect 6132 114 6166 148
rect 340 46 374 80
rect 6132 46 6166 80
rect 340 -22 374 12
rect 340 -90 374 -56
rect 340 -158 374 -124
rect 340 -226 374 -192
rect 6132 -22 6166 12
rect 6132 -90 6166 -56
rect 6132 -158 6166 -124
rect 340 -294 374 -260
rect 6132 -226 6166 -192
rect 6132 -294 6166 -260
rect 340 -362 374 -328
rect 340 -430 374 -396
rect 340 -498 374 -464
rect 6132 -362 6166 -328
rect 6132 -430 6166 -396
rect 6132 -498 6166 -464
rect 340 -566 374 -532
rect 340 -634 374 -600
rect 340 -702 374 -668
rect 340 -770 374 -736
rect 6132 -566 6166 -532
rect 6132 -634 6166 -600
rect 6132 -702 6166 -668
rect 6132 -770 6166 -736
rect 340 -838 374 -804
rect 340 -906 374 -872
rect 340 -974 374 -940
rect 6132 -838 6166 -804
rect 6132 -906 6166 -872
rect 340 -1042 374 -1008
rect 6132 -974 6166 -940
rect 6132 -1042 6166 -1008
rect 340 -1110 374 -1076
rect 340 -1154 374 -1144
rect 6132 -1110 6166 -1076
rect 6132 -1154 6166 -1144
rect 340 -1178 6166 -1154
rect 374 -1188 6132 -1178
rect 340 -1246 374 -1212
rect 340 -1314 374 -1280
rect 6132 -1246 6166 -1212
rect 340 -1382 374 -1348
rect 6132 -1314 6166 -1280
rect 340 -1450 374 -1416
rect 340 -1518 374 -1484
rect 340 -1586 374 -1552
rect 6132 -1382 6166 -1348
rect 6132 -1450 6166 -1416
rect 6132 -1518 6166 -1484
rect 6132 -1586 6166 -1552
rect 340 -1654 374 -1620
rect 340 -1722 374 -1688
rect 340 -1790 374 -1756
rect 340 -1858 374 -1824
rect 340 -1926 374 -1892
rect 340 -1994 374 -1960
rect 340 -2062 374 -2028
rect 340 -2130 374 -2096
rect 340 -2198 374 -2164
rect 340 -2266 374 -2232
rect 6132 -1654 6166 -1620
rect 6132 -1722 6166 -1688
rect 6132 -1790 6166 -1756
rect 6132 -1858 6166 -1824
rect 6132 -1926 6166 -1892
rect 6132 -1994 6166 -1960
rect 6132 -2062 6166 -2028
rect 6132 -2130 6166 -2096
rect 6132 -2198 6166 -2164
rect 6132 -2266 6166 -2232
rect 340 -2334 374 -2300
rect 340 -2402 374 -2368
rect 340 -2470 374 -2436
rect 6132 -2334 6166 -2300
rect 6132 -2402 6166 -2368
rect 6132 -2470 6166 -2436
rect 340 -2538 374 -2504
rect 340 -2606 374 -2572
rect 6132 -2538 6166 -2504
rect 340 -2674 374 -2640
rect 340 -2742 374 -2708
rect 340 -2810 374 -2776
rect 6132 -2606 6166 -2572
rect 6132 -2674 6166 -2640
rect 6132 -2742 6166 -2708
rect 340 -2878 374 -2844
rect 6132 -2810 6166 -2776
rect 6132 -2878 6166 -2844
rect 340 -2946 374 -2912
rect 340 -3014 374 -2980
rect 340 -3082 374 -3048
rect 6132 -2946 6166 -2912
rect 6132 -3014 6166 -2980
rect 6132 -3082 6166 -3048
rect 340 -3150 374 -3116
rect 340 -3218 374 -3184
rect 340 -3286 374 -3252
rect 340 -3354 374 -3320
rect 340 -3422 374 -3388
rect 340 -3490 374 -3456
rect 340 -3558 374 -3524
rect 340 -3626 374 -3592
rect 340 -3694 374 -3660
rect 340 -3762 374 -3728
rect 6132 -3150 6166 -3116
rect 6132 -3218 6166 -3184
rect 6132 -3286 6166 -3252
rect 6132 -3354 6166 -3320
rect 6132 -3422 6166 -3388
rect 6132 -3490 6166 -3456
rect 6132 -3558 6166 -3524
rect 6132 -3626 6166 -3592
rect 6132 -3694 6166 -3660
rect 6132 -3762 6166 -3728
rect 340 -3830 374 -3796
rect 340 -3898 374 -3864
rect 340 -3966 374 -3932
rect 6132 -3830 6166 -3796
rect 6132 -3898 6166 -3864
rect 6132 -3966 6166 -3932
rect 340 -4034 374 -4000
rect 340 -4102 374 -4068
rect 6132 -4034 6166 -4000
rect 340 -4170 374 -4136
rect 340 -4238 374 -4204
rect 340 -4306 374 -4272
rect 6132 -4102 6166 -4068
rect 6132 -4170 6166 -4136
rect 6132 -4238 6166 -4204
rect 340 -4374 374 -4340
rect 6132 -4306 6166 -4272
rect 6132 -4374 6166 -4340
rect 340 -4442 374 -4408
rect 340 -4510 374 -4476
rect 340 -4578 374 -4544
rect 6132 -4442 6166 -4408
rect 6132 -4510 6166 -4476
rect 6132 -4578 6166 -4544
rect 340 -4646 374 -4612
rect 340 -4714 374 -4680
rect 340 -4782 374 -4748
rect 340 -4850 374 -4816
rect 340 -4918 374 -4884
rect 340 -4986 374 -4952
rect 340 -5054 374 -5020
rect 340 -5122 374 -5088
rect 6132 -4646 6166 -4612
rect 6132 -4714 6166 -4680
rect 6132 -4782 6166 -4748
rect 6132 -4850 6166 -4816
rect 6132 -4918 6166 -4884
rect 6132 -4986 6166 -4952
rect 6132 -5054 6166 -5020
rect 6132 -5122 6166 -5088
rect 340 -5190 374 -5156
rect 340 -5258 374 -5224
rect 340 -5326 374 -5292
rect 6132 -5190 6166 -5156
rect 6132 -5258 6166 -5224
rect 6132 -5326 6166 -5292
rect 340 -5506 374 -5360
rect 6132 -5506 6166 -5360
rect 340 -5540 461 -5506
rect 495 -5540 529 -5506
rect 563 -5540 597 -5506
rect 631 -5540 665 -5506
rect 699 -5540 733 -5506
rect 767 -5540 801 -5506
rect 835 -5540 869 -5506
rect 903 -5540 937 -5506
rect 971 -5540 1005 -5506
rect 1039 -5540 1073 -5506
rect 1107 -5540 1141 -5506
rect 1175 -5540 1209 -5506
rect 1243 -5540 1277 -5506
rect 1311 -5540 1345 -5506
rect 1379 -5540 1413 -5506
rect 1447 -5540 1481 -5506
rect 1515 -5540 1549 -5506
rect 1583 -5540 1617 -5506
rect 1651 -5540 1685 -5506
rect 1719 -5540 1753 -5506
rect 1787 -5540 1821 -5506
rect 1855 -5540 1889 -5506
rect 1923 -5540 1957 -5506
rect 1991 -5540 2025 -5506
rect 2059 -5540 2093 -5506
rect 2127 -5540 2161 -5506
rect 2195 -5540 2229 -5506
rect 2263 -5540 2297 -5506
rect 2331 -5540 2365 -5506
rect 2399 -5540 2433 -5506
rect 2467 -5540 2501 -5506
rect 2535 -5540 2569 -5506
rect 2603 -5540 2637 -5506
rect 2671 -5540 2705 -5506
rect 2739 -5540 2773 -5506
rect 2807 -5540 2841 -5506
rect 2875 -5540 2909 -5506
rect 2943 -5540 2977 -5506
rect 3011 -5540 3045 -5506
rect 3079 -5540 3113 -5506
rect 3147 -5540 3181 -5506
rect 3215 -5540 3249 -5506
rect 3283 -5540 3317 -5506
rect 3351 -5540 3385 -5506
rect 3419 -5540 3453 -5506
rect 3487 -5540 3521 -5506
rect 3555 -5540 3589 -5506
rect 3623 -5540 3657 -5506
rect 3691 -5540 3725 -5506
rect 3759 -5540 3793 -5506
rect 3827 -5540 3861 -5506
rect 3895 -5540 3929 -5506
rect 3963 -5540 3997 -5506
rect 4031 -5540 4065 -5506
rect 4099 -5540 4133 -5506
rect 4167 -5540 4201 -5506
rect 4235 -5540 4269 -5506
rect 4303 -5540 4337 -5506
rect 4371 -5540 4405 -5506
rect 4439 -5540 4473 -5506
rect 4507 -5540 4541 -5506
rect 4575 -5540 4609 -5506
rect 4643 -5540 4677 -5506
rect 4711 -5540 4745 -5506
rect 4779 -5540 4813 -5506
rect 4847 -5540 4881 -5506
rect 4915 -5540 4949 -5506
rect 4983 -5540 5017 -5506
rect 5051 -5540 5085 -5506
rect 5119 -5540 5153 -5506
rect 5187 -5540 5221 -5506
rect 5255 -5540 5289 -5506
rect 5323 -5540 5357 -5506
rect 5391 -5540 5425 -5506
rect 5459 -5540 5493 -5506
rect 5527 -5540 5561 -5506
rect 5595 -5540 5629 -5506
rect 5663 -5540 5697 -5506
rect 5731 -5540 5765 -5506
rect 5799 -5540 5833 -5506
rect 5867 -5540 5901 -5506
rect 5935 -5540 5969 -5506
rect 6003 -5540 6166 -5506
<< nsubdiffcont >>
rect 461 5922 495 5956
rect 529 5922 563 5956
rect 597 5922 631 5956
rect 665 5922 699 5956
rect 733 5922 767 5956
rect 801 5922 835 5956
rect 869 5922 903 5956
rect 937 5922 971 5956
rect 1005 5922 1039 5956
rect 1073 5922 1107 5956
rect 1141 5922 1175 5956
rect 1209 5922 1243 5956
rect 1277 5922 1311 5956
rect 1345 5922 1379 5956
rect 1413 5922 1447 5956
rect 1481 5922 1515 5956
rect 1549 5922 1583 5956
rect 1617 5922 1651 5956
rect 1685 5922 1719 5956
rect 1753 5922 1787 5956
rect 1821 5922 1855 5956
rect 1889 5922 1923 5956
rect 1957 5922 1991 5956
rect 2025 5922 2059 5956
rect 2093 5922 2127 5956
rect 2161 5922 2195 5956
rect 2229 5922 2263 5956
rect 2297 5922 2331 5956
rect 2365 5922 2399 5956
rect 2433 5922 2467 5956
rect 2501 5922 2535 5956
rect 2569 5922 2603 5956
rect 2637 5922 2671 5956
rect 2705 5922 2739 5956
rect 2773 5922 2807 5956
rect 2841 5922 2875 5956
rect 2909 5922 2943 5956
rect 2977 5922 3011 5956
rect 3045 5922 3079 5956
rect 3113 5922 3147 5956
rect 3181 5922 3215 5956
rect 3249 5922 3283 5956
rect 3317 5922 3351 5956
rect 3385 5922 3419 5956
rect 3453 5922 3487 5956
rect 3521 5922 3555 5956
rect 3589 5922 3623 5956
rect 3657 5922 3691 5956
rect 3725 5922 3759 5956
rect 3793 5922 3827 5956
rect 3861 5922 3895 5956
rect 3929 5922 3963 5956
rect 3997 5922 4031 5956
rect 4065 5922 4099 5956
rect 4133 5922 4167 5956
rect 4201 5922 4235 5956
rect 4269 5922 4303 5956
rect 4337 5922 4371 5956
rect 4405 5922 4439 5956
rect 4473 5922 4507 5956
rect 4541 5922 4575 5956
rect 4609 5922 4643 5956
rect 4677 5922 4711 5956
rect 4745 5922 4779 5956
rect 4813 5922 4847 5956
rect 4881 5922 4915 5956
rect 4949 5922 4983 5956
rect 5017 5922 5051 5956
rect 5085 5922 5119 5956
rect 5153 5922 5187 5956
rect 5221 5922 5255 5956
rect 5289 5922 5323 5956
rect 5357 5922 5391 5956
rect 5425 5922 5459 5956
rect 5493 5922 5527 5956
rect 5561 5922 5595 5956
rect 5629 5922 5663 5956
rect 5697 5922 5731 5956
rect 5765 5922 5799 5956
rect 5833 5922 5867 5956
rect 5901 5922 5935 5956
rect 5969 5922 6003 5956
rect 340 5761 374 5795
rect 340 5693 374 5727
rect 340 5625 374 5659
rect 340 5557 374 5591
rect 6132 5761 6166 5795
rect 6132 5693 6166 5727
rect 6132 5625 6166 5659
rect 340 5489 374 5523
rect 6132 5557 6166 5591
rect 340 5421 374 5455
rect 340 5353 374 5387
rect 340 5285 374 5319
rect 6132 5489 6166 5523
rect 6132 5421 6166 5455
rect 6132 5353 6166 5387
rect 6132 5285 6166 5319
rect 340 5217 374 5251
rect 340 5149 374 5183
rect 6132 5217 6166 5251
rect 340 5081 374 5115
rect 340 5013 374 5047
rect 6132 5149 6166 5183
rect 6132 5081 6166 5115
rect 6132 5013 6166 5047
rect 340 4945 374 4979
rect 340 4877 374 4911
rect 340 4809 374 4843
rect 340 4741 374 4775
rect 340 4673 374 4707
rect 340 4605 374 4639
rect 340 4537 374 4571
rect 340 4469 374 4503
rect 340 4401 374 4435
rect 340 4333 374 4367
rect 6132 4945 6166 4979
rect 6132 4877 6166 4911
rect 6132 4809 6166 4843
rect 6132 4741 6166 4775
rect 6132 4673 6166 4707
rect 6132 4605 6166 4639
rect 6132 4537 6166 4571
rect 6132 4469 6166 4503
rect 6132 4401 6166 4435
rect 6132 4333 6166 4367
rect 340 4265 374 4299
rect 340 4197 374 4231
rect 340 4129 374 4163
rect 340 4061 374 4095
rect 6132 4265 6166 4299
rect 6132 4197 6166 4231
rect 6132 4129 6166 4163
rect 340 3993 374 4027
rect 6132 4061 6166 4095
rect 6132 3993 6166 4027
rect 340 3925 374 3959
rect 340 3857 374 3891
rect 340 3789 374 3823
rect 6132 3925 6166 3959
rect 6132 3857 6166 3891
rect 6132 3789 6166 3823
rect 340 3721 374 3755
rect 340 3653 374 3687
rect 6132 3721 6166 3755
rect 340 3585 374 3619
rect 340 3517 374 3551
rect 340 3449 374 3483
rect 6132 3653 6166 3687
rect 6132 3585 6166 3619
rect 6132 3517 6166 3551
rect 340 3381 374 3415
rect 340 3313 374 3347
rect 340 3245 374 3279
rect 340 3177 374 3211
rect 340 3109 374 3143
rect 340 3041 374 3075
rect 340 2973 374 3007
rect 340 2905 374 2939
rect 340 2837 374 2871
rect 6132 3449 6166 3483
rect 6132 3381 6166 3415
rect 6132 3313 6166 3347
rect 6132 3245 6166 3279
rect 6132 3177 6166 3211
rect 6132 3109 6166 3143
rect 6132 3041 6166 3075
rect 6132 2973 6166 3007
rect 6132 2905 6166 2939
rect 6132 2837 6166 2871
rect 340 2769 374 2803
rect 340 2701 374 2735
rect 340 2633 374 2667
rect 340 2565 374 2599
rect 6132 2769 6166 2803
rect 6132 2701 6166 2735
rect 6132 2633 6166 2667
rect 340 2497 374 2531
rect 6132 2565 6166 2599
rect 6132 2497 6166 2531
rect 340 2429 374 2463
rect 340 2361 374 2395
rect 340 2293 374 2327
rect 6132 2429 6166 2463
rect 6132 2361 6166 2395
rect 6132 2293 6166 2327
rect 340 2225 374 2259
rect 340 2157 374 2191
rect 6132 2225 6166 2259
rect 340 2089 374 2123
rect 6132 2157 6166 2191
rect 6132 2089 6166 2123
rect 340 1848 374 1882
rect 340 1780 374 1814
rect 340 1712 374 1746
rect 340 1644 374 1678
rect 340 1576 374 1610
rect 6132 1848 6166 1882
rect 6132 1780 6166 1814
rect 6132 1712 6166 1746
rect 6132 1644 6166 1678
rect 6132 1576 6166 1610
rect 340 1508 374 1542
rect 340 1440 374 1474
rect 6132 1508 6166 1542
rect 6132 1440 6166 1474
rect 340 1372 374 1406
rect 340 1304 374 1338
rect 340 1236 374 1270
rect 6132 1372 6166 1406
rect 6132 1304 6166 1338
rect 6132 1236 6166 1270
rect 340 1168 374 1202
rect 340 1100 374 1134
rect 6132 1168 6166 1202
rect 340 1032 374 1066
rect 340 964 374 998
rect 340 896 374 930
rect 6132 1100 6166 1134
rect 6132 1032 6166 1066
rect 6132 964 6166 998
rect 340 828 374 862
rect 6132 896 6166 930
rect 6132 828 6166 862
rect 340 760 374 794
rect 340 692 374 726
rect 340 624 374 658
rect 6132 760 6166 794
rect 6132 692 6166 726
rect 6132 624 6166 658
rect 340 556 374 590
rect 340 488 374 522
rect 340 420 374 454
rect 340 352 374 386
rect 6132 556 6166 590
rect 6132 488 6166 522
rect 6132 420 6166 454
rect 6132 352 6166 386
rect 340 284 374 318
rect 340 216 374 250
rect 340 148 374 182
rect 6132 284 6166 318
rect 6132 216 6166 250
rect 6132 148 6166 182
rect 340 80 374 114
rect 340 12 374 46
rect 6132 80 6166 114
rect 340 -56 374 -22
rect 340 -124 374 -90
rect 340 -192 374 -158
rect 6132 12 6166 46
rect 6132 -56 6166 -22
rect 6132 -124 6166 -90
rect 6132 -192 6166 -158
rect 340 -260 374 -226
rect 340 -328 374 -294
rect 6132 -260 6166 -226
rect 340 -396 374 -362
rect 340 -464 374 -430
rect 6132 -328 6166 -294
rect 6132 -396 6166 -362
rect 6132 -464 6166 -430
rect 340 -532 374 -498
rect 340 -600 374 -566
rect 340 -668 374 -634
rect 340 -736 374 -702
rect 6132 -532 6166 -498
rect 6132 -600 6166 -566
rect 6132 -668 6166 -634
rect 6132 -736 6166 -702
rect 340 -804 374 -770
rect 340 -872 374 -838
rect 340 -940 374 -906
rect 6132 -804 6166 -770
rect 6132 -872 6166 -838
rect 6132 -940 6166 -906
rect 340 -1008 374 -974
rect 340 -1076 374 -1042
rect 6132 -1008 6166 -974
rect 340 -1144 374 -1110
rect 6132 -1076 6166 -1042
rect 6132 -1144 6166 -1110
rect 340 -1212 374 -1178
rect 340 -1280 374 -1246
rect 6132 -1212 6166 -1178
rect 6132 -1280 6166 -1246
rect 340 -1348 374 -1314
rect 6132 -1348 6166 -1314
rect 340 -1416 374 -1382
rect 340 -1484 374 -1450
rect 340 -1552 374 -1518
rect 6132 -1416 6166 -1382
rect 6132 -1484 6166 -1450
rect 6132 -1552 6166 -1518
rect 340 -1620 374 -1586
rect 340 -1688 374 -1654
rect 340 -1756 374 -1722
rect 340 -1824 374 -1790
rect 340 -1892 374 -1858
rect 340 -1960 374 -1926
rect 340 -2028 374 -1994
rect 340 -2096 374 -2062
rect 340 -2164 374 -2130
rect 340 -2232 374 -2198
rect 6132 -1620 6166 -1586
rect 6132 -1688 6166 -1654
rect 6132 -1756 6166 -1722
rect 6132 -1824 6166 -1790
rect 6132 -1892 6166 -1858
rect 6132 -1960 6166 -1926
rect 6132 -2028 6166 -1994
rect 6132 -2096 6166 -2062
rect 6132 -2164 6166 -2130
rect 6132 -2232 6166 -2198
rect 340 -2300 374 -2266
rect 340 -2368 374 -2334
rect 340 -2436 374 -2402
rect 340 -2504 374 -2470
rect 6132 -2300 6166 -2266
rect 6132 -2368 6166 -2334
rect 6132 -2436 6166 -2402
rect 340 -2572 374 -2538
rect 6132 -2504 6166 -2470
rect 6132 -2572 6166 -2538
rect 340 -2640 374 -2606
rect 340 -2708 374 -2674
rect 340 -2776 374 -2742
rect 6132 -2640 6166 -2606
rect 6132 -2708 6166 -2674
rect 6132 -2776 6166 -2742
rect 340 -2844 374 -2810
rect 340 -2912 374 -2878
rect 6132 -2844 6166 -2810
rect 340 -2980 374 -2946
rect 340 -3048 374 -3014
rect 340 -3116 374 -3082
rect 6132 -2912 6166 -2878
rect 6132 -2980 6166 -2946
rect 6132 -3048 6166 -3014
rect 340 -3184 374 -3150
rect 340 -3252 374 -3218
rect 340 -3320 374 -3286
rect 340 -3388 374 -3354
rect 340 -3456 374 -3422
rect 340 -3524 374 -3490
rect 340 -3592 374 -3558
rect 340 -3660 374 -3626
rect 340 -3728 374 -3694
rect 6132 -3116 6166 -3082
rect 6132 -3184 6166 -3150
rect 6132 -3252 6166 -3218
rect 6132 -3320 6166 -3286
rect 6132 -3388 6166 -3354
rect 6132 -3456 6166 -3422
rect 6132 -3524 6166 -3490
rect 6132 -3592 6166 -3558
rect 6132 -3660 6166 -3626
rect 6132 -3728 6166 -3694
rect 340 -3796 374 -3762
rect 340 -3864 374 -3830
rect 340 -3932 374 -3898
rect 340 -4000 374 -3966
rect 6132 -3796 6166 -3762
rect 6132 -3864 6166 -3830
rect 6132 -3932 6166 -3898
rect 340 -4068 374 -4034
rect 6132 -4000 6166 -3966
rect 6132 -4068 6166 -4034
rect 340 -4136 374 -4102
rect 340 -4204 374 -4170
rect 340 -4272 374 -4238
rect 6132 -4136 6166 -4102
rect 6132 -4204 6166 -4170
rect 6132 -4272 6166 -4238
rect 340 -4340 374 -4306
rect 340 -4408 374 -4374
rect 6132 -4340 6166 -4306
rect 340 -4476 374 -4442
rect 340 -4544 374 -4510
rect 340 -4612 374 -4578
rect 6132 -4408 6166 -4374
rect 6132 -4476 6166 -4442
rect 6132 -4544 6166 -4510
rect 6132 -4612 6166 -4578
rect 340 -4680 374 -4646
rect 340 -4748 374 -4714
rect 340 -4816 374 -4782
rect 340 -4884 374 -4850
rect 340 -4952 374 -4918
rect 340 -5020 374 -4986
rect 340 -5088 374 -5054
rect 6132 -4680 6166 -4646
rect 6132 -4748 6166 -4714
rect 6132 -4816 6166 -4782
rect 6132 -4884 6166 -4850
rect 6132 -4952 6166 -4918
rect 6132 -5020 6166 -4986
rect 6132 -5088 6166 -5054
rect 340 -5156 374 -5122
rect 340 -5224 374 -5190
rect 340 -5292 374 -5258
rect 340 -5360 374 -5326
rect 6132 -5156 6166 -5122
rect 6132 -5224 6166 -5190
rect 6132 -5292 6166 -5258
rect 6132 -5360 6166 -5326
rect 461 -5540 495 -5506
rect 529 -5540 563 -5506
rect 597 -5540 631 -5506
rect 665 -5540 699 -5506
rect 733 -5540 767 -5506
rect 801 -5540 835 -5506
rect 869 -5540 903 -5506
rect 937 -5540 971 -5506
rect 1005 -5540 1039 -5506
rect 1073 -5540 1107 -5506
rect 1141 -5540 1175 -5506
rect 1209 -5540 1243 -5506
rect 1277 -5540 1311 -5506
rect 1345 -5540 1379 -5506
rect 1413 -5540 1447 -5506
rect 1481 -5540 1515 -5506
rect 1549 -5540 1583 -5506
rect 1617 -5540 1651 -5506
rect 1685 -5540 1719 -5506
rect 1753 -5540 1787 -5506
rect 1821 -5540 1855 -5506
rect 1889 -5540 1923 -5506
rect 1957 -5540 1991 -5506
rect 2025 -5540 2059 -5506
rect 2093 -5540 2127 -5506
rect 2161 -5540 2195 -5506
rect 2229 -5540 2263 -5506
rect 2297 -5540 2331 -5506
rect 2365 -5540 2399 -5506
rect 2433 -5540 2467 -5506
rect 2501 -5540 2535 -5506
rect 2569 -5540 2603 -5506
rect 2637 -5540 2671 -5506
rect 2705 -5540 2739 -5506
rect 2773 -5540 2807 -5506
rect 2841 -5540 2875 -5506
rect 2909 -5540 2943 -5506
rect 2977 -5540 3011 -5506
rect 3045 -5540 3079 -5506
rect 3113 -5540 3147 -5506
rect 3181 -5540 3215 -5506
rect 3249 -5540 3283 -5506
rect 3317 -5540 3351 -5506
rect 3385 -5540 3419 -5506
rect 3453 -5540 3487 -5506
rect 3521 -5540 3555 -5506
rect 3589 -5540 3623 -5506
rect 3657 -5540 3691 -5506
rect 3725 -5540 3759 -5506
rect 3793 -5540 3827 -5506
rect 3861 -5540 3895 -5506
rect 3929 -5540 3963 -5506
rect 3997 -5540 4031 -5506
rect 4065 -5540 4099 -5506
rect 4133 -5540 4167 -5506
rect 4201 -5540 4235 -5506
rect 4269 -5540 4303 -5506
rect 4337 -5540 4371 -5506
rect 4405 -5540 4439 -5506
rect 4473 -5540 4507 -5506
rect 4541 -5540 4575 -5506
rect 4609 -5540 4643 -5506
rect 4677 -5540 4711 -5506
rect 4745 -5540 4779 -5506
rect 4813 -5540 4847 -5506
rect 4881 -5540 4915 -5506
rect 4949 -5540 4983 -5506
rect 5017 -5540 5051 -5506
rect 5085 -5540 5119 -5506
rect 5153 -5540 5187 -5506
rect 5221 -5540 5255 -5506
rect 5289 -5540 5323 -5506
rect 5357 -5540 5391 -5506
rect 5425 -5540 5459 -5506
rect 5493 -5540 5527 -5506
rect 5561 -5540 5595 -5506
rect 5629 -5540 5663 -5506
rect 5697 -5540 5731 -5506
rect 5765 -5540 5799 -5506
rect 5833 -5540 5867 -5506
rect 5901 -5540 5935 -5506
rect 5969 -5540 6003 -5506
<< poly >>
rect 576 5789 776 5815
rect 834 5789 1034 5815
rect 1286 5789 1486 5815
rect 1544 5789 1744 5815
rect 1802 5789 2002 5815
rect 2060 5789 2260 5815
rect 2512 5789 2712 5815
rect 2770 5789 2970 5815
rect 3028 5789 3228 5815
rect 3286 5789 3486 5815
rect 3544 5789 3744 5815
rect 3802 5789 4002 5815
rect 4254 5789 4454 5815
rect 4512 5789 4712 5815
rect 4770 5789 4970 5815
rect 5028 5789 5228 5815
rect 5479 5789 5679 5815
rect 5737 5789 5937 5815
rect 576 5542 776 5589
rect 576 5508 625 5542
rect 659 5508 693 5542
rect 727 5508 776 5542
rect 576 5492 776 5508
rect 834 5542 1034 5589
rect 834 5508 883 5542
rect 917 5508 951 5542
rect 985 5508 1034 5542
rect 834 5492 1034 5508
rect 1286 5542 1486 5589
rect 1286 5508 1335 5542
rect 1369 5508 1403 5542
rect 1437 5508 1486 5542
rect 1286 5492 1486 5508
rect 1544 5542 1744 5589
rect 1544 5508 1593 5542
rect 1627 5508 1661 5542
rect 1695 5508 1744 5542
rect 1544 5492 1744 5508
rect 1802 5542 2002 5589
rect 1802 5508 1851 5542
rect 1885 5508 1919 5542
rect 1953 5508 2002 5542
rect 1802 5492 2002 5508
rect 2060 5542 2260 5589
rect 2060 5508 2109 5542
rect 2143 5508 2177 5542
rect 2211 5508 2260 5542
rect 2060 5492 2260 5508
rect 2512 5542 2712 5589
rect 2512 5508 2561 5542
rect 2595 5508 2629 5542
rect 2663 5508 2712 5542
rect 2512 5492 2712 5508
rect 2770 5542 2970 5589
rect 2770 5508 2819 5542
rect 2853 5508 2887 5542
rect 2921 5508 2970 5542
rect 2770 5492 2970 5508
rect 3028 5542 3228 5589
rect 3028 5508 3077 5542
rect 3111 5508 3145 5542
rect 3179 5508 3228 5542
rect 3028 5492 3228 5508
rect 3286 5542 3486 5589
rect 3286 5508 3335 5542
rect 3369 5508 3403 5542
rect 3437 5508 3486 5542
rect 3286 5492 3486 5508
rect 3544 5542 3744 5589
rect 3544 5508 3593 5542
rect 3627 5508 3661 5542
rect 3695 5508 3744 5542
rect 3544 5492 3744 5508
rect 3802 5542 4002 5589
rect 3802 5508 3851 5542
rect 3885 5508 3919 5542
rect 3953 5508 4002 5542
rect 3802 5492 4002 5508
rect 4254 5542 4454 5589
rect 4254 5508 4303 5542
rect 4337 5508 4371 5542
rect 4405 5508 4454 5542
rect 4254 5492 4454 5508
rect 4512 5542 4712 5589
rect 4512 5508 4561 5542
rect 4595 5508 4629 5542
rect 4663 5508 4712 5542
rect 4512 5492 4712 5508
rect 4770 5542 4970 5589
rect 4770 5508 4819 5542
rect 4853 5508 4887 5542
rect 4921 5508 4970 5542
rect 4770 5492 4970 5508
rect 5028 5542 5228 5589
rect 5028 5508 5077 5542
rect 5111 5508 5145 5542
rect 5179 5508 5228 5542
rect 5028 5492 5228 5508
rect 5479 5542 5679 5589
rect 5479 5508 5528 5542
rect 5562 5508 5596 5542
rect 5630 5508 5679 5542
rect 5479 5492 5679 5508
rect 5737 5542 5937 5589
rect 5737 5508 5786 5542
rect 5820 5508 5854 5542
rect 5888 5508 5937 5542
rect 5737 5492 5937 5508
rect 576 5261 776 5277
rect 576 5227 625 5261
rect 659 5227 693 5261
rect 727 5227 776 5261
rect 576 5180 776 5227
rect 834 5261 1034 5277
rect 834 5227 883 5261
rect 917 5227 951 5261
rect 985 5227 1034 5261
rect 834 5180 1034 5227
rect 5479 5261 5679 5277
rect 5479 5227 5528 5261
rect 5562 5227 5596 5261
rect 5630 5227 5679 5261
rect 5479 5180 5679 5227
rect 5737 5261 5937 5277
rect 5737 5227 5786 5261
rect 5820 5227 5854 5261
rect 5888 5227 5937 5261
rect 5737 5180 5937 5227
rect 576 4954 776 4980
rect 834 4954 1034 4980
rect 5479 4954 5679 4980
rect 5737 4954 5937 4980
rect 576 4285 776 4311
rect 834 4285 1034 4311
rect 5479 4285 5679 4311
rect 5737 4285 5937 4311
rect 576 4038 776 4085
rect 576 4004 625 4038
rect 659 4004 693 4038
rect 727 4004 776 4038
rect 576 3988 776 4004
rect 834 4038 1034 4085
rect 834 4004 883 4038
rect 917 4004 951 4038
rect 985 4004 1034 4038
rect 834 3988 1034 4004
rect 5479 4038 5679 4085
rect 5479 4004 5528 4038
rect 5562 4004 5596 4038
rect 5630 4004 5679 4038
rect 5479 3988 5679 4004
rect 5737 4038 5937 4085
rect 5737 4004 5786 4038
rect 5820 4004 5854 4038
rect 5888 4004 5937 4038
rect 5737 3988 5937 4004
rect 576 3757 776 3773
rect 576 3723 625 3757
rect 659 3723 693 3757
rect 727 3723 776 3757
rect 576 3676 776 3723
rect 834 3757 1034 3773
rect 834 3723 883 3757
rect 917 3723 951 3757
rect 985 3723 1034 3757
rect 834 3676 1034 3723
rect 5479 3757 5679 3773
rect 5479 3723 5528 3757
rect 5562 3723 5596 3757
rect 5630 3723 5679 3757
rect 5479 3676 5679 3723
rect 5737 3757 5937 3773
rect 5737 3723 5786 3757
rect 5820 3723 5854 3757
rect 5888 3723 5937 3757
rect 5737 3676 5937 3723
rect 576 3450 776 3476
rect 834 3450 1034 3476
rect 5479 3450 5679 3476
rect 5737 3450 5937 3476
rect 576 2778 776 2804
rect 834 2778 1034 2804
rect 5479 2778 5679 2804
rect 5737 2778 5937 2804
rect 576 2531 776 2578
rect 576 2497 625 2531
rect 659 2497 693 2531
rect 727 2497 776 2531
rect 576 2481 776 2497
rect 834 2531 1034 2578
rect 834 2497 883 2531
rect 917 2497 951 2531
rect 985 2497 1034 2531
rect 834 2481 1034 2497
rect 5479 2531 5679 2578
rect 5479 2497 5528 2531
rect 5562 2497 5596 2531
rect 5630 2497 5679 2531
rect 5479 2481 5679 2497
rect 5737 2531 5937 2578
rect 5737 2497 5786 2531
rect 5820 2497 5854 2531
rect 5888 2497 5937 2531
rect 5737 2481 5937 2497
rect 576 2250 776 2266
rect 576 2216 625 2250
rect 659 2216 693 2250
rect 727 2216 776 2250
rect 576 2169 776 2216
rect 834 2250 1034 2266
rect 834 2216 883 2250
rect 917 2216 951 2250
rect 985 2216 1034 2250
rect 834 2169 1034 2216
rect 5479 2250 5679 2266
rect 5479 2216 5528 2250
rect 5562 2216 5596 2250
rect 5630 2216 5679 2250
rect 5479 2169 5679 2216
rect 5737 2250 5937 2266
rect 5737 2216 5786 2250
rect 5820 2216 5854 2250
rect 5888 2216 5937 2250
rect 5737 2169 5937 2216
rect 576 1943 776 1969
rect 834 1943 1034 1969
rect 5479 1943 5679 1969
rect 5737 1943 5937 1969
rect 576 1409 776 1435
rect 834 1409 1034 1435
rect 5479 1409 5679 1435
rect 5737 1409 5937 1435
rect 576 1162 776 1209
rect 576 1128 625 1162
rect 659 1128 693 1162
rect 727 1128 776 1162
rect 576 1112 776 1128
rect 834 1162 1034 1209
rect 834 1128 883 1162
rect 917 1128 951 1162
rect 985 1128 1034 1162
rect 834 1112 1034 1128
rect 5479 1162 5679 1209
rect 5479 1128 5528 1162
rect 5562 1128 5596 1162
rect 5630 1128 5679 1162
rect 5479 1112 5679 1128
rect 5737 1162 5937 1209
rect 5737 1128 5786 1162
rect 5820 1128 5854 1162
rect 5888 1128 5937 1162
rect 5737 1112 5937 1128
rect 576 881 776 897
rect 576 847 625 881
rect 659 847 693 881
rect 727 847 776 881
rect 576 800 776 847
rect 834 881 1034 897
rect 834 847 883 881
rect 917 847 951 881
rect 985 847 1034 881
rect 834 800 1034 847
rect 5479 881 5679 897
rect 5479 847 5528 881
rect 5562 847 5596 881
rect 5630 847 5679 881
rect 5479 800 5679 847
rect 5737 881 5937 897
rect 5737 847 5786 881
rect 5820 847 5854 881
rect 5888 847 5937 881
rect 5737 800 5937 847
rect 576 574 776 600
rect 834 574 1034 600
rect 5479 574 5679 600
rect 5737 574 5937 600
rect 576 314 776 340
rect 834 314 1034 340
rect 5479 314 5679 340
rect 5737 314 5937 340
rect 576 67 776 114
rect 576 33 625 67
rect 659 33 693 67
rect 727 33 776 67
rect 576 17 776 33
rect 834 67 1034 114
rect 834 33 883 67
rect 917 33 951 67
rect 985 33 1034 67
rect 834 17 1034 33
rect 5479 67 5679 114
rect 5479 33 5528 67
rect 5562 33 5596 67
rect 5630 33 5679 67
rect 5479 17 5679 33
rect 5737 67 5937 114
rect 5737 33 5786 67
rect 5820 33 5854 67
rect 5888 33 5937 67
rect 5737 17 5937 33
rect 576 -214 776 -198
rect 576 -248 625 -214
rect 659 -248 693 -214
rect 727 -248 776 -214
rect 576 -295 776 -248
rect 834 -214 1034 -198
rect 834 -248 883 -214
rect 917 -248 951 -214
rect 985 -248 1034 -214
rect 834 -295 1034 -248
rect 5479 -214 5679 -198
rect 5479 -248 5528 -214
rect 5562 -248 5596 -214
rect 5630 -248 5679 -214
rect 5479 -295 5679 -248
rect 5737 -214 5937 -198
rect 5737 -248 5786 -214
rect 5820 -248 5854 -214
rect 5888 -248 5937 -214
rect 5737 -295 5937 -248
rect 576 -521 776 -495
rect 834 -521 1034 -495
rect 5479 -521 5679 -495
rect 5737 -521 5937 -495
rect 576 -772 776 -746
rect 834 -772 1034 -746
rect 5479 -772 5679 -746
rect 5737 -772 5937 -746
rect 576 -1019 776 -972
rect 576 -1053 625 -1019
rect 659 -1053 693 -1019
rect 727 -1053 776 -1019
rect 576 -1069 776 -1053
rect 834 -1019 1034 -972
rect 834 -1053 883 -1019
rect 917 -1053 951 -1019
rect 985 -1053 1034 -1019
rect 834 -1069 1034 -1053
rect 5479 -1019 5679 -972
rect 5479 -1053 5528 -1019
rect 5562 -1053 5596 -1019
rect 5630 -1053 5679 -1019
rect 5479 -1069 5679 -1053
rect 5737 -1019 5937 -972
rect 5737 -1053 5786 -1019
rect 5820 -1053 5854 -1019
rect 5888 -1053 5937 -1019
rect 5737 -1069 5937 -1053
rect 576 -1300 776 -1284
rect 576 -1334 625 -1300
rect 659 -1334 693 -1300
rect 727 -1334 776 -1300
rect 576 -1381 776 -1334
rect 834 -1300 1034 -1284
rect 834 -1334 883 -1300
rect 917 -1334 951 -1300
rect 985 -1334 1034 -1300
rect 834 -1381 1034 -1334
rect 5479 -1300 5679 -1284
rect 5479 -1334 5528 -1300
rect 5562 -1334 5596 -1300
rect 5630 -1334 5679 -1300
rect 5479 -1381 5679 -1334
rect 5737 -1300 5937 -1284
rect 5737 -1334 5786 -1300
rect 5820 -1334 5854 -1300
rect 5888 -1334 5937 -1300
rect 5737 -1381 5937 -1334
rect 576 -1607 776 -1581
rect 834 -1607 1034 -1581
rect 5479 -1607 5679 -1581
rect 5737 -1607 5937 -1581
rect 576 -2276 776 -2250
rect 834 -2276 1034 -2250
rect 5479 -2276 5679 -2250
rect 5737 -2276 5937 -2250
rect 576 -2523 776 -2476
rect 576 -2557 625 -2523
rect 659 -2557 693 -2523
rect 727 -2557 776 -2523
rect 576 -2573 776 -2557
rect 834 -2523 1034 -2476
rect 834 -2557 883 -2523
rect 917 -2557 951 -2523
rect 985 -2557 1034 -2523
rect 834 -2573 1034 -2557
rect 5479 -2523 5679 -2476
rect 5479 -2557 5528 -2523
rect 5562 -2557 5596 -2523
rect 5630 -2557 5679 -2523
rect 5479 -2573 5679 -2557
rect 5737 -2523 5937 -2476
rect 5737 -2557 5786 -2523
rect 5820 -2557 5854 -2523
rect 5888 -2557 5937 -2523
rect 5737 -2573 5937 -2557
rect 576 -2804 776 -2788
rect 576 -2838 625 -2804
rect 659 -2838 693 -2804
rect 727 -2838 776 -2804
rect 576 -2885 776 -2838
rect 834 -2804 1034 -2788
rect 834 -2838 883 -2804
rect 917 -2838 951 -2804
rect 985 -2838 1034 -2804
rect 834 -2885 1034 -2838
rect 5479 -2804 5679 -2788
rect 5479 -2838 5528 -2804
rect 5562 -2838 5596 -2804
rect 5630 -2838 5679 -2804
rect 5479 -2885 5679 -2838
rect 5737 -2804 5937 -2788
rect 5737 -2838 5786 -2804
rect 5820 -2838 5854 -2804
rect 5888 -2838 5937 -2804
rect 5737 -2885 5937 -2838
rect 576 -3111 776 -3085
rect 834 -3111 1034 -3085
rect 5479 -3111 5679 -3085
rect 5737 -3111 5937 -3085
rect 576 -3780 776 -3754
rect 834 -3780 1034 -3754
rect 5479 -3780 5679 -3754
rect 5737 -3780 5937 -3754
rect 576 -4027 776 -3980
rect 576 -4061 625 -4027
rect 659 -4061 693 -4027
rect 727 -4061 776 -4027
rect 576 -4077 776 -4061
rect 834 -4027 1034 -3980
rect 834 -4061 883 -4027
rect 917 -4061 951 -4027
rect 985 -4061 1034 -4027
rect 834 -4077 1034 -4061
rect 5479 -4027 5679 -3980
rect 5479 -4061 5528 -4027
rect 5562 -4061 5596 -4027
rect 5630 -4061 5679 -4027
rect 5479 -4077 5679 -4061
rect 5737 -4027 5937 -3980
rect 5737 -4061 5786 -4027
rect 5820 -4061 5854 -4027
rect 5888 -4061 5937 -4027
rect 5737 -4077 5937 -4061
rect 576 -4308 776 -4292
rect 576 -4342 625 -4308
rect 659 -4342 693 -4308
rect 727 -4342 776 -4308
rect 576 -4389 776 -4342
rect 834 -4308 1034 -4292
rect 834 -4342 883 -4308
rect 917 -4342 951 -4308
rect 985 -4342 1034 -4308
rect 834 -4389 1034 -4342
rect 5479 -4308 5679 -4292
rect 5479 -4342 5528 -4308
rect 5562 -4342 5596 -4308
rect 5630 -4342 5679 -4308
rect 5479 -4389 5679 -4342
rect 5737 -4308 5937 -4292
rect 5737 -4342 5786 -4308
rect 5820 -4342 5854 -4308
rect 5888 -4342 5937 -4308
rect 5737 -4389 5937 -4342
rect 576 -4615 776 -4589
rect 834 -4615 1034 -4589
rect 5479 -4615 5679 -4589
rect 5737 -4615 5937 -4589
rect 576 -5136 776 -5110
rect 834 -5136 1034 -5110
rect 1286 -5136 1486 -5110
rect 1544 -5136 1744 -5110
rect 1802 -5136 2002 -5110
rect 2060 -5136 2260 -5110
rect 2512 -5136 2712 -5110
rect 2770 -5136 2970 -5110
rect 3028 -5136 3228 -5110
rect 3286 -5136 3486 -5110
rect 3544 -5136 3744 -5110
rect 3802 -5136 4002 -5110
rect 4254 -5136 4454 -5110
rect 4512 -5136 4712 -5110
rect 4770 -5136 4970 -5110
rect 5028 -5136 5228 -5110
rect 5479 -5136 5679 -5110
rect 5737 -5136 5937 -5110
rect 576 -5383 776 -5336
rect 576 -5417 625 -5383
rect 659 -5417 693 -5383
rect 727 -5417 776 -5383
rect 576 -5433 776 -5417
rect 834 -5383 1034 -5336
rect 834 -5417 883 -5383
rect 917 -5417 951 -5383
rect 985 -5417 1034 -5383
rect 834 -5433 1034 -5417
rect 1286 -5383 1486 -5336
rect 1286 -5417 1335 -5383
rect 1369 -5417 1403 -5383
rect 1437 -5417 1486 -5383
rect 1286 -5433 1486 -5417
rect 1544 -5383 1744 -5336
rect 1544 -5417 1593 -5383
rect 1627 -5417 1661 -5383
rect 1695 -5417 1744 -5383
rect 1544 -5433 1744 -5417
rect 1802 -5383 2002 -5336
rect 1802 -5417 1851 -5383
rect 1885 -5417 1919 -5383
rect 1953 -5417 2002 -5383
rect 1802 -5433 2002 -5417
rect 2060 -5383 2260 -5336
rect 2060 -5417 2109 -5383
rect 2143 -5417 2177 -5383
rect 2211 -5417 2260 -5383
rect 2060 -5433 2260 -5417
rect 2512 -5383 2712 -5336
rect 2512 -5417 2561 -5383
rect 2595 -5417 2629 -5383
rect 2663 -5417 2712 -5383
rect 2512 -5433 2712 -5417
rect 2770 -5383 2970 -5336
rect 2770 -5417 2819 -5383
rect 2853 -5417 2887 -5383
rect 2921 -5417 2970 -5383
rect 2770 -5433 2970 -5417
rect 3028 -5383 3228 -5336
rect 3028 -5417 3077 -5383
rect 3111 -5417 3145 -5383
rect 3179 -5417 3228 -5383
rect 3028 -5433 3228 -5417
rect 3286 -5383 3486 -5336
rect 3286 -5417 3335 -5383
rect 3369 -5417 3403 -5383
rect 3437 -5417 3486 -5383
rect 3286 -5433 3486 -5417
rect 3544 -5383 3744 -5336
rect 3544 -5417 3593 -5383
rect 3627 -5417 3661 -5383
rect 3695 -5417 3744 -5383
rect 3544 -5433 3744 -5417
rect 3802 -5383 4002 -5336
rect 3802 -5417 3851 -5383
rect 3885 -5417 3919 -5383
rect 3953 -5417 4002 -5383
rect 3802 -5433 4002 -5417
rect 4254 -5383 4454 -5336
rect 4254 -5417 4303 -5383
rect 4337 -5417 4371 -5383
rect 4405 -5417 4454 -5383
rect 4254 -5433 4454 -5417
rect 4512 -5383 4712 -5336
rect 4512 -5417 4561 -5383
rect 4595 -5417 4629 -5383
rect 4663 -5417 4712 -5383
rect 4512 -5433 4712 -5417
rect 4770 -5383 4970 -5336
rect 4770 -5417 4819 -5383
rect 4853 -5417 4887 -5383
rect 4921 -5417 4970 -5383
rect 4770 -5433 4970 -5417
rect 5028 -5383 5228 -5336
rect 5028 -5417 5077 -5383
rect 5111 -5417 5145 -5383
rect 5179 -5417 5228 -5383
rect 5028 -5433 5228 -5417
rect 5479 -5383 5679 -5336
rect 5479 -5417 5528 -5383
rect 5562 -5417 5596 -5383
rect 5630 -5417 5679 -5383
rect 5479 -5433 5679 -5417
rect 5737 -5383 5937 -5336
rect 5737 -5417 5786 -5383
rect 5820 -5417 5854 -5383
rect 5888 -5417 5937 -5383
rect 5737 -5433 5937 -5417
<< polycont >>
rect 625 5508 659 5542
rect 693 5508 727 5542
rect 883 5508 917 5542
rect 951 5508 985 5542
rect 1335 5508 1369 5542
rect 1403 5508 1437 5542
rect 1593 5508 1627 5542
rect 1661 5508 1695 5542
rect 1851 5508 1885 5542
rect 1919 5508 1953 5542
rect 2109 5508 2143 5542
rect 2177 5508 2211 5542
rect 2561 5508 2595 5542
rect 2629 5508 2663 5542
rect 2819 5508 2853 5542
rect 2887 5508 2921 5542
rect 3077 5508 3111 5542
rect 3145 5508 3179 5542
rect 3335 5508 3369 5542
rect 3403 5508 3437 5542
rect 3593 5508 3627 5542
rect 3661 5508 3695 5542
rect 3851 5508 3885 5542
rect 3919 5508 3953 5542
rect 4303 5508 4337 5542
rect 4371 5508 4405 5542
rect 4561 5508 4595 5542
rect 4629 5508 4663 5542
rect 4819 5508 4853 5542
rect 4887 5508 4921 5542
rect 5077 5508 5111 5542
rect 5145 5508 5179 5542
rect 5528 5508 5562 5542
rect 5596 5508 5630 5542
rect 5786 5508 5820 5542
rect 5854 5508 5888 5542
rect 625 5227 659 5261
rect 693 5227 727 5261
rect 883 5227 917 5261
rect 951 5227 985 5261
rect 5528 5227 5562 5261
rect 5596 5227 5630 5261
rect 5786 5227 5820 5261
rect 5854 5227 5888 5261
rect 625 4004 659 4038
rect 693 4004 727 4038
rect 883 4004 917 4038
rect 951 4004 985 4038
rect 5528 4004 5562 4038
rect 5596 4004 5630 4038
rect 5786 4004 5820 4038
rect 5854 4004 5888 4038
rect 625 3723 659 3757
rect 693 3723 727 3757
rect 883 3723 917 3757
rect 951 3723 985 3757
rect 5528 3723 5562 3757
rect 5596 3723 5630 3757
rect 5786 3723 5820 3757
rect 5854 3723 5888 3757
rect 625 2497 659 2531
rect 693 2497 727 2531
rect 883 2497 917 2531
rect 951 2497 985 2531
rect 5528 2497 5562 2531
rect 5596 2497 5630 2531
rect 5786 2497 5820 2531
rect 5854 2497 5888 2531
rect 625 2216 659 2250
rect 693 2216 727 2250
rect 883 2216 917 2250
rect 951 2216 985 2250
rect 5528 2216 5562 2250
rect 5596 2216 5630 2250
rect 5786 2216 5820 2250
rect 5854 2216 5888 2250
rect 625 1128 659 1162
rect 693 1128 727 1162
rect 883 1128 917 1162
rect 951 1128 985 1162
rect 5528 1128 5562 1162
rect 5596 1128 5630 1162
rect 5786 1128 5820 1162
rect 5854 1128 5888 1162
rect 625 847 659 881
rect 693 847 727 881
rect 883 847 917 881
rect 951 847 985 881
rect 5528 847 5562 881
rect 5596 847 5630 881
rect 5786 847 5820 881
rect 5854 847 5888 881
rect 625 33 659 67
rect 693 33 727 67
rect 883 33 917 67
rect 951 33 985 67
rect 5528 33 5562 67
rect 5596 33 5630 67
rect 5786 33 5820 67
rect 5854 33 5888 67
rect 625 -248 659 -214
rect 693 -248 727 -214
rect 883 -248 917 -214
rect 951 -248 985 -214
rect 5528 -248 5562 -214
rect 5596 -248 5630 -214
rect 5786 -248 5820 -214
rect 5854 -248 5888 -214
rect 625 -1053 659 -1019
rect 693 -1053 727 -1019
rect 883 -1053 917 -1019
rect 951 -1053 985 -1019
rect 5528 -1053 5562 -1019
rect 5596 -1053 5630 -1019
rect 5786 -1053 5820 -1019
rect 5854 -1053 5888 -1019
rect 625 -1334 659 -1300
rect 693 -1334 727 -1300
rect 883 -1334 917 -1300
rect 951 -1334 985 -1300
rect 5528 -1334 5562 -1300
rect 5596 -1334 5630 -1300
rect 5786 -1334 5820 -1300
rect 5854 -1334 5888 -1300
rect 625 -2557 659 -2523
rect 693 -2557 727 -2523
rect 883 -2557 917 -2523
rect 951 -2557 985 -2523
rect 5528 -2557 5562 -2523
rect 5596 -2557 5630 -2523
rect 5786 -2557 5820 -2523
rect 5854 -2557 5888 -2523
rect 625 -2838 659 -2804
rect 693 -2838 727 -2804
rect 883 -2838 917 -2804
rect 951 -2838 985 -2804
rect 5528 -2838 5562 -2804
rect 5596 -2838 5630 -2804
rect 5786 -2838 5820 -2804
rect 5854 -2838 5888 -2804
rect 625 -4061 659 -4027
rect 693 -4061 727 -4027
rect 883 -4061 917 -4027
rect 951 -4061 985 -4027
rect 5528 -4061 5562 -4027
rect 5596 -4061 5630 -4027
rect 5786 -4061 5820 -4027
rect 5854 -4061 5888 -4027
rect 625 -4342 659 -4308
rect 693 -4342 727 -4308
rect 883 -4342 917 -4308
rect 951 -4342 985 -4308
rect 5528 -4342 5562 -4308
rect 5596 -4342 5630 -4308
rect 5786 -4342 5820 -4308
rect 5854 -4342 5888 -4308
rect 625 -5417 659 -5383
rect 693 -5417 727 -5383
rect 883 -5417 917 -5383
rect 951 -5417 985 -5383
rect 1335 -5417 1369 -5383
rect 1403 -5417 1437 -5383
rect 1593 -5417 1627 -5383
rect 1661 -5417 1695 -5383
rect 1851 -5417 1885 -5383
rect 1919 -5417 1953 -5383
rect 2109 -5417 2143 -5383
rect 2177 -5417 2211 -5383
rect 2561 -5417 2595 -5383
rect 2629 -5417 2663 -5383
rect 2819 -5417 2853 -5383
rect 2887 -5417 2921 -5383
rect 3077 -5417 3111 -5383
rect 3145 -5417 3179 -5383
rect 3335 -5417 3369 -5383
rect 3403 -5417 3437 -5383
rect 3593 -5417 3627 -5383
rect 3661 -5417 3695 -5383
rect 3851 -5417 3885 -5383
rect 3919 -5417 3953 -5383
rect 4303 -5417 4337 -5383
rect 4371 -5417 4405 -5383
rect 4561 -5417 4595 -5383
rect 4629 -5417 4663 -5383
rect 4819 -5417 4853 -5383
rect 4887 -5417 4921 -5383
rect 5077 -5417 5111 -5383
rect 5145 -5417 5179 -5383
rect 5528 -5417 5562 -5383
rect 5596 -5417 5630 -5383
rect 5786 -5417 5820 -5383
rect 5854 -5417 5888 -5383
<< locali >>
rect 340 5922 461 5956
rect 521 5922 529 5956
rect 593 5922 597 5956
rect 699 5922 703 5956
rect 767 5922 775 5956
rect 835 5922 847 5956
rect 903 5922 919 5956
rect 971 5922 991 5956
rect 1039 5922 1063 5956
rect 1107 5922 1135 5956
rect 1175 5922 1207 5956
rect 1243 5922 1277 5956
rect 1313 5922 1345 5956
rect 1385 5922 1413 5956
rect 1457 5922 1481 5956
rect 1529 5922 1549 5956
rect 1601 5922 1617 5956
rect 1673 5922 1685 5956
rect 1745 5922 1753 5956
rect 1817 5922 1821 5956
rect 1923 5922 1927 5956
rect 1991 5922 1999 5956
rect 2059 5922 2071 5956
rect 2127 5922 2143 5956
rect 2195 5922 2215 5956
rect 2263 5922 2287 5956
rect 2331 5922 2359 5956
rect 2399 5922 2431 5956
rect 2467 5922 2501 5956
rect 2537 5922 2569 5956
rect 2609 5922 2637 5956
rect 2681 5922 2705 5956
rect 2753 5922 2773 5956
rect 2825 5922 2841 5956
rect 2897 5922 2909 5956
rect 2969 5922 2977 5956
rect 3041 5922 3045 5956
rect 3147 5922 3151 5956
rect 3215 5922 3223 5956
rect 3283 5922 3295 5956
rect 3351 5922 3367 5956
rect 3419 5922 3439 5956
rect 3487 5922 3511 5956
rect 3555 5922 3583 5956
rect 3623 5922 3655 5956
rect 3691 5922 3725 5956
rect 3761 5922 3793 5956
rect 3833 5922 3861 5956
rect 3905 5922 3929 5956
rect 3977 5922 3997 5956
rect 4049 5922 4065 5956
rect 4121 5922 4133 5956
rect 4193 5922 4201 5956
rect 4265 5922 4269 5956
rect 4371 5922 4375 5956
rect 4439 5922 4447 5956
rect 4507 5922 4519 5956
rect 4575 5922 4591 5956
rect 4643 5922 4663 5956
rect 4711 5922 4735 5956
rect 4779 5922 4807 5956
rect 4847 5922 4879 5956
rect 4915 5922 4949 5956
rect 4985 5922 5017 5956
rect 5057 5922 5085 5956
rect 5129 5922 5153 5956
rect 5201 5922 5221 5956
rect 5273 5922 5289 5956
rect 5345 5922 5357 5956
rect 5417 5922 5425 5956
rect 5489 5922 5493 5956
rect 5595 5922 5599 5956
rect 5663 5922 5671 5956
rect 5731 5922 5743 5956
rect 5799 5922 5815 5956
rect 5867 5922 5887 5956
rect 5935 5922 5959 5956
rect 6003 5922 6166 5956
rect 340 5821 374 5922
rect 6132 5821 6166 5922
rect 340 5749 374 5761
rect 340 5677 374 5693
rect 340 5605 374 5625
rect 530 5774 564 5793
rect 530 5706 564 5708
rect 530 5670 564 5672
rect 530 5585 564 5604
rect 788 5774 822 5793
rect 788 5706 822 5708
rect 788 5670 822 5672
rect 788 5585 822 5604
rect 1046 5774 1080 5793
rect 1046 5706 1080 5708
rect 1046 5670 1080 5672
rect 1046 5585 1080 5604
rect 1240 5774 1274 5793
rect 1240 5706 1274 5708
rect 1240 5670 1274 5672
rect 1240 5585 1274 5604
rect 1498 5774 1532 5793
rect 1498 5706 1532 5708
rect 1498 5670 1532 5672
rect 1498 5585 1532 5604
rect 1756 5774 1790 5793
rect 1756 5706 1790 5708
rect 1756 5670 1790 5672
rect 1756 5585 1790 5604
rect 2014 5774 2048 5793
rect 2014 5706 2048 5708
rect 2014 5670 2048 5672
rect 2014 5585 2048 5604
rect 2272 5774 2306 5793
rect 2272 5706 2306 5708
rect 2272 5670 2306 5672
rect 2272 5585 2306 5604
rect 2466 5774 2500 5793
rect 2466 5706 2500 5708
rect 2466 5670 2500 5672
rect 2466 5585 2500 5604
rect 2724 5774 2758 5793
rect 2724 5706 2758 5708
rect 2724 5670 2758 5672
rect 2724 5585 2758 5604
rect 2982 5774 3016 5793
rect 2982 5706 3016 5708
rect 2982 5670 3016 5672
rect 2982 5585 3016 5604
rect 3240 5774 3274 5793
rect 3240 5706 3274 5708
rect 3240 5670 3274 5672
rect 3240 5585 3274 5604
rect 3498 5774 3532 5793
rect 3498 5706 3532 5708
rect 3498 5670 3532 5672
rect 3498 5585 3532 5604
rect 3756 5774 3790 5793
rect 3756 5706 3790 5708
rect 3756 5670 3790 5672
rect 3756 5585 3790 5604
rect 4014 5774 4048 5793
rect 4014 5706 4048 5708
rect 4014 5670 4048 5672
rect 4014 5585 4048 5604
rect 4208 5774 4242 5793
rect 4208 5706 4242 5708
rect 4208 5670 4242 5672
rect 4208 5585 4242 5604
rect 4466 5774 4500 5793
rect 4466 5706 4500 5708
rect 4466 5670 4500 5672
rect 4466 5585 4500 5604
rect 4724 5774 4758 5793
rect 4724 5706 4758 5708
rect 4724 5670 4758 5672
rect 4724 5585 4758 5604
rect 4982 5774 5016 5793
rect 4982 5706 5016 5708
rect 4982 5670 5016 5672
rect 4982 5585 5016 5604
rect 5240 5774 5274 5793
rect 5240 5706 5274 5708
rect 5240 5670 5274 5672
rect 5240 5585 5274 5604
rect 5433 5774 5467 5793
rect 5433 5706 5467 5708
rect 5433 5670 5467 5672
rect 5433 5585 5467 5604
rect 5691 5774 5725 5793
rect 5691 5706 5725 5708
rect 5691 5670 5725 5672
rect 5691 5585 5725 5604
rect 5949 5774 5983 5793
rect 5949 5706 5983 5708
rect 5949 5670 5983 5672
rect 5949 5585 5983 5604
rect 6132 5749 6166 5761
rect 6132 5677 6166 5693
rect 6132 5605 6166 5625
rect 340 5533 374 5557
rect 576 5508 623 5542
rect 659 5508 693 5542
rect 729 5508 776 5542
rect 834 5508 881 5542
rect 917 5508 951 5542
rect 987 5508 1034 5542
rect 1286 5508 1333 5542
rect 1369 5508 1403 5542
rect 1439 5508 1486 5542
rect 1544 5508 1591 5542
rect 1627 5508 1661 5542
rect 1697 5508 1744 5542
rect 1802 5508 1849 5542
rect 1885 5508 1919 5542
rect 1955 5508 2002 5542
rect 2060 5508 2107 5542
rect 2143 5508 2177 5542
rect 2213 5508 2260 5542
rect 2512 5508 2559 5542
rect 2595 5508 2629 5542
rect 2665 5508 2712 5542
rect 2770 5508 2817 5542
rect 2853 5508 2887 5542
rect 2923 5508 2970 5542
rect 3028 5508 3075 5542
rect 3111 5508 3145 5542
rect 3181 5508 3228 5542
rect 3286 5508 3333 5542
rect 3369 5508 3403 5542
rect 3439 5508 3486 5542
rect 3544 5508 3591 5542
rect 3627 5508 3661 5542
rect 3697 5508 3744 5542
rect 3802 5508 3849 5542
rect 3885 5508 3919 5542
rect 3955 5508 4002 5542
rect 4254 5508 4301 5542
rect 4337 5508 4371 5542
rect 4407 5508 4454 5542
rect 4512 5508 4559 5542
rect 4595 5508 4629 5542
rect 4665 5508 4712 5542
rect 4770 5508 4817 5542
rect 4853 5508 4887 5542
rect 4923 5508 4970 5542
rect 5028 5508 5075 5542
rect 5111 5508 5145 5542
rect 5181 5508 5228 5542
rect 5479 5508 5526 5542
rect 5562 5508 5596 5542
rect 5632 5508 5679 5542
rect 5737 5508 5784 5542
rect 5820 5508 5854 5542
rect 5890 5508 5937 5542
rect 6132 5533 6166 5557
rect 340 5461 374 5489
rect 340 5389 374 5421
rect 340 5319 374 5353
rect 340 5251 374 5283
rect 6132 5461 6166 5489
rect 6132 5389 6166 5421
rect 6132 5319 6166 5353
rect 576 5227 623 5261
rect 659 5227 693 5261
rect 729 5227 776 5261
rect 834 5227 881 5261
rect 917 5227 951 5261
rect 987 5227 1034 5261
rect 5479 5227 5526 5261
rect 5562 5227 5596 5261
rect 5632 5227 5679 5261
rect 5737 5227 5784 5261
rect 5820 5227 5854 5261
rect 5890 5227 5937 5261
rect 6132 5251 6166 5283
rect 340 5183 374 5211
rect 340 5115 374 5139
rect 340 5047 374 5067
rect 340 4979 374 4995
rect 530 5165 564 5184
rect 530 5097 564 5099
rect 530 5061 564 5063
rect 530 4976 564 4995
rect 788 5165 822 5184
rect 788 5097 822 5099
rect 788 5061 822 5063
rect 788 4976 822 4995
rect 1046 5165 1080 5184
rect 1046 5097 1080 5099
rect 1046 5061 1080 5063
rect 1046 4976 1080 4995
rect 5433 5165 5467 5184
rect 5433 5097 5467 5099
rect 5433 5061 5467 5063
rect 5433 4976 5467 4995
rect 5691 5165 5725 5184
rect 5691 5097 5725 5099
rect 5691 5061 5725 5063
rect 5691 4976 5725 4995
rect 5949 5165 5983 5184
rect 5949 5097 5983 5099
rect 5949 5061 5983 5063
rect 5949 4976 5983 4995
rect 6132 5183 6166 5211
rect 6132 5115 6166 5139
rect 6132 5047 6166 5067
rect 6132 4979 6166 4995
rect 340 4911 374 4923
rect 340 4843 374 4851
rect 340 4775 374 4779
rect 340 4669 374 4673
rect 340 4597 374 4605
rect 340 4525 374 4537
rect 340 4453 374 4469
rect 340 4381 374 4401
rect 340 4309 374 4333
rect 6132 4911 6166 4923
rect 6132 4843 6166 4851
rect 6132 4775 6166 4779
rect 6132 4669 6166 4673
rect 6132 4597 6166 4605
rect 6132 4525 6166 4537
rect 6132 4453 6166 4469
rect 6132 4381 6166 4401
rect 6132 4309 6166 4333
rect 340 4237 374 4265
rect 340 4165 374 4197
rect 340 4095 374 4129
rect 530 4270 564 4289
rect 530 4202 564 4204
rect 530 4166 564 4168
rect 530 4081 564 4100
rect 788 4270 822 4289
rect 788 4202 822 4204
rect 788 4166 822 4168
rect 788 4081 822 4100
rect 1046 4270 1080 4289
rect 1046 4202 1080 4204
rect 1046 4166 1080 4168
rect 1046 4081 1080 4100
rect 5433 4270 5467 4289
rect 5433 4202 5467 4204
rect 5433 4166 5467 4168
rect 5433 4081 5467 4100
rect 5691 4270 5725 4289
rect 5691 4202 5725 4204
rect 5691 4166 5725 4168
rect 5691 4081 5725 4100
rect 5949 4270 5983 4289
rect 5949 4202 5983 4204
rect 5949 4166 5983 4168
rect 5949 4081 5983 4100
rect 6132 4237 6166 4265
rect 6132 4165 6166 4197
rect 6132 4095 6166 4129
rect 340 4027 374 4059
rect 576 4004 623 4038
rect 659 4004 693 4038
rect 729 4004 776 4038
rect 834 4004 881 4038
rect 917 4004 951 4038
rect 987 4004 1034 4038
rect 5479 4004 5526 4038
rect 5562 4004 5596 4038
rect 5632 4004 5679 4038
rect 5737 4004 5784 4038
rect 5820 4004 5854 4038
rect 5890 4004 5937 4038
rect 6132 4027 6166 4059
rect 340 3959 374 3987
rect 340 3891 374 3915
rect 340 3823 374 3843
rect 340 3755 374 3771
rect 6132 3959 6166 3987
rect 6132 3891 6166 3915
rect 6132 3823 6166 3843
rect 576 3723 623 3757
rect 659 3723 693 3757
rect 729 3723 776 3757
rect 834 3723 881 3757
rect 917 3723 951 3757
rect 987 3723 1034 3757
rect 5479 3723 5526 3757
rect 5562 3723 5596 3757
rect 5632 3723 5679 3757
rect 5737 3723 5784 3757
rect 5820 3723 5854 3757
rect 5890 3723 5937 3757
rect 6132 3755 6166 3771
rect 340 3687 374 3699
rect 6132 3687 6166 3699
rect 340 3619 374 3627
rect 340 3551 374 3555
rect 530 3661 564 3680
rect 530 3593 564 3595
rect 530 3557 564 3559
rect 530 3472 564 3491
rect 788 3661 822 3680
rect 788 3593 822 3595
rect 788 3557 822 3559
rect 788 3472 822 3491
rect 1046 3661 1080 3680
rect 1046 3593 1080 3595
rect 1046 3557 1080 3559
rect 1046 3472 1080 3491
rect 5433 3661 5467 3680
rect 5433 3593 5467 3595
rect 5433 3557 5467 3559
rect 5433 3472 5467 3491
rect 5691 3661 5725 3680
rect 5691 3593 5725 3595
rect 5691 3557 5725 3559
rect 5691 3472 5725 3491
rect 5949 3661 5983 3680
rect 5949 3593 5983 3595
rect 5949 3557 5983 3559
rect 5949 3472 5983 3491
rect 6132 3619 6166 3627
rect 6132 3551 6166 3555
rect 340 3445 374 3449
rect 340 3373 374 3381
rect 340 3301 374 3313
rect 340 3229 374 3245
rect 340 3157 374 3177
rect 340 3085 374 3109
rect 340 3013 374 3041
rect 340 2941 374 2973
rect 340 2871 374 2905
rect 340 2803 374 2835
rect 6132 3445 6166 3449
rect 6132 3373 6166 3381
rect 6132 3301 6166 3313
rect 6132 3229 6166 3245
rect 6132 3157 6166 3177
rect 6132 3085 6166 3109
rect 6132 3013 6166 3041
rect 6132 2941 6166 2973
rect 6132 2871 6166 2905
rect 6132 2803 6166 2835
rect 340 2735 374 2763
rect 340 2667 374 2691
rect 340 2599 374 2619
rect 530 2763 564 2782
rect 530 2695 564 2697
rect 530 2659 564 2661
rect 530 2574 564 2593
rect 788 2763 822 2782
rect 788 2695 822 2697
rect 788 2659 822 2661
rect 788 2574 822 2593
rect 1046 2763 1080 2782
rect 1046 2695 1080 2697
rect 1046 2659 1080 2661
rect 1046 2574 1080 2593
rect 5433 2763 5467 2782
rect 5433 2695 5467 2697
rect 5433 2659 5467 2661
rect 5433 2574 5467 2593
rect 5691 2763 5725 2782
rect 5691 2695 5725 2697
rect 5691 2659 5725 2661
rect 5691 2574 5725 2593
rect 5949 2763 5983 2782
rect 5949 2695 5983 2697
rect 5949 2659 5983 2661
rect 5949 2574 5983 2593
rect 6132 2735 6166 2763
rect 6132 2667 6166 2691
rect 6132 2599 6166 2619
rect 340 2531 374 2547
rect 6132 2531 6166 2547
rect 576 2497 623 2531
rect 659 2497 693 2531
rect 729 2497 776 2531
rect 834 2497 881 2531
rect 917 2497 951 2531
rect 987 2497 1034 2531
rect 5479 2497 5526 2531
rect 5562 2497 5596 2531
rect 5632 2497 5679 2531
rect 5737 2497 5784 2531
rect 5820 2497 5854 2531
rect 5890 2497 5937 2531
rect 340 2463 374 2475
rect 340 2395 374 2403
rect 340 2327 374 2331
rect 6132 2463 6166 2475
rect 6132 2395 6166 2403
rect 6132 2327 6166 2331
rect 340 2221 374 2225
rect 576 2216 623 2250
rect 659 2216 693 2250
rect 729 2216 776 2250
rect 834 2216 881 2250
rect 917 2216 951 2250
rect 987 2216 1034 2250
rect 5479 2216 5526 2250
rect 5562 2216 5596 2250
rect 5632 2216 5679 2250
rect 5737 2216 5784 2250
rect 5820 2216 5854 2250
rect 5890 2216 5937 2250
rect 6132 2221 6166 2225
rect 340 2149 374 2157
rect 340 2077 374 2089
rect 340 1928 374 2043
rect 530 2154 564 2173
rect 530 2086 564 2088
rect 530 2050 564 2052
rect 530 1965 564 1984
rect 788 2154 822 2173
rect 788 2086 822 2088
rect 788 2050 822 2052
rect 788 1965 822 1984
rect 1046 2154 1080 2173
rect 1046 2086 1080 2088
rect 1046 2050 1080 2052
rect 1046 1965 1080 1984
rect 5433 2154 5467 2173
rect 5433 2086 5467 2088
rect 5433 2050 5467 2052
rect 5433 1965 5467 1984
rect 5691 2154 5725 2173
rect 5691 2086 5725 2088
rect 5691 2050 5725 2052
rect 5691 1965 5725 1984
rect 5949 2154 5983 2173
rect 5949 2086 5983 2088
rect 5949 2050 5983 2052
rect 5949 1965 5983 1984
rect 6132 2149 6166 2157
rect 6132 2077 6166 2089
rect 340 1882 374 1894
rect 340 1814 374 1822
rect 340 1746 374 1750
rect 340 1640 374 1644
rect 340 1570 374 1576
rect 6132 1928 6166 2043
rect 6132 1882 6166 1894
rect 6132 1814 6166 1822
rect 6132 1746 6166 1750
rect 6132 1640 6166 1644
rect 6132 1570 6166 1576
rect 340 1568 6166 1570
rect 374 1536 6132 1568
rect 340 1496 374 1508
rect 340 1424 374 1440
rect 6132 1496 6166 1508
rect 6132 1424 6166 1440
rect 340 1352 374 1372
rect 340 1280 374 1304
rect 340 1208 374 1236
rect 530 1394 564 1413
rect 530 1326 564 1328
rect 530 1290 564 1292
rect 530 1205 564 1224
rect 788 1394 822 1413
rect 788 1326 822 1328
rect 788 1290 822 1292
rect 788 1205 822 1224
rect 1046 1394 1080 1413
rect 1046 1326 1080 1328
rect 1046 1290 1080 1292
rect 1046 1205 1080 1224
rect 5433 1394 5467 1413
rect 5433 1326 5467 1328
rect 5433 1290 5467 1292
rect 5433 1205 5467 1224
rect 5691 1394 5725 1413
rect 5691 1326 5725 1328
rect 5691 1290 5725 1292
rect 5691 1205 5725 1224
rect 5949 1394 5983 1413
rect 5949 1326 5983 1328
rect 5949 1290 5983 1292
rect 5949 1205 5983 1224
rect 6132 1352 6166 1372
rect 6132 1280 6166 1304
rect 6132 1208 6166 1236
rect 340 1136 374 1168
rect 576 1128 623 1162
rect 659 1128 693 1162
rect 729 1128 776 1162
rect 834 1128 881 1162
rect 917 1128 951 1162
rect 987 1128 1034 1162
rect 5479 1128 5526 1162
rect 5562 1128 5596 1162
rect 5632 1128 5679 1162
rect 5737 1128 5784 1162
rect 5820 1128 5854 1162
rect 5890 1128 5937 1162
rect 6132 1136 6166 1168
rect 340 1066 374 1100
rect 340 998 374 1030
rect 340 930 374 958
rect 340 862 374 886
rect 6132 1066 6166 1100
rect 6132 998 6166 1030
rect 6132 930 6166 958
rect 576 847 623 881
rect 659 847 693 881
rect 729 847 776 881
rect 834 847 881 881
rect 917 847 951 881
rect 987 847 1034 881
rect 5479 847 5526 881
rect 5562 847 5596 881
rect 5632 847 5679 881
rect 5737 847 5784 881
rect 5820 847 5854 881
rect 5890 847 5937 881
rect 6132 862 6166 886
rect 340 794 374 814
rect 340 726 374 742
rect 340 658 374 670
rect 340 590 374 598
rect 530 785 564 804
rect 530 717 564 719
rect 530 681 564 683
rect 530 596 564 615
rect 788 785 822 804
rect 788 717 822 719
rect 788 681 822 683
rect 788 596 822 615
rect 1046 785 1080 804
rect 1046 717 1080 719
rect 1046 681 1080 683
rect 1046 596 1080 615
rect 5433 785 5467 804
rect 5433 717 5467 719
rect 5433 681 5467 683
rect 5433 596 5467 615
rect 5691 785 5725 804
rect 5691 717 5725 719
rect 5691 681 5725 683
rect 5691 596 5725 615
rect 5949 785 5983 804
rect 5949 717 5983 719
rect 5949 681 5983 683
rect 5949 596 5983 615
rect 6132 794 6166 814
rect 6132 726 6166 742
rect 6132 658 6166 670
rect 340 522 374 526
rect 340 416 374 420
rect 340 344 374 352
rect 6132 590 6166 598
rect 6132 522 6166 526
rect 6132 416 6166 420
rect 6132 344 6166 352
rect 340 272 374 284
rect 340 200 374 216
rect 340 128 374 148
rect 530 299 564 318
rect 530 231 564 233
rect 530 195 564 197
rect 530 110 564 129
rect 788 299 822 318
rect 788 231 822 233
rect 788 195 822 197
rect 788 110 822 129
rect 1046 299 1080 318
rect 1046 231 1080 233
rect 1046 195 1080 197
rect 1046 110 1080 129
rect 5433 299 5467 318
rect 5433 231 5467 233
rect 5433 195 5467 197
rect 5433 110 5467 129
rect 5691 299 5725 318
rect 5691 231 5725 233
rect 5691 195 5725 197
rect 5691 110 5725 129
rect 5949 299 5983 318
rect 5949 231 5983 233
rect 5949 195 5983 197
rect 5949 110 5983 129
rect 6132 272 6166 284
rect 6132 200 6166 216
rect 6132 128 6166 148
rect 340 56 374 80
rect 576 33 623 67
rect 659 33 693 67
rect 729 33 776 67
rect 834 33 881 67
rect 917 33 951 67
rect 987 33 1034 67
rect 5479 33 5526 67
rect 5562 33 5596 67
rect 5632 33 5679 67
rect 5737 33 5784 67
rect 5820 33 5854 67
rect 5890 33 5937 67
rect 6132 56 6166 80
rect 340 -16 374 12
rect 340 -88 374 -56
rect 340 -158 374 -124
rect 340 -226 374 -194
rect 6132 -16 6166 12
rect 6132 -88 6166 -56
rect 6132 -158 6166 -124
rect 576 -248 623 -214
rect 659 -248 693 -214
rect 729 -248 776 -214
rect 834 -248 881 -214
rect 917 -248 951 -214
rect 987 -248 1034 -214
rect 5479 -248 5526 -214
rect 5562 -248 5596 -214
rect 5632 -248 5679 -214
rect 5737 -248 5784 -214
rect 5820 -248 5854 -214
rect 5890 -248 5937 -214
rect 6132 -226 6166 -194
rect 340 -294 374 -266
rect 340 -362 374 -338
rect 340 -430 374 -410
rect 340 -498 374 -482
rect 530 -310 564 -291
rect 530 -378 564 -376
rect 530 -414 564 -412
rect 530 -499 564 -480
rect 788 -310 822 -291
rect 788 -378 822 -376
rect 788 -414 822 -412
rect 788 -499 822 -480
rect 1046 -310 1080 -291
rect 1046 -378 1080 -376
rect 1046 -414 1080 -412
rect 1046 -499 1080 -480
rect 5433 -310 5467 -291
rect 5433 -378 5467 -376
rect 5433 -414 5467 -412
rect 5433 -499 5467 -480
rect 5691 -310 5725 -291
rect 5691 -378 5725 -376
rect 5691 -414 5725 -412
rect 5691 -499 5725 -480
rect 5949 -310 5983 -291
rect 5949 -378 5983 -376
rect 5949 -414 5983 -412
rect 5949 -499 5983 -480
rect 6132 -294 6166 -266
rect 6132 -362 6166 -338
rect 6132 -430 6166 -410
rect 6132 -498 6166 -482
rect 340 -566 374 -554
rect 340 -634 374 -626
rect 340 -702 374 -698
rect 6132 -566 6166 -554
rect 6132 -634 6166 -626
rect 6132 -702 6166 -698
rect 340 -808 374 -804
rect 340 -880 374 -872
rect 340 -952 374 -940
rect 530 -787 564 -768
rect 530 -855 564 -853
rect 530 -891 564 -889
rect 530 -976 564 -957
rect 788 -787 822 -768
rect 788 -855 822 -853
rect 788 -891 822 -889
rect 788 -976 822 -957
rect 1046 -787 1080 -768
rect 1046 -855 1080 -853
rect 1046 -891 1080 -889
rect 1046 -976 1080 -957
rect 5433 -787 5467 -768
rect 5433 -855 5467 -853
rect 5433 -891 5467 -889
rect 5433 -976 5467 -957
rect 5691 -787 5725 -768
rect 5691 -855 5725 -853
rect 5691 -891 5725 -889
rect 5691 -976 5725 -957
rect 5949 -787 5983 -768
rect 5949 -855 5983 -853
rect 5949 -891 5983 -889
rect 5949 -976 5983 -957
rect 6132 -808 6166 -804
rect 6132 -880 6166 -872
rect 6132 -952 6166 -940
rect 340 -1024 374 -1008
rect 576 -1053 623 -1019
rect 659 -1053 693 -1019
rect 729 -1053 776 -1019
rect 834 -1053 881 -1019
rect 917 -1053 951 -1019
rect 987 -1053 1034 -1019
rect 5479 -1053 5526 -1019
rect 5562 -1053 5596 -1019
rect 5632 -1053 5679 -1019
rect 5737 -1053 5784 -1019
rect 5820 -1053 5854 -1019
rect 5890 -1053 5937 -1019
rect 6132 -1024 6166 -1008
rect 340 -1096 374 -1076
rect 340 -1154 374 -1144
rect 6132 -1096 6166 -1076
rect 6132 -1154 6166 -1144
rect 340 -1168 6166 -1154
rect 374 -1188 6132 -1168
rect 340 -1240 374 -1212
rect 340 -1312 374 -1280
rect 6132 -1240 6166 -1212
rect 576 -1334 623 -1300
rect 659 -1334 693 -1300
rect 729 -1334 776 -1300
rect 834 -1334 881 -1300
rect 917 -1334 951 -1300
rect 987 -1334 1034 -1300
rect 5479 -1334 5526 -1300
rect 5562 -1334 5596 -1300
rect 5632 -1334 5679 -1300
rect 5737 -1334 5784 -1300
rect 5820 -1334 5854 -1300
rect 5890 -1334 5937 -1300
rect 6132 -1312 6166 -1280
rect 340 -1382 374 -1348
rect 340 -1450 374 -1418
rect 340 -1518 374 -1490
rect 340 -1586 374 -1562
rect 530 -1396 564 -1377
rect 530 -1464 564 -1462
rect 530 -1500 564 -1498
rect 530 -1585 564 -1566
rect 788 -1396 822 -1377
rect 788 -1464 822 -1462
rect 788 -1500 822 -1498
rect 788 -1585 822 -1566
rect 1046 -1396 1080 -1377
rect 1046 -1464 1080 -1462
rect 1046 -1500 1080 -1498
rect 1046 -1585 1080 -1566
rect 5433 -1396 5467 -1377
rect 5433 -1464 5467 -1462
rect 5433 -1500 5467 -1498
rect 5433 -1585 5467 -1566
rect 5691 -1396 5725 -1377
rect 5691 -1464 5725 -1462
rect 5691 -1500 5725 -1498
rect 5691 -1585 5725 -1566
rect 5949 -1396 5983 -1377
rect 5949 -1464 5983 -1462
rect 5949 -1500 5983 -1498
rect 5949 -1585 5983 -1566
rect 6132 -1382 6166 -1348
rect 6132 -1450 6166 -1418
rect 6132 -1518 6166 -1490
rect 340 -1654 374 -1634
rect 340 -1722 374 -1706
rect 340 -1790 374 -1778
rect 340 -1858 374 -1850
rect 340 -1926 374 -1922
rect 340 -2032 374 -2028
rect 340 -2104 374 -2096
rect 340 -2176 374 -2164
rect 340 -2248 374 -2232
rect 6132 -1586 6166 -1562
rect 6132 -1654 6166 -1634
rect 6132 -1722 6166 -1706
rect 6132 -1790 6166 -1778
rect 6132 -1858 6166 -1850
rect 6132 -1926 6166 -1922
rect 6132 -2032 6166 -2028
rect 6132 -2104 6166 -2096
rect 6132 -2176 6166 -2164
rect 6132 -2248 6166 -2232
rect 340 -2320 374 -2300
rect 340 -2392 374 -2368
rect 340 -2464 374 -2436
rect 530 -2291 564 -2272
rect 530 -2359 564 -2357
rect 530 -2395 564 -2393
rect 530 -2480 564 -2461
rect 788 -2291 822 -2272
rect 788 -2359 822 -2357
rect 788 -2395 822 -2393
rect 788 -2480 822 -2461
rect 1046 -2291 1080 -2272
rect 1046 -2359 1080 -2357
rect 1046 -2395 1080 -2393
rect 1046 -2480 1080 -2461
rect 5433 -2291 5467 -2272
rect 5433 -2359 5467 -2357
rect 5433 -2395 5467 -2393
rect 5433 -2480 5467 -2461
rect 5691 -2291 5725 -2272
rect 5691 -2359 5725 -2357
rect 5691 -2395 5725 -2393
rect 5691 -2480 5725 -2461
rect 5949 -2291 5983 -2272
rect 5949 -2359 5983 -2357
rect 5949 -2395 5983 -2393
rect 5949 -2480 5983 -2461
rect 6132 -2320 6166 -2300
rect 6132 -2392 6166 -2368
rect 6132 -2464 6166 -2436
rect 340 -2536 374 -2504
rect 576 -2557 623 -2523
rect 659 -2557 693 -2523
rect 729 -2557 776 -2523
rect 834 -2557 881 -2523
rect 917 -2557 951 -2523
rect 987 -2557 1034 -2523
rect 5479 -2557 5526 -2523
rect 5562 -2557 5596 -2523
rect 5632 -2557 5679 -2523
rect 5737 -2557 5784 -2523
rect 5820 -2557 5854 -2523
rect 5890 -2557 5937 -2523
rect 6132 -2536 6166 -2504
rect 340 -2606 374 -2572
rect 340 -2674 374 -2642
rect 340 -2742 374 -2714
rect 340 -2810 374 -2786
rect 6132 -2606 6166 -2572
rect 6132 -2674 6166 -2642
rect 6132 -2742 6166 -2714
rect 576 -2838 623 -2804
rect 659 -2838 693 -2804
rect 729 -2838 776 -2804
rect 834 -2838 881 -2804
rect 917 -2838 951 -2804
rect 987 -2838 1034 -2804
rect 5479 -2838 5526 -2804
rect 5562 -2838 5596 -2804
rect 5632 -2838 5679 -2804
rect 5737 -2838 5784 -2804
rect 5820 -2838 5854 -2804
rect 5890 -2838 5937 -2804
rect 6132 -2810 6166 -2786
rect 340 -2878 374 -2858
rect 6132 -2878 6166 -2858
rect 340 -2946 374 -2930
rect 340 -3014 374 -3002
rect 340 -3082 374 -3074
rect 530 -2900 564 -2881
rect 530 -2968 564 -2966
rect 530 -3004 564 -3002
rect 530 -3089 564 -3070
rect 788 -2900 822 -2881
rect 788 -2968 822 -2966
rect 788 -3004 822 -3002
rect 788 -3089 822 -3070
rect 1046 -2900 1080 -2881
rect 1046 -2968 1080 -2966
rect 1046 -3004 1080 -3002
rect 1046 -3089 1080 -3070
rect 5433 -2900 5467 -2881
rect 5433 -2968 5467 -2966
rect 5433 -3004 5467 -3002
rect 5433 -3089 5467 -3070
rect 5691 -2900 5725 -2881
rect 5691 -2968 5725 -2966
rect 5691 -3004 5725 -3002
rect 5691 -3089 5725 -3070
rect 5949 -2900 5983 -2881
rect 5949 -2968 5983 -2966
rect 5949 -3004 5983 -3002
rect 5949 -3089 5983 -3070
rect 6132 -2946 6166 -2930
rect 6132 -3014 6166 -3002
rect 6132 -3082 6166 -3074
rect 340 -3150 374 -3146
rect 340 -3256 374 -3252
rect 340 -3328 374 -3320
rect 340 -3400 374 -3388
rect 340 -3472 374 -3456
rect 340 -3544 374 -3524
rect 340 -3616 374 -3592
rect 340 -3688 374 -3660
rect 340 -3760 374 -3728
rect 6132 -3150 6166 -3146
rect 6132 -3256 6166 -3252
rect 6132 -3328 6166 -3320
rect 6132 -3400 6166 -3388
rect 6132 -3472 6166 -3456
rect 6132 -3544 6166 -3524
rect 6132 -3616 6166 -3592
rect 6132 -3688 6166 -3660
rect 6132 -3760 6166 -3728
rect 340 -3830 374 -3796
rect 340 -3898 374 -3866
rect 340 -3966 374 -3938
rect 530 -3795 564 -3776
rect 530 -3863 564 -3861
rect 530 -3899 564 -3897
rect 530 -3984 564 -3965
rect 788 -3795 822 -3776
rect 788 -3863 822 -3861
rect 788 -3899 822 -3897
rect 788 -3984 822 -3965
rect 1046 -3795 1080 -3776
rect 1046 -3863 1080 -3861
rect 1046 -3899 1080 -3897
rect 1046 -3984 1080 -3965
rect 5433 -3795 5467 -3776
rect 5433 -3863 5467 -3861
rect 5433 -3899 5467 -3897
rect 5433 -3984 5467 -3965
rect 5691 -3795 5725 -3776
rect 5691 -3863 5725 -3861
rect 5691 -3899 5725 -3897
rect 5691 -3984 5725 -3965
rect 5949 -3795 5983 -3776
rect 5949 -3863 5983 -3861
rect 5949 -3899 5983 -3897
rect 5949 -3984 5983 -3965
rect 6132 -3830 6166 -3796
rect 6132 -3898 6166 -3866
rect 6132 -3966 6166 -3938
rect 340 -4034 374 -4010
rect 576 -4061 623 -4027
rect 659 -4061 693 -4027
rect 729 -4061 776 -4027
rect 834 -4061 881 -4027
rect 917 -4061 951 -4027
rect 987 -4061 1034 -4027
rect 5479 -4061 5526 -4027
rect 5562 -4061 5596 -4027
rect 5632 -4061 5679 -4027
rect 5737 -4061 5784 -4027
rect 5820 -4061 5854 -4027
rect 5890 -4061 5937 -4027
rect 6132 -4034 6166 -4010
rect 340 -4102 374 -4082
rect 340 -4170 374 -4154
rect 340 -4238 374 -4226
rect 340 -4306 374 -4298
rect 6132 -4102 6166 -4082
rect 6132 -4170 6166 -4154
rect 6132 -4238 6166 -4226
rect 6132 -4306 6166 -4298
rect 576 -4342 623 -4308
rect 659 -4342 693 -4308
rect 729 -4342 776 -4308
rect 834 -4342 881 -4308
rect 917 -4342 951 -4308
rect 987 -4342 1034 -4308
rect 5479 -4342 5526 -4308
rect 5562 -4342 5596 -4308
rect 5632 -4342 5679 -4308
rect 5737 -4342 5784 -4308
rect 5820 -4342 5854 -4308
rect 5890 -4342 5937 -4308
rect 340 -4374 374 -4370
rect 6132 -4374 6166 -4370
rect 340 -4480 374 -4476
rect 340 -4552 374 -4544
rect 530 -4404 564 -4385
rect 530 -4472 564 -4470
rect 530 -4508 564 -4506
rect 530 -4593 564 -4574
rect 788 -4404 822 -4385
rect 788 -4472 822 -4470
rect 788 -4508 822 -4506
rect 788 -4593 822 -4574
rect 1046 -4404 1080 -4385
rect 1046 -4472 1080 -4470
rect 1046 -4508 1080 -4506
rect 1046 -4593 1080 -4574
rect 5433 -4404 5467 -4385
rect 5433 -4472 5467 -4470
rect 5433 -4508 5467 -4506
rect 5433 -4593 5467 -4574
rect 5691 -4404 5725 -4385
rect 5691 -4472 5725 -4470
rect 5691 -4508 5725 -4506
rect 5691 -4593 5725 -4574
rect 5949 -4404 5983 -4385
rect 5949 -4472 5983 -4470
rect 5949 -4508 5983 -4506
rect 5949 -4593 5983 -4574
rect 6132 -4480 6166 -4476
rect 6132 -4552 6166 -4544
rect 340 -4624 374 -4612
rect 340 -4696 374 -4680
rect 340 -4768 374 -4748
rect 340 -4840 374 -4816
rect 340 -4912 374 -4884
rect 340 -4984 374 -4952
rect 340 -5054 374 -5020
rect 340 -5122 374 -5090
rect 6132 -4624 6166 -4612
rect 6132 -4696 6166 -4680
rect 6132 -4768 6166 -4748
rect 6132 -4840 6166 -4816
rect 6132 -4912 6166 -4884
rect 6132 -4984 6166 -4952
rect 6132 -5054 6166 -5020
rect 6132 -5122 6166 -5090
rect 340 -5190 374 -5162
rect 340 -5258 374 -5234
rect 340 -5326 374 -5306
rect 530 -5151 564 -5132
rect 530 -5219 564 -5217
rect 530 -5255 564 -5253
rect 530 -5340 564 -5321
rect 788 -5151 822 -5132
rect 788 -5219 822 -5217
rect 788 -5255 822 -5253
rect 788 -5340 822 -5321
rect 1046 -5151 1080 -5132
rect 1046 -5219 1080 -5217
rect 1046 -5255 1080 -5253
rect 1046 -5340 1080 -5321
rect 1240 -5151 1274 -5132
rect 1240 -5219 1274 -5217
rect 1240 -5255 1274 -5253
rect 1240 -5340 1274 -5321
rect 1498 -5151 1532 -5132
rect 1498 -5219 1532 -5217
rect 1498 -5255 1532 -5253
rect 1498 -5340 1532 -5321
rect 1756 -5151 1790 -5132
rect 1756 -5219 1790 -5217
rect 1756 -5255 1790 -5253
rect 1756 -5340 1790 -5321
rect 2014 -5151 2048 -5132
rect 2014 -5219 2048 -5217
rect 2014 -5255 2048 -5253
rect 2014 -5340 2048 -5321
rect 2272 -5151 2306 -5132
rect 2272 -5219 2306 -5217
rect 2272 -5255 2306 -5253
rect 2272 -5340 2306 -5321
rect 2466 -5151 2500 -5132
rect 2466 -5219 2500 -5217
rect 2466 -5255 2500 -5253
rect 2466 -5340 2500 -5321
rect 2724 -5151 2758 -5132
rect 2724 -5219 2758 -5217
rect 2724 -5255 2758 -5253
rect 2724 -5340 2758 -5321
rect 2982 -5151 3016 -5132
rect 2982 -5219 3016 -5217
rect 2982 -5255 3016 -5253
rect 2982 -5340 3016 -5321
rect 3240 -5151 3274 -5132
rect 3240 -5219 3274 -5217
rect 3240 -5255 3274 -5253
rect 3240 -5340 3274 -5321
rect 3498 -5151 3532 -5132
rect 3498 -5219 3532 -5217
rect 3498 -5255 3532 -5253
rect 3498 -5340 3532 -5321
rect 3756 -5151 3790 -5132
rect 3756 -5219 3790 -5217
rect 3756 -5255 3790 -5253
rect 3756 -5340 3790 -5321
rect 4014 -5151 4048 -5132
rect 4014 -5219 4048 -5217
rect 4014 -5255 4048 -5253
rect 4014 -5340 4048 -5321
rect 4208 -5151 4242 -5132
rect 4208 -5219 4242 -5217
rect 4208 -5255 4242 -5253
rect 4208 -5340 4242 -5321
rect 4466 -5151 4500 -5132
rect 4466 -5219 4500 -5217
rect 4466 -5255 4500 -5253
rect 4466 -5340 4500 -5321
rect 4724 -5151 4758 -5132
rect 4724 -5219 4758 -5217
rect 4724 -5255 4758 -5253
rect 4724 -5340 4758 -5321
rect 4982 -5151 5016 -5132
rect 4982 -5219 5016 -5217
rect 4982 -5255 5016 -5253
rect 4982 -5340 5016 -5321
rect 5240 -5151 5274 -5132
rect 5240 -5219 5274 -5217
rect 5240 -5255 5274 -5253
rect 5240 -5340 5274 -5321
rect 5433 -5151 5467 -5132
rect 5433 -5219 5467 -5217
rect 5433 -5255 5467 -5253
rect 5433 -5340 5467 -5321
rect 5691 -5151 5725 -5132
rect 5691 -5219 5725 -5217
rect 5691 -5255 5725 -5253
rect 5691 -5340 5725 -5321
rect 5949 -5151 5983 -5132
rect 5949 -5219 5983 -5217
rect 5949 -5255 5983 -5253
rect 5949 -5340 5983 -5321
rect 6132 -5190 6166 -5162
rect 6132 -5258 6166 -5234
rect 6132 -5326 6166 -5306
rect 340 -5506 374 -5378
rect 576 -5417 623 -5383
rect 659 -5417 693 -5383
rect 729 -5417 776 -5383
rect 834 -5417 881 -5383
rect 917 -5417 951 -5383
rect 987 -5417 1034 -5383
rect 1286 -5417 1333 -5383
rect 1369 -5417 1403 -5383
rect 1439 -5417 1486 -5383
rect 1544 -5417 1591 -5383
rect 1627 -5417 1661 -5383
rect 1697 -5417 1744 -5383
rect 1802 -5417 1849 -5383
rect 1885 -5417 1919 -5383
rect 1955 -5417 2002 -5383
rect 2060 -5417 2107 -5383
rect 2143 -5417 2177 -5383
rect 2213 -5417 2260 -5383
rect 2512 -5417 2559 -5383
rect 2595 -5417 2629 -5383
rect 2665 -5417 2712 -5383
rect 2770 -5417 2817 -5383
rect 2853 -5417 2887 -5383
rect 2923 -5417 2970 -5383
rect 3028 -5417 3075 -5383
rect 3111 -5417 3145 -5383
rect 3181 -5417 3228 -5383
rect 3286 -5417 3333 -5383
rect 3369 -5417 3403 -5383
rect 3439 -5417 3486 -5383
rect 3544 -5417 3591 -5383
rect 3627 -5417 3661 -5383
rect 3697 -5417 3744 -5383
rect 3802 -5417 3849 -5383
rect 3885 -5417 3919 -5383
rect 3955 -5417 4002 -5383
rect 4254 -5417 4301 -5383
rect 4337 -5417 4371 -5383
rect 4407 -5417 4454 -5383
rect 4512 -5417 4559 -5383
rect 4595 -5417 4629 -5383
rect 4665 -5417 4712 -5383
rect 4770 -5417 4817 -5383
rect 4853 -5417 4887 -5383
rect 4923 -5417 4970 -5383
rect 5028 -5417 5075 -5383
rect 5111 -5417 5145 -5383
rect 5181 -5417 5228 -5383
rect 5479 -5417 5526 -5383
rect 5562 -5417 5596 -5383
rect 5632 -5417 5679 -5383
rect 5737 -5417 5784 -5383
rect 5820 -5417 5854 -5383
rect 5890 -5417 5937 -5383
rect 6132 -5506 6166 -5378
rect 340 -5540 461 -5506
rect 521 -5540 529 -5506
rect 593 -5540 597 -5506
rect 699 -5540 703 -5506
rect 767 -5540 775 -5506
rect 835 -5540 847 -5506
rect 903 -5540 919 -5506
rect 971 -5540 991 -5506
rect 1039 -5540 1063 -5506
rect 1107 -5540 1135 -5506
rect 1175 -5540 1207 -5506
rect 1243 -5540 1277 -5506
rect 1313 -5540 1345 -5506
rect 1385 -5540 1413 -5506
rect 1457 -5540 1481 -5506
rect 1529 -5540 1549 -5506
rect 1601 -5540 1617 -5506
rect 1673 -5540 1685 -5506
rect 1745 -5540 1753 -5506
rect 1817 -5540 1821 -5506
rect 1923 -5540 1927 -5506
rect 1991 -5540 1999 -5506
rect 2059 -5540 2071 -5506
rect 2127 -5540 2143 -5506
rect 2195 -5540 2215 -5506
rect 2263 -5540 2287 -5506
rect 2331 -5540 2359 -5506
rect 2399 -5540 2431 -5506
rect 2467 -5540 2501 -5506
rect 2537 -5540 2569 -5506
rect 2609 -5540 2637 -5506
rect 2681 -5540 2705 -5506
rect 2753 -5540 2773 -5506
rect 2825 -5540 2841 -5506
rect 2897 -5540 2909 -5506
rect 2969 -5540 2977 -5506
rect 3041 -5540 3045 -5506
rect 3147 -5540 3151 -5506
rect 3215 -5540 3223 -5506
rect 3283 -5540 3295 -5506
rect 3351 -5540 3367 -5506
rect 3419 -5540 3439 -5506
rect 3487 -5540 3511 -5506
rect 3555 -5540 3583 -5506
rect 3623 -5540 3655 -5506
rect 3691 -5540 3725 -5506
rect 3761 -5540 3793 -5506
rect 3833 -5540 3861 -5506
rect 3905 -5540 3929 -5506
rect 3977 -5540 3997 -5506
rect 4049 -5540 4065 -5506
rect 4121 -5540 4133 -5506
rect 4193 -5540 4201 -5506
rect 4265 -5540 4269 -5506
rect 4371 -5540 4375 -5506
rect 4439 -5540 4447 -5506
rect 4507 -5540 4519 -5506
rect 4575 -5540 4591 -5506
rect 4643 -5540 4663 -5506
rect 4711 -5540 4735 -5506
rect 4779 -5540 4807 -5506
rect 4847 -5540 4879 -5506
rect 4915 -5540 4949 -5506
rect 4985 -5540 5017 -5506
rect 5057 -5540 5085 -5506
rect 5129 -5540 5153 -5506
rect 5201 -5540 5221 -5506
rect 5273 -5540 5289 -5506
rect 5345 -5540 5357 -5506
rect 5417 -5540 5425 -5506
rect 5489 -5540 5493 -5506
rect 5595 -5540 5599 -5506
rect 5663 -5540 5671 -5506
rect 5731 -5540 5743 -5506
rect 5799 -5540 5815 -5506
rect 5867 -5540 5887 -5506
rect 5935 -5540 5959 -5506
rect 6003 -5540 6166 -5506
<< viali >>
rect 487 5922 495 5956
rect 495 5922 521 5956
rect 559 5922 563 5956
rect 563 5922 593 5956
rect 631 5922 665 5956
rect 703 5922 733 5956
rect 733 5922 737 5956
rect 775 5922 801 5956
rect 801 5922 809 5956
rect 847 5922 869 5956
rect 869 5922 881 5956
rect 919 5922 937 5956
rect 937 5922 953 5956
rect 991 5922 1005 5956
rect 1005 5922 1025 5956
rect 1063 5922 1073 5956
rect 1073 5922 1097 5956
rect 1135 5922 1141 5956
rect 1141 5922 1169 5956
rect 1207 5922 1209 5956
rect 1209 5922 1241 5956
rect 1279 5922 1311 5956
rect 1311 5922 1313 5956
rect 1351 5922 1379 5956
rect 1379 5922 1385 5956
rect 1423 5922 1447 5956
rect 1447 5922 1457 5956
rect 1495 5922 1515 5956
rect 1515 5922 1529 5956
rect 1567 5922 1583 5956
rect 1583 5922 1601 5956
rect 1639 5922 1651 5956
rect 1651 5922 1673 5956
rect 1711 5922 1719 5956
rect 1719 5922 1745 5956
rect 1783 5922 1787 5956
rect 1787 5922 1817 5956
rect 1855 5922 1889 5956
rect 1927 5922 1957 5956
rect 1957 5922 1961 5956
rect 1999 5922 2025 5956
rect 2025 5922 2033 5956
rect 2071 5922 2093 5956
rect 2093 5922 2105 5956
rect 2143 5922 2161 5956
rect 2161 5922 2177 5956
rect 2215 5922 2229 5956
rect 2229 5922 2249 5956
rect 2287 5922 2297 5956
rect 2297 5922 2321 5956
rect 2359 5922 2365 5956
rect 2365 5922 2393 5956
rect 2431 5922 2433 5956
rect 2433 5922 2465 5956
rect 2503 5922 2535 5956
rect 2535 5922 2537 5956
rect 2575 5922 2603 5956
rect 2603 5922 2609 5956
rect 2647 5922 2671 5956
rect 2671 5922 2681 5956
rect 2719 5922 2739 5956
rect 2739 5922 2753 5956
rect 2791 5922 2807 5956
rect 2807 5922 2825 5956
rect 2863 5922 2875 5956
rect 2875 5922 2897 5956
rect 2935 5922 2943 5956
rect 2943 5922 2969 5956
rect 3007 5922 3011 5956
rect 3011 5922 3041 5956
rect 3079 5922 3113 5956
rect 3151 5922 3181 5956
rect 3181 5922 3185 5956
rect 3223 5922 3249 5956
rect 3249 5922 3257 5956
rect 3295 5922 3317 5956
rect 3317 5922 3329 5956
rect 3367 5922 3385 5956
rect 3385 5922 3401 5956
rect 3439 5922 3453 5956
rect 3453 5922 3473 5956
rect 3511 5922 3521 5956
rect 3521 5922 3545 5956
rect 3583 5922 3589 5956
rect 3589 5922 3617 5956
rect 3655 5922 3657 5956
rect 3657 5922 3689 5956
rect 3727 5922 3759 5956
rect 3759 5922 3761 5956
rect 3799 5922 3827 5956
rect 3827 5922 3833 5956
rect 3871 5922 3895 5956
rect 3895 5922 3905 5956
rect 3943 5922 3963 5956
rect 3963 5922 3977 5956
rect 4015 5922 4031 5956
rect 4031 5922 4049 5956
rect 4087 5922 4099 5956
rect 4099 5922 4121 5956
rect 4159 5922 4167 5956
rect 4167 5922 4193 5956
rect 4231 5922 4235 5956
rect 4235 5922 4265 5956
rect 4303 5922 4337 5956
rect 4375 5922 4405 5956
rect 4405 5922 4409 5956
rect 4447 5922 4473 5956
rect 4473 5922 4481 5956
rect 4519 5922 4541 5956
rect 4541 5922 4553 5956
rect 4591 5922 4609 5956
rect 4609 5922 4625 5956
rect 4663 5922 4677 5956
rect 4677 5922 4697 5956
rect 4735 5922 4745 5956
rect 4745 5922 4769 5956
rect 4807 5922 4813 5956
rect 4813 5922 4841 5956
rect 4879 5922 4881 5956
rect 4881 5922 4913 5956
rect 4951 5922 4983 5956
rect 4983 5922 4985 5956
rect 5023 5922 5051 5956
rect 5051 5922 5057 5956
rect 5095 5922 5119 5956
rect 5119 5922 5129 5956
rect 5167 5922 5187 5956
rect 5187 5922 5201 5956
rect 5239 5922 5255 5956
rect 5255 5922 5273 5956
rect 5311 5922 5323 5956
rect 5323 5922 5345 5956
rect 5383 5922 5391 5956
rect 5391 5922 5417 5956
rect 5455 5922 5459 5956
rect 5459 5922 5489 5956
rect 5527 5922 5561 5956
rect 5599 5922 5629 5956
rect 5629 5922 5633 5956
rect 5671 5922 5697 5956
rect 5697 5922 5705 5956
rect 5743 5922 5765 5956
rect 5765 5922 5777 5956
rect 5815 5922 5833 5956
rect 5833 5922 5849 5956
rect 5887 5922 5901 5956
rect 5901 5922 5921 5956
rect 5959 5922 5969 5956
rect 5969 5922 5993 5956
rect 340 5795 374 5821
rect 340 5787 374 5795
rect 6132 5795 6166 5821
rect 340 5727 374 5749
rect 340 5715 374 5727
rect 340 5659 374 5677
rect 340 5643 374 5659
rect 340 5591 374 5605
rect 340 5571 374 5591
rect 530 5740 564 5742
rect 530 5708 564 5740
rect 530 5638 564 5670
rect 530 5636 564 5638
rect 788 5740 822 5742
rect 788 5708 822 5740
rect 788 5638 822 5670
rect 788 5636 822 5638
rect 1046 5740 1080 5742
rect 1046 5708 1080 5740
rect 1046 5638 1080 5670
rect 1046 5636 1080 5638
rect 1240 5740 1274 5742
rect 1240 5708 1274 5740
rect 1240 5638 1274 5670
rect 1240 5636 1274 5638
rect 1498 5740 1532 5742
rect 1498 5708 1532 5740
rect 1498 5638 1532 5670
rect 1498 5636 1532 5638
rect 1756 5740 1790 5742
rect 1756 5708 1790 5740
rect 1756 5638 1790 5670
rect 1756 5636 1790 5638
rect 2014 5740 2048 5742
rect 2014 5708 2048 5740
rect 2014 5638 2048 5670
rect 2014 5636 2048 5638
rect 2272 5740 2306 5742
rect 2272 5708 2306 5740
rect 2272 5638 2306 5670
rect 2272 5636 2306 5638
rect 2466 5740 2500 5742
rect 2466 5708 2500 5740
rect 2466 5638 2500 5670
rect 2466 5636 2500 5638
rect 2724 5740 2758 5742
rect 2724 5708 2758 5740
rect 2724 5638 2758 5670
rect 2724 5636 2758 5638
rect 2982 5740 3016 5742
rect 2982 5708 3016 5740
rect 2982 5638 3016 5670
rect 2982 5636 3016 5638
rect 3240 5740 3274 5742
rect 3240 5708 3274 5740
rect 3240 5638 3274 5670
rect 3240 5636 3274 5638
rect 3498 5740 3532 5742
rect 3498 5708 3532 5740
rect 3498 5638 3532 5670
rect 3498 5636 3532 5638
rect 3756 5740 3790 5742
rect 3756 5708 3790 5740
rect 3756 5638 3790 5670
rect 3756 5636 3790 5638
rect 4014 5740 4048 5742
rect 4014 5708 4048 5740
rect 4014 5638 4048 5670
rect 4014 5636 4048 5638
rect 4208 5740 4242 5742
rect 4208 5708 4242 5740
rect 4208 5638 4242 5670
rect 4208 5636 4242 5638
rect 4466 5740 4500 5742
rect 4466 5708 4500 5740
rect 4466 5638 4500 5670
rect 4466 5636 4500 5638
rect 4724 5740 4758 5742
rect 4724 5708 4758 5740
rect 4724 5638 4758 5670
rect 4724 5636 4758 5638
rect 4982 5740 5016 5742
rect 4982 5708 5016 5740
rect 4982 5638 5016 5670
rect 4982 5636 5016 5638
rect 5240 5740 5274 5742
rect 5240 5708 5274 5740
rect 5240 5638 5274 5670
rect 5240 5636 5274 5638
rect 5433 5740 5467 5742
rect 5433 5708 5467 5740
rect 5433 5638 5467 5670
rect 5433 5636 5467 5638
rect 5691 5740 5725 5742
rect 5691 5708 5725 5740
rect 5691 5638 5725 5670
rect 5691 5636 5725 5638
rect 5949 5740 5983 5742
rect 5949 5708 5983 5740
rect 5949 5638 5983 5670
rect 5949 5636 5983 5638
rect 6132 5787 6166 5795
rect 6132 5727 6166 5749
rect 6132 5715 6166 5727
rect 6132 5659 6166 5677
rect 6132 5643 6166 5659
rect 6132 5591 6166 5605
rect 6132 5571 6166 5591
rect 340 5523 374 5533
rect 340 5499 374 5523
rect 623 5508 625 5542
rect 625 5508 657 5542
rect 695 5508 727 5542
rect 727 5508 729 5542
rect 881 5508 883 5542
rect 883 5508 915 5542
rect 953 5508 985 5542
rect 985 5508 987 5542
rect 1333 5508 1335 5542
rect 1335 5508 1367 5542
rect 1405 5508 1437 5542
rect 1437 5508 1439 5542
rect 1591 5508 1593 5542
rect 1593 5508 1625 5542
rect 1663 5508 1695 5542
rect 1695 5508 1697 5542
rect 1849 5508 1851 5542
rect 1851 5508 1883 5542
rect 1921 5508 1953 5542
rect 1953 5508 1955 5542
rect 2107 5508 2109 5542
rect 2109 5508 2141 5542
rect 2179 5508 2211 5542
rect 2211 5508 2213 5542
rect 2559 5508 2561 5542
rect 2561 5508 2593 5542
rect 2631 5508 2663 5542
rect 2663 5508 2665 5542
rect 2817 5508 2819 5542
rect 2819 5508 2851 5542
rect 2889 5508 2921 5542
rect 2921 5508 2923 5542
rect 3075 5508 3077 5542
rect 3077 5508 3109 5542
rect 3147 5508 3179 5542
rect 3179 5508 3181 5542
rect 3333 5508 3335 5542
rect 3335 5508 3367 5542
rect 3405 5508 3437 5542
rect 3437 5508 3439 5542
rect 3591 5508 3593 5542
rect 3593 5508 3625 5542
rect 3663 5508 3695 5542
rect 3695 5508 3697 5542
rect 3849 5508 3851 5542
rect 3851 5508 3883 5542
rect 3921 5508 3953 5542
rect 3953 5508 3955 5542
rect 4301 5508 4303 5542
rect 4303 5508 4335 5542
rect 4373 5508 4405 5542
rect 4405 5508 4407 5542
rect 4559 5508 4561 5542
rect 4561 5508 4593 5542
rect 4631 5508 4663 5542
rect 4663 5508 4665 5542
rect 4817 5508 4819 5542
rect 4819 5508 4851 5542
rect 4889 5508 4921 5542
rect 4921 5508 4923 5542
rect 5075 5508 5077 5542
rect 5077 5508 5109 5542
rect 5147 5508 5179 5542
rect 5179 5508 5181 5542
rect 5526 5508 5528 5542
rect 5528 5508 5560 5542
rect 5598 5508 5630 5542
rect 5630 5508 5632 5542
rect 5784 5508 5786 5542
rect 5786 5508 5818 5542
rect 5856 5508 5888 5542
rect 5888 5508 5890 5542
rect 6132 5523 6166 5533
rect 340 5455 374 5461
rect 340 5427 374 5455
rect 340 5387 374 5389
rect 340 5355 374 5387
rect 340 5285 374 5317
rect 340 5283 374 5285
rect 6132 5499 6166 5523
rect 6132 5455 6166 5461
rect 6132 5427 6166 5455
rect 6132 5387 6166 5389
rect 6132 5355 6166 5387
rect 6132 5285 6166 5317
rect 6132 5283 6166 5285
rect 340 5217 374 5245
rect 623 5227 625 5261
rect 625 5227 657 5261
rect 695 5227 727 5261
rect 727 5227 729 5261
rect 881 5227 883 5261
rect 883 5227 915 5261
rect 953 5227 985 5261
rect 985 5227 987 5261
rect 5526 5227 5528 5261
rect 5528 5227 5560 5261
rect 5598 5227 5630 5261
rect 5630 5227 5632 5261
rect 5784 5227 5786 5261
rect 5786 5227 5818 5261
rect 5856 5227 5888 5261
rect 5888 5227 5890 5261
rect 340 5211 374 5217
rect 6132 5217 6166 5245
rect 6132 5211 6166 5217
rect 340 5149 374 5173
rect 340 5139 374 5149
rect 340 5081 374 5101
rect 340 5067 374 5081
rect 340 5013 374 5029
rect 340 4995 374 5013
rect 530 5131 564 5133
rect 530 5099 564 5131
rect 530 5029 564 5061
rect 530 5027 564 5029
rect 788 5131 822 5133
rect 788 5099 822 5131
rect 788 5029 822 5061
rect 788 5027 822 5029
rect 1046 5131 1080 5133
rect 1046 5099 1080 5131
rect 1046 5029 1080 5061
rect 1046 5027 1080 5029
rect 5433 5131 5467 5133
rect 5433 5099 5467 5131
rect 5433 5029 5467 5061
rect 5433 5027 5467 5029
rect 5691 5131 5725 5133
rect 5691 5099 5725 5131
rect 5691 5029 5725 5061
rect 5691 5027 5725 5029
rect 5949 5131 5983 5133
rect 5949 5099 5983 5131
rect 5949 5029 5983 5061
rect 5949 5027 5983 5029
rect 6132 5149 6166 5173
rect 6132 5139 6166 5149
rect 6132 5081 6166 5101
rect 6132 5067 6166 5081
rect 6132 5013 6166 5029
rect 6132 4995 6166 5013
rect 340 4945 374 4957
rect 340 4923 374 4945
rect 340 4877 374 4885
rect 340 4851 374 4877
rect 340 4809 374 4813
rect 340 4779 374 4809
rect 340 4707 374 4741
rect 340 4639 374 4669
rect 340 4635 374 4639
rect 340 4571 374 4597
rect 340 4563 374 4571
rect 340 4503 374 4525
rect 340 4491 374 4503
rect 340 4435 374 4453
rect 340 4419 374 4435
rect 340 4367 374 4381
rect 340 4347 374 4367
rect 340 4299 374 4309
rect 340 4275 374 4299
rect 6132 4945 6166 4957
rect 6132 4923 6166 4945
rect 6132 4877 6166 4885
rect 6132 4851 6166 4877
rect 6132 4809 6166 4813
rect 6132 4779 6166 4809
rect 6132 4707 6166 4741
rect 6132 4639 6166 4669
rect 6132 4635 6166 4639
rect 6132 4571 6166 4597
rect 6132 4563 6166 4571
rect 6132 4503 6166 4525
rect 6132 4491 6166 4503
rect 6132 4435 6166 4453
rect 6132 4419 6166 4435
rect 6132 4367 6166 4381
rect 6132 4347 6166 4367
rect 6132 4299 6166 4309
rect 340 4231 374 4237
rect 340 4203 374 4231
rect 340 4163 374 4165
rect 340 4131 374 4163
rect 340 4061 374 4093
rect 530 4236 564 4238
rect 530 4204 564 4236
rect 530 4134 564 4166
rect 530 4132 564 4134
rect 788 4236 822 4238
rect 788 4204 822 4236
rect 788 4134 822 4166
rect 788 4132 822 4134
rect 1046 4236 1080 4238
rect 1046 4204 1080 4236
rect 1046 4134 1080 4166
rect 1046 4132 1080 4134
rect 5433 4236 5467 4238
rect 5433 4204 5467 4236
rect 5433 4134 5467 4166
rect 5433 4132 5467 4134
rect 5691 4236 5725 4238
rect 5691 4204 5725 4236
rect 5691 4134 5725 4166
rect 5691 4132 5725 4134
rect 5949 4236 5983 4238
rect 5949 4204 5983 4236
rect 5949 4134 5983 4166
rect 5949 4132 5983 4134
rect 6132 4275 6166 4299
rect 6132 4231 6166 4237
rect 6132 4203 6166 4231
rect 6132 4163 6166 4165
rect 6132 4131 6166 4163
rect 340 4059 374 4061
rect 6132 4061 6166 4093
rect 6132 4059 6166 4061
rect 340 3993 374 4021
rect 623 4004 625 4038
rect 625 4004 657 4038
rect 695 4004 727 4038
rect 727 4004 729 4038
rect 881 4004 883 4038
rect 883 4004 915 4038
rect 953 4004 985 4038
rect 985 4004 987 4038
rect 5526 4004 5528 4038
rect 5528 4004 5560 4038
rect 5598 4004 5630 4038
rect 5630 4004 5632 4038
rect 5784 4004 5786 4038
rect 5786 4004 5818 4038
rect 5856 4004 5888 4038
rect 5888 4004 5890 4038
rect 340 3987 374 3993
rect 340 3925 374 3949
rect 340 3915 374 3925
rect 340 3857 374 3877
rect 340 3843 374 3857
rect 340 3789 374 3805
rect 340 3771 374 3789
rect 6132 3993 6166 4021
rect 6132 3987 6166 3993
rect 6132 3925 6166 3949
rect 6132 3915 6166 3925
rect 6132 3857 6166 3877
rect 6132 3843 6166 3857
rect 6132 3789 6166 3805
rect 6132 3771 6166 3789
rect 340 3721 374 3733
rect 623 3723 625 3757
rect 625 3723 657 3757
rect 695 3723 727 3757
rect 727 3723 729 3757
rect 881 3723 883 3757
rect 883 3723 915 3757
rect 953 3723 985 3757
rect 985 3723 987 3757
rect 5526 3723 5528 3757
rect 5528 3723 5560 3757
rect 5598 3723 5630 3757
rect 5630 3723 5632 3757
rect 5784 3723 5786 3757
rect 5786 3723 5818 3757
rect 5856 3723 5888 3757
rect 5888 3723 5890 3757
rect 340 3699 374 3721
rect 6132 3721 6166 3733
rect 6132 3699 6166 3721
rect 340 3653 374 3661
rect 340 3627 374 3653
rect 340 3585 374 3589
rect 340 3555 374 3585
rect 340 3483 374 3517
rect 530 3627 564 3629
rect 530 3595 564 3627
rect 530 3525 564 3557
rect 530 3523 564 3525
rect 788 3627 822 3629
rect 788 3595 822 3627
rect 788 3525 822 3557
rect 788 3523 822 3525
rect 1046 3627 1080 3629
rect 1046 3595 1080 3627
rect 1046 3525 1080 3557
rect 1046 3523 1080 3525
rect 5433 3627 5467 3629
rect 5433 3595 5467 3627
rect 5433 3525 5467 3557
rect 5433 3523 5467 3525
rect 5691 3627 5725 3629
rect 5691 3595 5725 3627
rect 5691 3525 5725 3557
rect 5691 3523 5725 3525
rect 5949 3627 5983 3629
rect 5949 3595 5983 3627
rect 5949 3525 5983 3557
rect 5949 3523 5983 3525
rect 6132 3653 6166 3661
rect 6132 3627 6166 3653
rect 6132 3585 6166 3589
rect 6132 3555 6166 3585
rect 6132 3483 6166 3517
rect 340 3415 374 3445
rect 340 3411 374 3415
rect 340 3347 374 3373
rect 340 3339 374 3347
rect 340 3279 374 3301
rect 340 3267 374 3279
rect 340 3211 374 3229
rect 340 3195 374 3211
rect 340 3143 374 3157
rect 340 3123 374 3143
rect 340 3075 374 3085
rect 340 3051 374 3075
rect 340 3007 374 3013
rect 340 2979 374 3007
rect 340 2939 374 2941
rect 340 2907 374 2939
rect 340 2837 374 2869
rect 340 2835 374 2837
rect 340 2769 374 2797
rect 6132 3415 6166 3445
rect 6132 3411 6166 3415
rect 6132 3347 6166 3373
rect 6132 3339 6166 3347
rect 6132 3279 6166 3301
rect 6132 3267 6166 3279
rect 6132 3211 6166 3229
rect 6132 3195 6166 3211
rect 6132 3143 6166 3157
rect 6132 3123 6166 3143
rect 6132 3075 6166 3085
rect 6132 3051 6166 3075
rect 6132 3007 6166 3013
rect 6132 2979 6166 3007
rect 6132 2939 6166 2941
rect 6132 2907 6166 2939
rect 6132 2837 6166 2869
rect 6132 2835 6166 2837
rect 340 2763 374 2769
rect 340 2701 374 2725
rect 340 2691 374 2701
rect 340 2633 374 2653
rect 340 2619 374 2633
rect 340 2565 374 2581
rect 530 2729 564 2731
rect 530 2697 564 2729
rect 530 2627 564 2659
rect 530 2625 564 2627
rect 788 2729 822 2731
rect 788 2697 822 2729
rect 788 2627 822 2659
rect 788 2625 822 2627
rect 1046 2729 1080 2731
rect 1046 2697 1080 2729
rect 1046 2627 1080 2659
rect 1046 2625 1080 2627
rect 5433 2729 5467 2731
rect 5433 2697 5467 2729
rect 5433 2627 5467 2659
rect 5433 2625 5467 2627
rect 5691 2729 5725 2731
rect 5691 2697 5725 2729
rect 5691 2627 5725 2659
rect 5691 2625 5725 2627
rect 5949 2729 5983 2731
rect 5949 2697 5983 2729
rect 5949 2627 5983 2659
rect 5949 2625 5983 2627
rect 6132 2769 6166 2797
rect 6132 2763 6166 2769
rect 6132 2701 6166 2725
rect 6132 2691 6166 2701
rect 6132 2633 6166 2653
rect 6132 2619 6166 2633
rect 340 2547 374 2565
rect 6132 2565 6166 2581
rect 6132 2547 6166 2565
rect 340 2497 374 2509
rect 623 2497 625 2531
rect 625 2497 657 2531
rect 695 2497 727 2531
rect 727 2497 729 2531
rect 881 2497 883 2531
rect 883 2497 915 2531
rect 953 2497 985 2531
rect 985 2497 987 2531
rect 5526 2497 5528 2531
rect 5528 2497 5560 2531
rect 5598 2497 5630 2531
rect 5630 2497 5632 2531
rect 5784 2497 5786 2531
rect 5786 2497 5818 2531
rect 5856 2497 5888 2531
rect 5888 2497 5890 2531
rect 6132 2497 6166 2509
rect 340 2475 374 2497
rect 340 2429 374 2437
rect 340 2403 374 2429
rect 340 2361 374 2365
rect 340 2331 374 2361
rect 340 2259 374 2293
rect 6132 2475 6166 2497
rect 6132 2429 6166 2437
rect 6132 2403 6166 2429
rect 6132 2361 6166 2365
rect 6132 2331 6166 2361
rect 6132 2259 6166 2293
rect 340 2191 374 2221
rect 623 2216 625 2250
rect 625 2216 657 2250
rect 695 2216 727 2250
rect 727 2216 729 2250
rect 881 2216 883 2250
rect 883 2216 915 2250
rect 953 2216 985 2250
rect 985 2216 987 2250
rect 5526 2216 5528 2250
rect 5528 2216 5560 2250
rect 5598 2216 5630 2250
rect 5630 2216 5632 2250
rect 5784 2216 5786 2250
rect 5786 2216 5818 2250
rect 5856 2216 5888 2250
rect 5888 2216 5890 2250
rect 340 2187 374 2191
rect 6132 2191 6166 2221
rect 6132 2187 6166 2191
rect 340 2123 374 2149
rect 340 2115 374 2123
rect 340 2043 374 2077
rect 530 2120 564 2122
rect 530 2088 564 2120
rect 530 2018 564 2050
rect 530 2016 564 2018
rect 788 2120 822 2122
rect 788 2088 822 2120
rect 788 2018 822 2050
rect 788 2016 822 2018
rect 1046 2120 1080 2122
rect 1046 2088 1080 2120
rect 1046 2018 1080 2050
rect 1046 2016 1080 2018
rect 5433 2120 5467 2122
rect 5433 2088 5467 2120
rect 5433 2018 5467 2050
rect 5433 2016 5467 2018
rect 5691 2120 5725 2122
rect 5691 2088 5725 2120
rect 5691 2018 5725 2050
rect 5691 2016 5725 2018
rect 5949 2120 5983 2122
rect 5949 2088 5983 2120
rect 5949 2018 5983 2050
rect 5949 2016 5983 2018
rect 6132 2123 6166 2149
rect 6132 2115 6166 2123
rect 6132 2043 6166 2077
rect 340 1894 374 1928
rect 340 1848 374 1856
rect 340 1822 374 1848
rect 340 1780 374 1784
rect 340 1750 374 1780
rect 340 1678 374 1712
rect 340 1610 374 1640
rect 340 1606 374 1610
rect 6132 1894 6166 1928
rect 6132 1848 6166 1856
rect 6132 1822 6166 1848
rect 6132 1780 6166 1784
rect 6132 1750 6166 1780
rect 6132 1678 6166 1712
rect 6132 1610 6166 1640
rect 6132 1606 6166 1610
rect 340 1542 374 1568
rect 340 1534 374 1542
rect 6132 1542 6166 1568
rect 340 1474 374 1496
rect 340 1462 374 1474
rect 340 1406 374 1424
rect 6132 1534 6166 1542
rect 6132 1474 6166 1496
rect 6132 1462 6166 1474
rect 340 1390 374 1406
rect 340 1338 374 1352
rect 340 1318 374 1338
rect 340 1270 374 1280
rect 340 1246 374 1270
rect 340 1202 374 1208
rect 530 1360 564 1362
rect 530 1328 564 1360
rect 530 1258 564 1290
rect 530 1256 564 1258
rect 788 1360 822 1362
rect 788 1328 822 1360
rect 788 1258 822 1290
rect 788 1256 822 1258
rect 1046 1360 1080 1362
rect 1046 1328 1080 1360
rect 1046 1258 1080 1290
rect 1046 1256 1080 1258
rect 5433 1360 5467 1362
rect 5433 1328 5467 1360
rect 5433 1258 5467 1290
rect 5433 1256 5467 1258
rect 5691 1360 5725 1362
rect 5691 1328 5725 1360
rect 5691 1258 5725 1290
rect 5691 1256 5725 1258
rect 5949 1360 5983 1362
rect 5949 1328 5983 1360
rect 5949 1258 5983 1290
rect 5949 1256 5983 1258
rect 6132 1406 6166 1424
rect 6132 1390 6166 1406
rect 6132 1338 6166 1352
rect 6132 1318 6166 1338
rect 6132 1270 6166 1280
rect 6132 1246 6166 1270
rect 340 1174 374 1202
rect 6132 1202 6166 1208
rect 6132 1174 6166 1202
rect 340 1134 374 1136
rect 340 1102 374 1134
rect 623 1128 625 1162
rect 625 1128 657 1162
rect 695 1128 727 1162
rect 727 1128 729 1162
rect 881 1128 883 1162
rect 883 1128 915 1162
rect 953 1128 985 1162
rect 985 1128 987 1162
rect 5526 1128 5528 1162
rect 5528 1128 5560 1162
rect 5598 1128 5630 1162
rect 5630 1128 5632 1162
rect 5784 1128 5786 1162
rect 5786 1128 5818 1162
rect 5856 1128 5888 1162
rect 5888 1128 5890 1162
rect 6132 1134 6166 1136
rect 340 1032 374 1064
rect 340 1030 374 1032
rect 340 964 374 992
rect 340 958 374 964
rect 340 896 374 920
rect 340 886 374 896
rect 6132 1102 6166 1134
rect 6132 1032 6166 1064
rect 6132 1030 6166 1032
rect 6132 964 6166 992
rect 6132 958 6166 964
rect 6132 896 6166 920
rect 6132 886 6166 896
rect 340 828 374 848
rect 623 847 625 881
rect 625 847 657 881
rect 695 847 727 881
rect 727 847 729 881
rect 881 847 883 881
rect 883 847 915 881
rect 953 847 985 881
rect 985 847 987 881
rect 5526 847 5528 881
rect 5528 847 5560 881
rect 5598 847 5630 881
rect 5630 847 5632 881
rect 5784 847 5786 881
rect 5786 847 5818 881
rect 5856 847 5888 881
rect 5888 847 5890 881
rect 340 814 374 828
rect 6132 828 6166 848
rect 6132 814 6166 828
rect 340 760 374 776
rect 340 742 374 760
rect 340 692 374 704
rect 340 670 374 692
rect 340 624 374 632
rect 340 598 374 624
rect 530 751 564 753
rect 530 719 564 751
rect 530 649 564 681
rect 530 647 564 649
rect 788 751 822 753
rect 788 719 822 751
rect 788 649 822 681
rect 788 647 822 649
rect 1046 751 1080 753
rect 1046 719 1080 751
rect 1046 649 1080 681
rect 1046 647 1080 649
rect 5433 751 5467 753
rect 5433 719 5467 751
rect 5433 649 5467 681
rect 5433 647 5467 649
rect 5691 751 5725 753
rect 5691 719 5725 751
rect 5691 649 5725 681
rect 5691 647 5725 649
rect 5949 751 5983 753
rect 5949 719 5983 751
rect 5949 649 5983 681
rect 5949 647 5983 649
rect 6132 760 6166 776
rect 6132 742 6166 760
rect 6132 692 6166 704
rect 6132 670 6166 692
rect 6132 624 6166 632
rect 6132 598 6166 624
rect 340 556 374 560
rect 340 526 374 556
rect 340 454 374 488
rect 340 386 374 416
rect 340 382 374 386
rect 340 318 374 344
rect 6132 556 6166 560
rect 6132 526 6166 556
rect 6132 454 6166 488
rect 6132 386 6166 416
rect 6132 382 6166 386
rect 6132 318 6166 344
rect 340 310 374 318
rect 340 250 374 272
rect 340 238 374 250
rect 340 182 374 200
rect 340 166 374 182
rect 340 114 374 128
rect 340 94 374 114
rect 530 265 564 267
rect 530 233 564 265
rect 530 163 564 195
rect 530 161 564 163
rect 788 265 822 267
rect 788 233 822 265
rect 788 163 822 195
rect 788 161 822 163
rect 1046 265 1080 267
rect 1046 233 1080 265
rect 1046 163 1080 195
rect 1046 161 1080 163
rect 5433 265 5467 267
rect 5433 233 5467 265
rect 5433 163 5467 195
rect 5433 161 5467 163
rect 5691 265 5725 267
rect 5691 233 5725 265
rect 5691 163 5725 195
rect 5691 161 5725 163
rect 5949 265 5983 267
rect 5949 233 5983 265
rect 5949 163 5983 195
rect 5949 161 5983 163
rect 6132 310 6166 318
rect 6132 250 6166 272
rect 6132 238 6166 250
rect 6132 182 6166 200
rect 6132 166 6166 182
rect 6132 114 6166 128
rect 6132 94 6166 114
rect 340 46 374 56
rect 340 22 374 46
rect 623 33 625 67
rect 625 33 657 67
rect 695 33 727 67
rect 727 33 729 67
rect 881 33 883 67
rect 883 33 915 67
rect 953 33 985 67
rect 985 33 987 67
rect 5526 33 5528 67
rect 5528 33 5560 67
rect 5598 33 5630 67
rect 5630 33 5632 67
rect 5784 33 5786 67
rect 5786 33 5818 67
rect 5856 33 5888 67
rect 5888 33 5890 67
rect 6132 46 6166 56
rect 340 -22 374 -16
rect 340 -50 374 -22
rect 340 -90 374 -88
rect 340 -122 374 -90
rect 340 -192 374 -160
rect 340 -194 374 -192
rect 6132 22 6166 46
rect 6132 -22 6166 -16
rect 6132 -50 6166 -22
rect 6132 -90 6166 -88
rect 6132 -122 6166 -90
rect 6132 -192 6166 -160
rect 6132 -194 6166 -192
rect 340 -260 374 -232
rect 623 -248 625 -214
rect 625 -248 657 -214
rect 695 -248 727 -214
rect 727 -248 729 -214
rect 881 -248 883 -214
rect 883 -248 915 -214
rect 953 -248 985 -214
rect 985 -248 987 -214
rect 5526 -248 5528 -214
rect 5528 -248 5560 -214
rect 5598 -248 5630 -214
rect 5630 -248 5632 -214
rect 5784 -248 5786 -214
rect 5786 -248 5818 -214
rect 5856 -248 5888 -214
rect 5888 -248 5890 -214
rect 340 -266 374 -260
rect 6132 -260 6166 -232
rect 6132 -266 6166 -260
rect 340 -328 374 -304
rect 340 -338 374 -328
rect 340 -396 374 -376
rect 340 -410 374 -396
rect 340 -464 374 -448
rect 340 -482 374 -464
rect 530 -344 564 -342
rect 530 -376 564 -344
rect 530 -446 564 -414
rect 530 -448 564 -446
rect 788 -344 822 -342
rect 788 -376 822 -344
rect 788 -446 822 -414
rect 788 -448 822 -446
rect 1046 -344 1080 -342
rect 1046 -376 1080 -344
rect 1046 -446 1080 -414
rect 1046 -448 1080 -446
rect 5433 -344 5467 -342
rect 5433 -376 5467 -344
rect 5433 -446 5467 -414
rect 5433 -448 5467 -446
rect 5691 -344 5725 -342
rect 5691 -376 5725 -344
rect 5691 -446 5725 -414
rect 5691 -448 5725 -446
rect 5949 -344 5983 -342
rect 5949 -376 5983 -344
rect 5949 -446 5983 -414
rect 5949 -448 5983 -446
rect 6132 -328 6166 -304
rect 6132 -338 6166 -328
rect 6132 -396 6166 -376
rect 6132 -410 6166 -396
rect 6132 -464 6166 -448
rect 6132 -482 6166 -464
rect 340 -532 374 -520
rect 340 -554 374 -532
rect 340 -600 374 -592
rect 340 -626 374 -600
rect 340 -668 374 -664
rect 340 -698 374 -668
rect 340 -770 374 -736
rect 6132 -532 6166 -520
rect 6132 -554 6166 -532
rect 6132 -600 6166 -592
rect 6132 -626 6166 -600
rect 6132 -668 6166 -664
rect 6132 -698 6166 -668
rect 340 -838 374 -808
rect 340 -842 374 -838
rect 340 -906 374 -880
rect 340 -914 374 -906
rect 340 -974 374 -952
rect 340 -986 374 -974
rect 530 -821 564 -819
rect 530 -853 564 -821
rect 530 -923 564 -891
rect 530 -925 564 -923
rect 788 -821 822 -819
rect 788 -853 822 -821
rect 788 -923 822 -891
rect 788 -925 822 -923
rect 1046 -821 1080 -819
rect 1046 -853 1080 -821
rect 1046 -923 1080 -891
rect 1046 -925 1080 -923
rect 5433 -821 5467 -819
rect 5433 -853 5467 -821
rect 5433 -923 5467 -891
rect 5433 -925 5467 -923
rect 5691 -821 5725 -819
rect 5691 -853 5725 -821
rect 5691 -923 5725 -891
rect 5691 -925 5725 -923
rect 5949 -821 5983 -819
rect 5949 -853 5983 -821
rect 5949 -923 5983 -891
rect 5949 -925 5983 -923
rect 6132 -770 6166 -736
rect 6132 -838 6166 -808
rect 6132 -842 6166 -838
rect 6132 -906 6166 -880
rect 6132 -914 6166 -906
rect 6132 -974 6166 -952
rect 6132 -986 6166 -974
rect 340 -1042 374 -1024
rect 340 -1058 374 -1042
rect 623 -1053 625 -1019
rect 625 -1053 657 -1019
rect 695 -1053 727 -1019
rect 727 -1053 729 -1019
rect 881 -1053 883 -1019
rect 883 -1053 915 -1019
rect 953 -1053 985 -1019
rect 985 -1053 987 -1019
rect 5526 -1053 5528 -1019
rect 5528 -1053 5560 -1019
rect 5598 -1053 5630 -1019
rect 5630 -1053 5632 -1019
rect 5784 -1053 5786 -1019
rect 5786 -1053 5818 -1019
rect 5856 -1053 5888 -1019
rect 5888 -1053 5890 -1019
rect 6132 -1042 6166 -1024
rect 340 -1110 374 -1096
rect 340 -1130 374 -1110
rect 6132 -1058 6166 -1042
rect 6132 -1110 6166 -1096
rect 6132 -1130 6166 -1110
rect 340 -1178 374 -1168
rect 340 -1202 374 -1178
rect 6132 -1178 6166 -1168
rect 340 -1246 374 -1240
rect 340 -1274 374 -1246
rect 6132 -1202 6166 -1178
rect 6132 -1246 6166 -1240
rect 6132 -1274 6166 -1246
rect 340 -1314 374 -1312
rect 340 -1346 374 -1314
rect 623 -1334 625 -1300
rect 625 -1334 657 -1300
rect 695 -1334 727 -1300
rect 727 -1334 729 -1300
rect 881 -1334 883 -1300
rect 883 -1334 915 -1300
rect 953 -1334 985 -1300
rect 985 -1334 987 -1300
rect 5526 -1334 5528 -1300
rect 5528 -1334 5560 -1300
rect 5598 -1334 5630 -1300
rect 5630 -1334 5632 -1300
rect 5784 -1334 5786 -1300
rect 5786 -1334 5818 -1300
rect 5856 -1334 5888 -1300
rect 5888 -1334 5890 -1300
rect 6132 -1314 6166 -1312
rect 6132 -1346 6166 -1314
rect 340 -1416 374 -1384
rect 340 -1418 374 -1416
rect 340 -1484 374 -1456
rect 340 -1490 374 -1484
rect 340 -1552 374 -1528
rect 340 -1562 374 -1552
rect 530 -1430 564 -1428
rect 530 -1462 564 -1430
rect 530 -1532 564 -1500
rect 530 -1534 564 -1532
rect 788 -1430 822 -1428
rect 788 -1462 822 -1430
rect 788 -1532 822 -1500
rect 788 -1534 822 -1532
rect 1046 -1430 1080 -1428
rect 1046 -1462 1080 -1430
rect 1046 -1532 1080 -1500
rect 1046 -1534 1080 -1532
rect 5433 -1430 5467 -1428
rect 5433 -1462 5467 -1430
rect 5433 -1532 5467 -1500
rect 5433 -1534 5467 -1532
rect 5691 -1430 5725 -1428
rect 5691 -1462 5725 -1430
rect 5691 -1532 5725 -1500
rect 5691 -1534 5725 -1532
rect 5949 -1430 5983 -1428
rect 5949 -1462 5983 -1430
rect 5949 -1532 5983 -1500
rect 5949 -1534 5983 -1532
rect 6132 -1416 6166 -1384
rect 6132 -1418 6166 -1416
rect 6132 -1484 6166 -1456
rect 6132 -1490 6166 -1484
rect 6132 -1552 6166 -1528
rect 6132 -1562 6166 -1552
rect 340 -1620 374 -1600
rect 340 -1634 374 -1620
rect 340 -1688 374 -1672
rect 340 -1706 374 -1688
rect 340 -1756 374 -1744
rect 340 -1778 374 -1756
rect 340 -1824 374 -1816
rect 340 -1850 374 -1824
rect 340 -1892 374 -1888
rect 340 -1922 374 -1892
rect 340 -1994 374 -1960
rect 340 -2062 374 -2032
rect 340 -2066 374 -2062
rect 340 -2130 374 -2104
rect 340 -2138 374 -2130
rect 340 -2198 374 -2176
rect 340 -2210 374 -2198
rect 340 -2266 374 -2248
rect 340 -2282 374 -2266
rect 6132 -1620 6166 -1600
rect 6132 -1634 6166 -1620
rect 6132 -1688 6166 -1672
rect 6132 -1706 6166 -1688
rect 6132 -1756 6166 -1744
rect 6132 -1778 6166 -1756
rect 6132 -1824 6166 -1816
rect 6132 -1850 6166 -1824
rect 6132 -1892 6166 -1888
rect 6132 -1922 6166 -1892
rect 6132 -1994 6166 -1960
rect 6132 -2062 6166 -2032
rect 6132 -2066 6166 -2062
rect 6132 -2130 6166 -2104
rect 6132 -2138 6166 -2130
rect 6132 -2198 6166 -2176
rect 6132 -2210 6166 -2198
rect 6132 -2266 6166 -2248
rect 340 -2334 374 -2320
rect 340 -2354 374 -2334
rect 340 -2402 374 -2392
rect 340 -2426 374 -2402
rect 340 -2470 374 -2464
rect 340 -2498 374 -2470
rect 530 -2325 564 -2323
rect 530 -2357 564 -2325
rect 530 -2427 564 -2395
rect 530 -2429 564 -2427
rect 788 -2325 822 -2323
rect 788 -2357 822 -2325
rect 788 -2427 822 -2395
rect 788 -2429 822 -2427
rect 1046 -2325 1080 -2323
rect 1046 -2357 1080 -2325
rect 1046 -2427 1080 -2395
rect 1046 -2429 1080 -2427
rect 5433 -2325 5467 -2323
rect 5433 -2357 5467 -2325
rect 5433 -2427 5467 -2395
rect 5433 -2429 5467 -2427
rect 5691 -2325 5725 -2323
rect 5691 -2357 5725 -2325
rect 5691 -2427 5725 -2395
rect 5691 -2429 5725 -2427
rect 5949 -2325 5983 -2323
rect 5949 -2357 5983 -2325
rect 5949 -2427 5983 -2395
rect 5949 -2429 5983 -2427
rect 6132 -2282 6166 -2266
rect 6132 -2334 6166 -2320
rect 6132 -2354 6166 -2334
rect 6132 -2402 6166 -2392
rect 6132 -2426 6166 -2402
rect 6132 -2470 6166 -2464
rect 6132 -2498 6166 -2470
rect 340 -2538 374 -2536
rect 340 -2570 374 -2538
rect 623 -2557 625 -2523
rect 625 -2557 657 -2523
rect 695 -2557 727 -2523
rect 727 -2557 729 -2523
rect 881 -2557 883 -2523
rect 883 -2557 915 -2523
rect 953 -2557 985 -2523
rect 985 -2557 987 -2523
rect 5526 -2557 5528 -2523
rect 5528 -2557 5560 -2523
rect 5598 -2557 5630 -2523
rect 5630 -2557 5632 -2523
rect 5784 -2557 5786 -2523
rect 5786 -2557 5818 -2523
rect 5856 -2557 5888 -2523
rect 5888 -2557 5890 -2523
rect 6132 -2538 6166 -2536
rect 340 -2640 374 -2608
rect 340 -2642 374 -2640
rect 340 -2708 374 -2680
rect 340 -2714 374 -2708
rect 340 -2776 374 -2752
rect 340 -2786 374 -2776
rect 6132 -2570 6166 -2538
rect 6132 -2640 6166 -2608
rect 6132 -2642 6166 -2640
rect 6132 -2708 6166 -2680
rect 6132 -2714 6166 -2708
rect 6132 -2776 6166 -2752
rect 6132 -2786 6166 -2776
rect 340 -2844 374 -2824
rect 623 -2838 625 -2804
rect 625 -2838 657 -2804
rect 695 -2838 727 -2804
rect 727 -2838 729 -2804
rect 881 -2838 883 -2804
rect 883 -2838 915 -2804
rect 953 -2838 985 -2804
rect 985 -2838 987 -2804
rect 5526 -2838 5528 -2804
rect 5528 -2838 5560 -2804
rect 5598 -2838 5630 -2804
rect 5630 -2838 5632 -2804
rect 5784 -2838 5786 -2804
rect 5786 -2838 5818 -2804
rect 5856 -2838 5888 -2804
rect 5888 -2838 5890 -2804
rect 340 -2858 374 -2844
rect 6132 -2844 6166 -2824
rect 6132 -2858 6166 -2844
rect 340 -2912 374 -2896
rect 340 -2930 374 -2912
rect 340 -2980 374 -2968
rect 340 -3002 374 -2980
rect 340 -3048 374 -3040
rect 340 -3074 374 -3048
rect 530 -2934 564 -2932
rect 530 -2966 564 -2934
rect 530 -3036 564 -3004
rect 530 -3038 564 -3036
rect 788 -2934 822 -2932
rect 788 -2966 822 -2934
rect 788 -3036 822 -3004
rect 788 -3038 822 -3036
rect 1046 -2934 1080 -2932
rect 1046 -2966 1080 -2934
rect 1046 -3036 1080 -3004
rect 1046 -3038 1080 -3036
rect 5433 -2934 5467 -2932
rect 5433 -2966 5467 -2934
rect 5433 -3036 5467 -3004
rect 5433 -3038 5467 -3036
rect 5691 -2934 5725 -2932
rect 5691 -2966 5725 -2934
rect 5691 -3036 5725 -3004
rect 5691 -3038 5725 -3036
rect 5949 -2934 5983 -2932
rect 5949 -2966 5983 -2934
rect 5949 -3036 5983 -3004
rect 5949 -3038 5983 -3036
rect 6132 -2912 6166 -2896
rect 6132 -2930 6166 -2912
rect 6132 -2980 6166 -2968
rect 6132 -3002 6166 -2980
rect 6132 -3048 6166 -3040
rect 6132 -3074 6166 -3048
rect 340 -3116 374 -3112
rect 340 -3146 374 -3116
rect 340 -3218 374 -3184
rect 340 -3286 374 -3256
rect 340 -3290 374 -3286
rect 340 -3354 374 -3328
rect 340 -3362 374 -3354
rect 340 -3422 374 -3400
rect 340 -3434 374 -3422
rect 340 -3490 374 -3472
rect 340 -3506 374 -3490
rect 340 -3558 374 -3544
rect 340 -3578 374 -3558
rect 340 -3626 374 -3616
rect 340 -3650 374 -3626
rect 340 -3694 374 -3688
rect 340 -3722 374 -3694
rect 340 -3762 374 -3760
rect 340 -3794 374 -3762
rect 6132 -3116 6166 -3112
rect 6132 -3146 6166 -3116
rect 6132 -3218 6166 -3184
rect 6132 -3286 6166 -3256
rect 6132 -3290 6166 -3286
rect 6132 -3354 6166 -3328
rect 6132 -3362 6166 -3354
rect 6132 -3422 6166 -3400
rect 6132 -3434 6166 -3422
rect 6132 -3490 6166 -3472
rect 6132 -3506 6166 -3490
rect 6132 -3558 6166 -3544
rect 6132 -3578 6166 -3558
rect 6132 -3626 6166 -3616
rect 6132 -3650 6166 -3626
rect 6132 -3694 6166 -3688
rect 6132 -3722 6166 -3694
rect 6132 -3762 6166 -3760
rect 340 -3864 374 -3832
rect 340 -3866 374 -3864
rect 340 -3932 374 -3904
rect 340 -3938 374 -3932
rect 340 -4000 374 -3976
rect 530 -3829 564 -3827
rect 530 -3861 564 -3829
rect 530 -3931 564 -3899
rect 530 -3933 564 -3931
rect 788 -3829 822 -3827
rect 788 -3861 822 -3829
rect 788 -3931 822 -3899
rect 788 -3933 822 -3931
rect 1046 -3829 1080 -3827
rect 1046 -3861 1080 -3829
rect 1046 -3931 1080 -3899
rect 1046 -3933 1080 -3931
rect 5433 -3829 5467 -3827
rect 5433 -3861 5467 -3829
rect 5433 -3931 5467 -3899
rect 5433 -3933 5467 -3931
rect 5691 -3829 5725 -3827
rect 5691 -3861 5725 -3829
rect 5691 -3931 5725 -3899
rect 5691 -3933 5725 -3931
rect 5949 -3829 5983 -3827
rect 5949 -3861 5983 -3829
rect 5949 -3931 5983 -3899
rect 5949 -3933 5983 -3931
rect 6132 -3794 6166 -3762
rect 6132 -3864 6166 -3832
rect 6132 -3866 6166 -3864
rect 6132 -3932 6166 -3904
rect 6132 -3938 6166 -3932
rect 340 -4010 374 -4000
rect 6132 -4000 6166 -3976
rect 6132 -4010 6166 -4000
rect 340 -4068 374 -4048
rect 623 -4061 625 -4027
rect 625 -4061 657 -4027
rect 695 -4061 727 -4027
rect 727 -4061 729 -4027
rect 881 -4061 883 -4027
rect 883 -4061 915 -4027
rect 953 -4061 985 -4027
rect 985 -4061 987 -4027
rect 5526 -4061 5528 -4027
rect 5528 -4061 5560 -4027
rect 5598 -4061 5630 -4027
rect 5630 -4061 5632 -4027
rect 5784 -4061 5786 -4027
rect 5786 -4061 5818 -4027
rect 5856 -4061 5888 -4027
rect 5888 -4061 5890 -4027
rect 340 -4082 374 -4068
rect 340 -4136 374 -4120
rect 340 -4154 374 -4136
rect 340 -4204 374 -4192
rect 340 -4226 374 -4204
rect 340 -4272 374 -4264
rect 340 -4298 374 -4272
rect 6132 -4068 6166 -4048
rect 6132 -4082 6166 -4068
rect 6132 -4136 6166 -4120
rect 6132 -4154 6166 -4136
rect 6132 -4204 6166 -4192
rect 6132 -4226 6166 -4204
rect 6132 -4272 6166 -4264
rect 6132 -4298 6166 -4272
rect 340 -4340 374 -4336
rect 340 -4370 374 -4340
rect 623 -4342 625 -4308
rect 625 -4342 657 -4308
rect 695 -4342 727 -4308
rect 727 -4342 729 -4308
rect 881 -4342 883 -4308
rect 883 -4342 915 -4308
rect 953 -4342 985 -4308
rect 985 -4342 987 -4308
rect 5526 -4342 5528 -4308
rect 5528 -4342 5560 -4308
rect 5598 -4342 5630 -4308
rect 5630 -4342 5632 -4308
rect 5784 -4342 5786 -4308
rect 5786 -4342 5818 -4308
rect 5856 -4342 5888 -4308
rect 5888 -4342 5890 -4308
rect 6132 -4340 6166 -4336
rect 6132 -4370 6166 -4340
rect 340 -4442 374 -4408
rect 340 -4510 374 -4480
rect 340 -4514 374 -4510
rect 340 -4578 374 -4552
rect 340 -4586 374 -4578
rect 530 -4438 564 -4436
rect 530 -4470 564 -4438
rect 530 -4540 564 -4508
rect 530 -4542 564 -4540
rect 788 -4438 822 -4436
rect 788 -4470 822 -4438
rect 788 -4540 822 -4508
rect 788 -4542 822 -4540
rect 1046 -4438 1080 -4436
rect 1046 -4470 1080 -4438
rect 1046 -4540 1080 -4508
rect 1046 -4542 1080 -4540
rect 5433 -4438 5467 -4436
rect 5433 -4470 5467 -4438
rect 5433 -4540 5467 -4508
rect 5433 -4542 5467 -4540
rect 5691 -4438 5725 -4436
rect 5691 -4470 5725 -4438
rect 5691 -4540 5725 -4508
rect 5691 -4542 5725 -4540
rect 5949 -4438 5983 -4436
rect 5949 -4470 5983 -4438
rect 5949 -4540 5983 -4508
rect 5949 -4542 5983 -4540
rect 6132 -4442 6166 -4408
rect 6132 -4510 6166 -4480
rect 6132 -4514 6166 -4510
rect 6132 -4578 6166 -4552
rect 6132 -4586 6166 -4578
rect 340 -4646 374 -4624
rect 340 -4658 374 -4646
rect 340 -4714 374 -4696
rect 340 -4730 374 -4714
rect 340 -4782 374 -4768
rect 340 -4802 374 -4782
rect 340 -4850 374 -4840
rect 340 -4874 374 -4850
rect 340 -4918 374 -4912
rect 340 -4946 374 -4918
rect 340 -4986 374 -4984
rect 340 -5018 374 -4986
rect 340 -5088 374 -5056
rect 340 -5090 374 -5088
rect 340 -5156 374 -5128
rect 6132 -4646 6166 -4624
rect 6132 -4658 6166 -4646
rect 6132 -4714 6166 -4696
rect 6132 -4730 6166 -4714
rect 6132 -4782 6166 -4768
rect 6132 -4802 6166 -4782
rect 6132 -4850 6166 -4840
rect 6132 -4874 6166 -4850
rect 6132 -4918 6166 -4912
rect 6132 -4946 6166 -4918
rect 6132 -4986 6166 -4984
rect 6132 -5018 6166 -4986
rect 6132 -5088 6166 -5056
rect 6132 -5090 6166 -5088
rect 340 -5162 374 -5156
rect 340 -5224 374 -5200
rect 340 -5234 374 -5224
rect 340 -5292 374 -5272
rect 340 -5306 374 -5292
rect 530 -5185 564 -5183
rect 530 -5217 564 -5185
rect 530 -5287 564 -5255
rect 530 -5289 564 -5287
rect 788 -5185 822 -5183
rect 788 -5217 822 -5185
rect 788 -5287 822 -5255
rect 788 -5289 822 -5287
rect 1046 -5185 1080 -5183
rect 1046 -5217 1080 -5185
rect 1046 -5287 1080 -5255
rect 1046 -5289 1080 -5287
rect 1240 -5185 1274 -5183
rect 1240 -5217 1274 -5185
rect 1240 -5287 1274 -5255
rect 1240 -5289 1274 -5287
rect 1498 -5185 1532 -5183
rect 1498 -5217 1532 -5185
rect 1498 -5287 1532 -5255
rect 1498 -5289 1532 -5287
rect 1756 -5185 1790 -5183
rect 1756 -5217 1790 -5185
rect 1756 -5287 1790 -5255
rect 1756 -5289 1790 -5287
rect 2014 -5185 2048 -5183
rect 2014 -5217 2048 -5185
rect 2014 -5287 2048 -5255
rect 2014 -5289 2048 -5287
rect 2272 -5185 2306 -5183
rect 2272 -5217 2306 -5185
rect 2272 -5287 2306 -5255
rect 2272 -5289 2306 -5287
rect 2466 -5185 2500 -5183
rect 2466 -5217 2500 -5185
rect 2466 -5287 2500 -5255
rect 2466 -5289 2500 -5287
rect 2724 -5185 2758 -5183
rect 2724 -5217 2758 -5185
rect 2724 -5287 2758 -5255
rect 2724 -5289 2758 -5287
rect 2982 -5185 3016 -5183
rect 2982 -5217 3016 -5185
rect 2982 -5287 3016 -5255
rect 2982 -5289 3016 -5287
rect 3240 -5185 3274 -5183
rect 3240 -5217 3274 -5185
rect 3240 -5287 3274 -5255
rect 3240 -5289 3274 -5287
rect 3498 -5185 3532 -5183
rect 3498 -5217 3532 -5185
rect 3498 -5287 3532 -5255
rect 3498 -5289 3532 -5287
rect 3756 -5185 3790 -5183
rect 3756 -5217 3790 -5185
rect 3756 -5287 3790 -5255
rect 3756 -5289 3790 -5287
rect 4014 -5185 4048 -5183
rect 4014 -5217 4048 -5185
rect 4014 -5287 4048 -5255
rect 4014 -5289 4048 -5287
rect 4208 -5185 4242 -5183
rect 4208 -5217 4242 -5185
rect 4208 -5287 4242 -5255
rect 4208 -5289 4242 -5287
rect 4466 -5185 4500 -5183
rect 4466 -5217 4500 -5185
rect 4466 -5287 4500 -5255
rect 4466 -5289 4500 -5287
rect 4724 -5185 4758 -5183
rect 4724 -5217 4758 -5185
rect 4724 -5287 4758 -5255
rect 4724 -5289 4758 -5287
rect 4982 -5185 5016 -5183
rect 4982 -5217 5016 -5185
rect 4982 -5287 5016 -5255
rect 4982 -5289 5016 -5287
rect 5240 -5185 5274 -5183
rect 5240 -5217 5274 -5185
rect 5240 -5287 5274 -5255
rect 5240 -5289 5274 -5287
rect 5433 -5185 5467 -5183
rect 5433 -5217 5467 -5185
rect 5433 -5287 5467 -5255
rect 5433 -5289 5467 -5287
rect 5691 -5185 5725 -5183
rect 5691 -5217 5725 -5185
rect 5691 -5287 5725 -5255
rect 5691 -5289 5725 -5287
rect 5949 -5185 5983 -5183
rect 5949 -5217 5983 -5185
rect 5949 -5287 5983 -5255
rect 5949 -5289 5983 -5287
rect 6132 -5156 6166 -5128
rect 6132 -5162 6166 -5156
rect 6132 -5224 6166 -5200
rect 6132 -5234 6166 -5224
rect 6132 -5292 6166 -5272
rect 6132 -5306 6166 -5292
rect 340 -5360 374 -5344
rect 340 -5378 374 -5360
rect 6132 -5360 6166 -5344
rect 6132 -5378 6166 -5360
rect 623 -5417 625 -5383
rect 625 -5417 657 -5383
rect 695 -5417 727 -5383
rect 727 -5417 729 -5383
rect 881 -5417 883 -5383
rect 883 -5417 915 -5383
rect 953 -5417 985 -5383
rect 985 -5417 987 -5383
rect 1333 -5417 1335 -5383
rect 1335 -5417 1367 -5383
rect 1405 -5417 1437 -5383
rect 1437 -5417 1439 -5383
rect 1591 -5417 1593 -5383
rect 1593 -5417 1625 -5383
rect 1663 -5417 1695 -5383
rect 1695 -5417 1697 -5383
rect 1849 -5417 1851 -5383
rect 1851 -5417 1883 -5383
rect 1921 -5417 1953 -5383
rect 1953 -5417 1955 -5383
rect 2107 -5417 2109 -5383
rect 2109 -5417 2141 -5383
rect 2179 -5417 2211 -5383
rect 2211 -5417 2213 -5383
rect 2559 -5417 2561 -5383
rect 2561 -5417 2593 -5383
rect 2631 -5417 2663 -5383
rect 2663 -5417 2665 -5383
rect 2817 -5417 2819 -5383
rect 2819 -5417 2851 -5383
rect 2889 -5417 2921 -5383
rect 2921 -5417 2923 -5383
rect 3075 -5417 3077 -5383
rect 3077 -5417 3109 -5383
rect 3147 -5417 3179 -5383
rect 3179 -5417 3181 -5383
rect 3333 -5417 3335 -5383
rect 3335 -5417 3367 -5383
rect 3405 -5417 3437 -5383
rect 3437 -5417 3439 -5383
rect 3591 -5417 3593 -5383
rect 3593 -5417 3625 -5383
rect 3663 -5417 3695 -5383
rect 3695 -5417 3697 -5383
rect 3849 -5417 3851 -5383
rect 3851 -5417 3883 -5383
rect 3921 -5417 3953 -5383
rect 3953 -5417 3955 -5383
rect 4301 -5417 4303 -5383
rect 4303 -5417 4335 -5383
rect 4373 -5417 4405 -5383
rect 4405 -5417 4407 -5383
rect 4559 -5417 4561 -5383
rect 4561 -5417 4593 -5383
rect 4631 -5417 4663 -5383
rect 4663 -5417 4665 -5383
rect 4817 -5417 4819 -5383
rect 4819 -5417 4851 -5383
rect 4889 -5417 4921 -5383
rect 4921 -5417 4923 -5383
rect 5075 -5417 5077 -5383
rect 5077 -5417 5109 -5383
rect 5147 -5417 5179 -5383
rect 5179 -5417 5181 -5383
rect 5526 -5417 5528 -5383
rect 5528 -5417 5560 -5383
rect 5598 -5417 5630 -5383
rect 5630 -5417 5632 -5383
rect 5784 -5417 5786 -5383
rect 5786 -5417 5818 -5383
rect 5856 -5417 5888 -5383
rect 5888 -5417 5890 -5383
rect 487 -5540 495 -5506
rect 495 -5540 521 -5506
rect 559 -5540 563 -5506
rect 563 -5540 593 -5506
rect 631 -5540 665 -5506
rect 703 -5540 733 -5506
rect 733 -5540 737 -5506
rect 775 -5540 801 -5506
rect 801 -5540 809 -5506
rect 847 -5540 869 -5506
rect 869 -5540 881 -5506
rect 919 -5540 937 -5506
rect 937 -5540 953 -5506
rect 991 -5540 1005 -5506
rect 1005 -5540 1025 -5506
rect 1063 -5540 1073 -5506
rect 1073 -5540 1097 -5506
rect 1135 -5540 1141 -5506
rect 1141 -5540 1169 -5506
rect 1207 -5540 1209 -5506
rect 1209 -5540 1241 -5506
rect 1279 -5540 1311 -5506
rect 1311 -5540 1313 -5506
rect 1351 -5540 1379 -5506
rect 1379 -5540 1385 -5506
rect 1423 -5540 1447 -5506
rect 1447 -5540 1457 -5506
rect 1495 -5540 1515 -5506
rect 1515 -5540 1529 -5506
rect 1567 -5540 1583 -5506
rect 1583 -5540 1601 -5506
rect 1639 -5540 1651 -5506
rect 1651 -5540 1673 -5506
rect 1711 -5540 1719 -5506
rect 1719 -5540 1745 -5506
rect 1783 -5540 1787 -5506
rect 1787 -5540 1817 -5506
rect 1855 -5540 1889 -5506
rect 1927 -5540 1957 -5506
rect 1957 -5540 1961 -5506
rect 1999 -5540 2025 -5506
rect 2025 -5540 2033 -5506
rect 2071 -5540 2093 -5506
rect 2093 -5540 2105 -5506
rect 2143 -5540 2161 -5506
rect 2161 -5540 2177 -5506
rect 2215 -5540 2229 -5506
rect 2229 -5540 2249 -5506
rect 2287 -5540 2297 -5506
rect 2297 -5540 2321 -5506
rect 2359 -5540 2365 -5506
rect 2365 -5540 2393 -5506
rect 2431 -5540 2433 -5506
rect 2433 -5540 2465 -5506
rect 2503 -5540 2535 -5506
rect 2535 -5540 2537 -5506
rect 2575 -5540 2603 -5506
rect 2603 -5540 2609 -5506
rect 2647 -5540 2671 -5506
rect 2671 -5540 2681 -5506
rect 2719 -5540 2739 -5506
rect 2739 -5540 2753 -5506
rect 2791 -5540 2807 -5506
rect 2807 -5540 2825 -5506
rect 2863 -5540 2875 -5506
rect 2875 -5540 2897 -5506
rect 2935 -5540 2943 -5506
rect 2943 -5540 2969 -5506
rect 3007 -5540 3011 -5506
rect 3011 -5540 3041 -5506
rect 3079 -5540 3113 -5506
rect 3151 -5540 3181 -5506
rect 3181 -5540 3185 -5506
rect 3223 -5540 3249 -5506
rect 3249 -5540 3257 -5506
rect 3295 -5540 3317 -5506
rect 3317 -5540 3329 -5506
rect 3367 -5540 3385 -5506
rect 3385 -5540 3401 -5506
rect 3439 -5540 3453 -5506
rect 3453 -5540 3473 -5506
rect 3511 -5540 3521 -5506
rect 3521 -5540 3545 -5506
rect 3583 -5540 3589 -5506
rect 3589 -5540 3617 -5506
rect 3655 -5540 3657 -5506
rect 3657 -5540 3689 -5506
rect 3727 -5540 3759 -5506
rect 3759 -5540 3761 -5506
rect 3799 -5540 3827 -5506
rect 3827 -5540 3833 -5506
rect 3871 -5540 3895 -5506
rect 3895 -5540 3905 -5506
rect 3943 -5540 3963 -5506
rect 3963 -5540 3977 -5506
rect 4015 -5540 4031 -5506
rect 4031 -5540 4049 -5506
rect 4087 -5540 4099 -5506
rect 4099 -5540 4121 -5506
rect 4159 -5540 4167 -5506
rect 4167 -5540 4193 -5506
rect 4231 -5540 4235 -5506
rect 4235 -5540 4265 -5506
rect 4303 -5540 4337 -5506
rect 4375 -5540 4405 -5506
rect 4405 -5540 4409 -5506
rect 4447 -5540 4473 -5506
rect 4473 -5540 4481 -5506
rect 4519 -5540 4541 -5506
rect 4541 -5540 4553 -5506
rect 4591 -5540 4609 -5506
rect 4609 -5540 4625 -5506
rect 4663 -5540 4677 -5506
rect 4677 -5540 4697 -5506
rect 4735 -5540 4745 -5506
rect 4745 -5540 4769 -5506
rect 4807 -5540 4813 -5506
rect 4813 -5540 4841 -5506
rect 4879 -5540 4881 -5506
rect 4881 -5540 4913 -5506
rect 4951 -5540 4983 -5506
rect 4983 -5540 4985 -5506
rect 5023 -5540 5051 -5506
rect 5051 -5540 5057 -5506
rect 5095 -5540 5119 -5506
rect 5119 -5540 5129 -5506
rect 5167 -5540 5187 -5506
rect 5187 -5540 5201 -5506
rect 5239 -5540 5255 -5506
rect 5255 -5540 5273 -5506
rect 5311 -5540 5323 -5506
rect 5323 -5540 5345 -5506
rect 5383 -5540 5391 -5506
rect 5391 -5540 5417 -5506
rect 5455 -5540 5459 -5506
rect 5459 -5540 5489 -5506
rect 5527 -5540 5561 -5506
rect 5599 -5540 5629 -5506
rect 5629 -5540 5633 -5506
rect 5671 -5540 5697 -5506
rect 5697 -5540 5705 -5506
rect 5743 -5540 5765 -5506
rect 5765 -5540 5777 -5506
rect 5815 -5540 5833 -5506
rect 5833 -5540 5849 -5506
rect 5887 -5540 5901 -5506
rect 5901 -5540 5921 -5506
rect 5959 -5540 5969 -5506
rect 5969 -5540 5993 -5506
<< metal1 >>
rect 315 5956 6191 5981
rect 315 5922 487 5956
rect 521 5922 559 5956
rect 593 5922 631 5956
rect 665 5922 703 5956
rect 737 5922 775 5956
rect 809 5922 847 5956
rect 881 5922 919 5956
rect 953 5922 991 5956
rect 1025 5922 1063 5956
rect 1097 5922 1135 5956
rect 1169 5922 1207 5956
rect 1241 5922 1279 5956
rect 1313 5922 1351 5956
rect 1385 5922 1423 5956
rect 1457 5922 1495 5956
rect 1529 5922 1567 5956
rect 1601 5922 1639 5956
rect 1673 5922 1711 5956
rect 1745 5922 1783 5956
rect 1817 5922 1855 5956
rect 1889 5922 1927 5956
rect 1961 5922 1999 5956
rect 2033 5922 2071 5956
rect 2105 5922 2143 5956
rect 2177 5922 2215 5956
rect 2249 5922 2287 5956
rect 2321 5922 2359 5956
rect 2393 5922 2431 5956
rect 2465 5922 2503 5956
rect 2537 5922 2575 5956
rect 2609 5922 2647 5956
rect 2681 5922 2719 5956
rect 2753 5922 2791 5956
rect 2825 5922 2863 5956
rect 2897 5922 2935 5956
rect 2969 5922 3007 5956
rect 3041 5922 3079 5956
rect 3113 5922 3151 5956
rect 3185 5922 3223 5956
rect 3257 5922 3295 5956
rect 3329 5922 3367 5956
rect 3401 5922 3439 5956
rect 3473 5922 3511 5956
rect 3545 5922 3583 5956
rect 3617 5922 3655 5956
rect 3689 5922 3727 5956
rect 3761 5922 3799 5956
rect 3833 5922 3871 5956
rect 3905 5922 3943 5956
rect 3977 5922 4015 5956
rect 4049 5922 4087 5956
rect 4121 5922 4159 5956
rect 4193 5922 4231 5956
rect 4265 5922 4303 5956
rect 4337 5922 4375 5956
rect 4409 5922 4447 5956
rect 4481 5922 4519 5956
rect 4553 5922 4591 5956
rect 4625 5922 4663 5956
rect 4697 5922 4735 5956
rect 4769 5922 4807 5956
rect 4841 5922 4879 5956
rect 4913 5922 4951 5956
rect 4985 5922 5023 5956
rect 5057 5922 5095 5956
rect 5129 5922 5167 5956
rect 5201 5922 5239 5956
rect 5273 5922 5311 5956
rect 5345 5922 5383 5956
rect 5417 5922 5455 5956
rect 5489 5922 5527 5956
rect 5561 5922 5599 5956
rect 5633 5922 5671 5956
rect 5705 5922 5743 5956
rect 5777 5922 5815 5956
rect 5849 5922 5887 5956
rect 5921 5922 5959 5956
rect 5993 5922 6191 5956
rect 315 5821 6191 5922
rect 315 5787 340 5821
rect 374 5787 6132 5821
rect 6166 5787 6191 5821
rect 315 5749 6191 5787
rect 315 5715 340 5749
rect 374 5742 6132 5749
rect 374 5715 530 5742
rect 315 5708 530 5715
rect 564 5708 788 5742
rect 822 5708 1046 5742
rect 1080 5708 1240 5742
rect 1274 5708 1498 5742
rect 1532 5708 1756 5742
rect 1790 5708 2014 5742
rect 2048 5708 2272 5742
rect 2306 5708 2466 5742
rect 2500 5708 2724 5742
rect 2758 5708 2982 5742
rect 3016 5708 3240 5742
rect 3274 5708 3498 5742
rect 3532 5708 3756 5742
rect 3790 5708 4014 5742
rect 4048 5708 4208 5742
rect 4242 5708 4466 5742
rect 4500 5708 4724 5742
rect 4758 5708 4982 5742
rect 5016 5708 5240 5742
rect 5274 5708 5433 5742
rect 5467 5708 5691 5742
rect 5725 5708 5949 5742
rect 5983 5715 6132 5742
rect 6166 5715 6191 5749
rect 5983 5708 6191 5715
rect 315 5677 6191 5708
rect 315 5643 340 5677
rect 374 5670 6132 5677
rect 374 5643 530 5670
rect 315 5636 530 5643
rect 564 5636 788 5670
rect 822 5636 1046 5670
rect 1080 5636 1240 5670
rect 1274 5636 1498 5670
rect 1532 5636 1756 5670
rect 1790 5636 2014 5670
rect 2048 5636 2272 5670
rect 2306 5636 2466 5670
rect 2500 5636 2724 5670
rect 2758 5636 2982 5670
rect 3016 5636 3240 5670
rect 3274 5636 3498 5670
rect 3532 5636 3756 5670
rect 3790 5636 4014 5670
rect 4048 5636 4208 5670
rect 4242 5636 4466 5670
rect 4500 5636 4724 5670
rect 4758 5636 4982 5670
rect 5016 5636 5240 5670
rect 5274 5636 5433 5670
rect 5467 5636 5691 5670
rect 5725 5636 5949 5670
rect 5983 5643 6132 5670
rect 6166 5643 6191 5677
rect 5983 5636 6191 5643
rect 315 5605 6191 5636
rect 315 5571 340 5605
rect 374 5571 6132 5605
rect 6166 5571 6191 5605
rect 315 5542 6191 5571
rect 315 5533 623 5542
rect 315 5499 340 5533
rect 374 5508 623 5533
rect 657 5508 695 5542
rect 729 5508 881 5542
rect 915 5508 953 5542
rect 987 5508 1333 5542
rect 1367 5508 1405 5542
rect 1439 5508 1591 5542
rect 1625 5508 1663 5542
rect 1697 5508 1849 5542
rect 1883 5508 1921 5542
rect 1955 5508 2107 5542
rect 2141 5508 2179 5542
rect 2213 5508 2559 5542
rect 2593 5508 2631 5542
rect 2665 5508 2817 5542
rect 2851 5508 2889 5542
rect 2923 5508 3075 5542
rect 3109 5508 3147 5542
rect 3181 5508 3333 5542
rect 3367 5508 3405 5542
rect 3439 5508 3591 5542
rect 3625 5508 3663 5542
rect 3697 5508 3849 5542
rect 3883 5508 3921 5542
rect 3955 5508 4301 5542
rect 4335 5508 4373 5542
rect 4407 5508 4559 5542
rect 4593 5508 4631 5542
rect 4665 5508 4817 5542
rect 4851 5508 4889 5542
rect 4923 5508 5075 5542
rect 5109 5508 5147 5542
rect 5181 5508 5526 5542
rect 5560 5508 5598 5542
rect 5632 5508 5784 5542
rect 5818 5508 5856 5542
rect 5890 5533 6191 5542
rect 5890 5508 6132 5533
rect 374 5502 6132 5508
rect 374 5499 1098 5502
rect 315 5461 1098 5499
rect 315 5427 340 5461
rect 374 5427 1098 5461
rect 315 5389 1098 5427
rect 315 5355 340 5389
rect 374 5355 1098 5389
rect 5427 5499 6132 5502
rect 6166 5499 6191 5533
rect 5427 5461 6191 5499
rect 5427 5427 6132 5461
rect 6166 5427 6191 5461
rect 5427 5389 6191 5427
rect 315 5317 1098 5355
rect 315 5283 340 5317
rect 374 5283 1098 5317
rect 315 5261 1098 5283
rect 315 5245 623 5261
rect 315 5211 340 5245
rect 374 5227 623 5245
rect 657 5227 695 5261
rect 729 5227 881 5261
rect 915 5227 953 5261
rect 987 5227 1098 5261
rect 374 5211 1098 5227
rect 1290 5348 1740 5356
rect 1290 5296 1421 5348
rect 1473 5296 1485 5348
rect 1537 5296 1549 5348
rect 1601 5296 1740 5348
rect 1290 5224 1740 5296
rect 1806 5348 2256 5356
rect 1806 5296 1937 5348
rect 1989 5296 2001 5348
rect 2053 5296 2065 5348
rect 2117 5296 2256 5348
rect 1806 5224 2256 5296
rect 2516 5348 2966 5356
rect 2516 5296 2647 5348
rect 2699 5296 2711 5348
rect 2763 5296 2775 5348
rect 2827 5296 2966 5348
rect 2516 5224 2966 5296
rect 3032 5348 3482 5356
rect 3032 5296 3163 5348
rect 3215 5296 3227 5348
rect 3279 5296 3291 5348
rect 3343 5296 3482 5348
rect 3032 5224 3482 5296
rect 3548 5348 3998 5356
rect 3548 5296 3679 5348
rect 3731 5296 3743 5348
rect 3795 5296 3807 5348
rect 3859 5296 3998 5348
rect 3548 5224 3998 5296
rect 4258 5348 4708 5356
rect 4258 5296 4389 5348
rect 4441 5296 4453 5348
rect 4505 5296 4517 5348
rect 4569 5296 4708 5348
rect 4258 5224 4708 5296
rect 4774 5348 5224 5356
rect 4774 5296 4905 5348
rect 4957 5296 4969 5348
rect 5021 5296 5033 5348
rect 5085 5296 5224 5348
rect 4774 5224 5224 5296
rect 5427 5355 6132 5389
rect 6166 5355 6191 5389
rect 5427 5317 6191 5355
rect 5427 5283 6132 5317
rect 6166 5283 6191 5317
rect 5427 5261 6191 5283
rect 5427 5227 5526 5261
rect 5560 5227 5598 5261
rect 5632 5227 5784 5261
rect 5818 5227 5856 5261
rect 5890 5245 6191 5261
rect 5890 5227 6132 5245
rect 315 5173 1098 5211
rect 315 5139 340 5173
rect 374 5139 1098 5173
rect 315 5133 1098 5139
rect 315 5101 530 5133
rect 315 5067 340 5101
rect 374 5099 530 5101
rect 564 5099 788 5133
rect 822 5099 1046 5133
rect 1080 5099 1098 5133
rect 374 5067 1098 5099
rect 5427 5211 6132 5227
rect 6166 5211 6191 5245
rect 5427 5173 6191 5211
rect 5427 5139 6132 5173
rect 6166 5139 6191 5173
rect 5427 5133 6191 5139
rect 5427 5099 5433 5133
rect 5467 5099 5691 5133
rect 5725 5099 5949 5133
rect 5983 5101 6191 5133
rect 5983 5099 6132 5101
rect 315 5061 1098 5067
rect 315 5029 530 5061
rect 315 4995 340 5029
rect 374 5027 530 5029
rect 564 5027 788 5061
rect 822 5027 1046 5061
rect 1080 5027 1098 5061
rect 374 4995 1098 5027
rect 315 4957 1098 4995
rect 315 4923 340 4957
rect 374 4923 1098 4957
rect 315 4885 1098 4923
rect 315 4851 340 4885
rect 374 4851 1098 4885
rect 315 4813 1098 4851
rect 315 4779 340 4813
rect 374 4779 1098 4813
rect 315 4741 1098 4779
rect 315 4707 340 4741
rect 374 4707 1098 4741
rect 315 4672 1098 4707
rect 1234 4672 1280 4990
rect 1750 4951 1796 5081
rect 1672 4943 1868 4951
rect 1672 4891 1681 4943
rect 1733 4891 1745 4943
rect 1797 4891 1809 4943
rect 1861 4891 1868 4943
rect 1672 4881 1868 4891
rect 2266 4672 2312 4990
rect 2460 4811 2506 5081
rect 2460 4803 2656 4811
rect 2460 4751 2469 4803
rect 2521 4751 2533 4803
rect 2585 4751 2597 4803
rect 2649 4751 2656 4803
rect 2460 4741 2656 4751
rect 2976 4672 3022 4990
rect 3492 4811 3538 5081
rect 3417 4803 3613 4811
rect 3417 4751 3424 4803
rect 3476 4751 3488 4803
rect 3540 4751 3552 4803
rect 3604 4751 3613 4803
rect 3417 4741 3613 4751
rect 4008 4672 4054 4990
rect 4202 4672 4248 4990
rect 4718 4951 4764 5081
rect 5427 5067 6132 5099
rect 6166 5067 6191 5101
rect 5427 5061 6191 5067
rect 5427 5027 5433 5061
rect 5467 5027 5691 5061
rect 5725 5027 5949 5061
rect 5983 5029 6191 5061
rect 5983 5027 6132 5029
rect 5427 4995 6132 5027
rect 6166 4995 6191 5029
rect 4642 4943 4838 4951
rect 4642 4891 4651 4943
rect 4703 4891 4715 4943
rect 4767 4891 4779 4943
rect 4831 4891 4838 4943
rect 4642 4881 4838 4891
rect 315 4669 1280 4672
rect 315 4635 340 4669
rect 374 4662 1280 4669
rect 374 4635 1074 4662
rect 315 4610 1074 4635
rect 1126 4610 1138 4662
rect 1190 4610 1202 4662
rect 1254 4610 1280 4662
rect 315 4602 1280 4610
rect 2108 4662 2312 4672
rect 2108 4610 2117 4662
rect 2169 4610 2181 4662
rect 2233 4610 2245 4662
rect 2297 4610 2312 4662
rect 2108 4602 2312 4610
rect 2914 4662 3110 4672
rect 2914 4610 2921 4662
rect 2973 4610 2985 4662
rect 3037 4610 3049 4662
rect 3101 4610 3110 4662
rect 2914 4602 3110 4610
rect 4008 4662 4248 4672
rect 4008 4610 4034 4662
rect 4086 4610 4098 4662
rect 4150 4610 4162 4662
rect 4214 4610 4248 4662
rect 4008 4602 4248 4610
rect 315 4597 1098 4602
rect 315 4563 340 4597
rect 374 4563 1098 4597
rect 315 4525 1098 4563
rect 315 4491 340 4525
rect 374 4491 1098 4525
rect 315 4453 1098 4491
rect 315 4419 340 4453
rect 374 4419 1098 4453
rect 315 4381 1098 4419
rect 315 4347 340 4381
rect 374 4347 1098 4381
rect 315 4309 1098 4347
rect 315 4275 340 4309
rect 374 4275 1098 4309
rect 315 4238 1098 4275
rect 315 4237 530 4238
rect 315 4203 340 4237
rect 374 4204 530 4237
rect 564 4204 788 4238
rect 822 4204 1046 4238
rect 1080 4204 1098 4238
rect 374 4203 1098 4204
rect 315 4166 1098 4203
rect 315 4165 530 4166
rect 315 4131 340 4165
rect 374 4132 530 4165
rect 564 4132 788 4166
rect 822 4132 1046 4166
rect 1080 4132 1098 4166
rect 1234 4164 1280 4602
rect 1672 4383 1868 4393
rect 1672 4331 1681 4383
rect 1733 4331 1745 4383
rect 1797 4331 1809 4383
rect 1861 4331 1868 4383
rect 1672 4323 1868 4331
rect 1750 4193 1796 4323
rect 2266 4164 2312 4602
rect 2460 4524 2656 4532
rect 2460 4472 2469 4524
rect 2521 4472 2533 4524
rect 2585 4472 2597 4524
rect 2649 4472 2656 4524
rect 2460 4462 2656 4472
rect 2460 4193 2506 4462
rect 2976 4164 3022 4602
rect 3417 4524 3613 4532
rect 3417 4472 3424 4524
rect 3476 4472 3488 4524
rect 3540 4472 3552 4524
rect 3604 4472 3613 4524
rect 3417 4462 3613 4472
rect 3492 4193 3538 4462
rect 4008 4165 4054 4602
rect 4202 4165 4248 4602
rect 5234 4672 5280 4990
rect 5427 4957 6191 4995
rect 5427 4923 6132 4957
rect 6166 4923 6191 4957
rect 5427 4885 6191 4923
rect 5427 4851 6132 4885
rect 6166 4851 6191 4885
rect 5427 4813 6191 4851
rect 5427 4779 6132 4813
rect 6166 4779 6191 4813
rect 5427 4741 6191 4779
rect 5427 4707 6132 4741
rect 6166 4707 6191 4741
rect 5427 4672 6191 4707
rect 5234 4669 6191 4672
rect 5234 4662 6132 4669
rect 5234 4610 5262 4662
rect 5314 4610 5326 4662
rect 5378 4610 5390 4662
rect 5442 4635 6132 4662
rect 6166 4635 6191 4669
rect 5442 4610 6191 4635
rect 5234 4602 6191 4610
rect 4642 4383 4838 4393
rect 4642 4331 4651 4383
rect 4703 4331 4715 4383
rect 4767 4331 4779 4383
rect 4831 4331 4838 4383
rect 4642 4323 4838 4331
rect 4718 4193 4764 4323
rect 5234 4165 5280 4602
rect 5427 4597 6191 4602
rect 5427 4563 6132 4597
rect 6166 4563 6191 4597
rect 5427 4525 6191 4563
rect 5427 4491 6132 4525
rect 6166 4491 6191 4525
rect 5427 4453 6191 4491
rect 5427 4419 6132 4453
rect 6166 4419 6191 4453
rect 5427 4381 6191 4419
rect 5427 4347 6132 4381
rect 6166 4347 6191 4381
rect 5427 4309 6191 4347
rect 5427 4275 6132 4309
rect 6166 4275 6191 4309
rect 5427 4238 6191 4275
rect 5427 4204 5433 4238
rect 5467 4204 5691 4238
rect 5725 4204 5949 4238
rect 5983 4237 6191 4238
rect 5983 4204 6132 4237
rect 5427 4203 6132 4204
rect 6166 4203 6191 4237
rect 5427 4166 6191 4203
rect 374 4131 1098 4132
rect 315 4093 1098 4131
rect 315 4059 340 4093
rect 374 4059 1098 4093
rect 315 4038 1098 4059
rect 5427 4132 5433 4166
rect 5467 4132 5691 4166
rect 5725 4132 5949 4166
rect 5983 4165 6191 4166
rect 5983 4132 6132 4165
rect 5427 4131 6132 4132
rect 6166 4131 6191 4165
rect 5427 4093 6191 4131
rect 5427 4059 6132 4093
rect 6166 4059 6191 4093
rect 315 4021 623 4038
rect 315 3987 340 4021
rect 374 4004 623 4021
rect 657 4004 695 4038
rect 729 4004 881 4038
rect 915 4004 953 4038
rect 987 4004 1098 4038
rect 374 3987 1098 4004
rect 315 3949 1098 3987
rect 315 3915 340 3949
rect 374 3915 1098 3949
rect 1290 3982 1740 4054
rect 1290 3930 1421 3982
rect 1473 3930 1485 3982
rect 1537 3930 1549 3982
rect 1601 3930 1740 3982
rect 1290 3922 1740 3930
rect 1806 3982 2256 4054
rect 1806 3930 1937 3982
rect 1989 3930 2001 3982
rect 2053 3930 2065 3982
rect 2117 3930 2256 3982
rect 1806 3922 2256 3930
rect 2516 3982 2966 4054
rect 2516 3930 2647 3982
rect 2699 3930 2711 3982
rect 2763 3930 2775 3982
rect 2827 3930 2966 3982
rect 2516 3922 2966 3930
rect 3032 3982 3482 4054
rect 3032 3930 3163 3982
rect 3215 3930 3227 3982
rect 3279 3930 3291 3982
rect 3343 3930 3482 3982
rect 3032 3922 3482 3930
rect 3548 3982 3998 4054
rect 3548 3930 3679 3982
rect 3731 3930 3743 3982
rect 3795 3930 3807 3982
rect 3859 3930 3998 3982
rect 3548 3922 3998 3930
rect 4258 3982 4708 4054
rect 4258 3930 4389 3982
rect 4441 3930 4453 3982
rect 4505 3930 4517 3982
rect 4569 3930 4708 3982
rect 4258 3922 4708 3930
rect 4774 3982 5224 4054
rect 4774 3930 4905 3982
rect 4957 3930 4969 3982
rect 5021 3930 5033 3982
rect 5085 3930 5224 3982
rect 4774 3922 5224 3930
rect 5427 4038 6191 4059
rect 5427 4004 5526 4038
rect 5560 4004 5598 4038
rect 5632 4004 5784 4038
rect 5818 4004 5856 4038
rect 5890 4021 6191 4038
rect 5890 4004 6132 4021
rect 5427 3987 6132 4004
rect 6166 3987 6191 4021
rect 5427 3949 6191 3987
rect 315 3877 1098 3915
rect 315 3843 340 3877
rect 374 3843 1098 3877
rect 5427 3915 6132 3949
rect 6166 3915 6191 3949
rect 5427 3877 6191 3915
rect 315 3805 1098 3843
rect 315 3771 340 3805
rect 374 3771 1098 3805
rect 315 3757 1098 3771
rect 315 3733 623 3757
rect 315 3699 340 3733
rect 374 3723 623 3733
rect 657 3723 695 3757
rect 729 3723 881 3757
rect 915 3723 953 3757
rect 987 3723 1098 3757
rect 374 3699 1098 3723
rect 1290 3844 1740 3852
rect 1290 3792 1421 3844
rect 1473 3792 1485 3844
rect 1537 3792 1549 3844
rect 1601 3792 1740 3844
rect 1290 3720 1740 3792
rect 1806 3844 2256 3852
rect 1806 3792 1937 3844
rect 1989 3792 2001 3844
rect 2053 3792 2065 3844
rect 2117 3792 2256 3844
rect 1806 3720 2256 3792
rect 2516 3844 2966 3852
rect 2516 3792 2647 3844
rect 2699 3792 2711 3844
rect 2763 3792 2775 3844
rect 2827 3792 2966 3844
rect 2516 3720 2966 3792
rect 3032 3844 3482 3852
rect 3032 3792 3163 3844
rect 3215 3792 3227 3844
rect 3279 3792 3291 3844
rect 3343 3792 3482 3844
rect 3032 3720 3482 3792
rect 3548 3844 3998 3852
rect 3548 3792 3679 3844
rect 3731 3792 3743 3844
rect 3795 3792 3807 3844
rect 3859 3792 3998 3844
rect 3548 3720 3998 3792
rect 4258 3844 4708 3852
rect 4258 3792 4389 3844
rect 4441 3792 4453 3844
rect 4505 3792 4517 3844
rect 4569 3792 4708 3844
rect 4258 3720 4708 3792
rect 4774 3844 5224 3852
rect 4774 3792 4905 3844
rect 4957 3792 4969 3844
rect 5021 3792 5033 3844
rect 5085 3792 5224 3844
rect 4774 3720 5224 3792
rect 5427 3843 6132 3877
rect 6166 3843 6191 3877
rect 5427 3805 6191 3843
rect 5427 3771 6132 3805
rect 6166 3771 6191 3805
rect 5427 3757 6191 3771
rect 5427 3723 5526 3757
rect 5560 3723 5598 3757
rect 5632 3723 5784 3757
rect 5818 3723 5856 3757
rect 5890 3733 6191 3757
rect 5890 3723 6132 3733
rect 315 3661 1098 3699
rect 315 3627 340 3661
rect 374 3629 1098 3661
rect 374 3627 530 3629
rect 315 3595 530 3627
rect 564 3595 788 3629
rect 822 3595 1046 3629
rect 1080 3595 1098 3629
rect 315 3589 1098 3595
rect 315 3555 340 3589
rect 374 3557 1098 3589
rect 5427 3699 6132 3723
rect 6166 3699 6191 3733
rect 5427 3661 6191 3699
rect 5427 3629 6132 3661
rect 5427 3595 5433 3629
rect 5467 3595 5691 3629
rect 5725 3595 5949 3629
rect 5983 3627 6132 3629
rect 6166 3627 6191 3661
rect 5983 3595 6191 3627
rect 5427 3589 6191 3595
rect 374 3555 530 3557
rect 315 3523 530 3555
rect 564 3523 788 3557
rect 822 3523 1046 3557
rect 1080 3523 1098 3557
rect 315 3517 1098 3523
rect 315 3483 340 3517
rect 374 3483 1098 3517
rect 315 3445 1098 3483
rect 315 3411 340 3445
rect 374 3411 1098 3445
rect 315 3373 1098 3411
rect 315 3339 340 3373
rect 374 3339 1098 3373
rect 315 3301 1098 3339
rect 315 3267 340 3301
rect 374 3267 1098 3301
rect 315 3229 1098 3267
rect 315 3195 340 3229
rect 374 3195 1098 3229
rect 315 3168 1098 3195
rect 1234 3168 1280 3486
rect 1750 3447 1796 3577
rect 1672 3439 1868 3447
rect 1672 3387 1681 3439
rect 1733 3387 1745 3439
rect 1797 3387 1809 3439
rect 1861 3387 1868 3439
rect 1672 3377 1868 3387
rect 2266 3168 2312 3486
rect 2460 3307 2506 3577
rect 2460 3299 2656 3307
rect 2460 3247 2469 3299
rect 2521 3247 2533 3299
rect 2585 3247 2597 3299
rect 2649 3247 2656 3299
rect 2460 3237 2656 3247
rect 2976 3168 3022 3486
rect 3492 3307 3538 3577
rect 3417 3299 3613 3307
rect 3417 3247 3424 3299
rect 3476 3247 3488 3299
rect 3540 3247 3552 3299
rect 3604 3247 3613 3299
rect 3417 3237 3613 3247
rect 4008 3168 4054 3486
rect 4202 3168 4248 3486
rect 4718 3447 4764 3577
rect 5427 3557 6132 3589
rect 5427 3523 5433 3557
rect 5467 3523 5691 3557
rect 5725 3523 5949 3557
rect 5983 3555 6132 3557
rect 6166 3555 6191 3589
rect 5983 3523 6191 3555
rect 5427 3517 6191 3523
rect 4642 3439 4838 3447
rect 4642 3387 4651 3439
rect 4703 3387 4715 3439
rect 4767 3387 4779 3439
rect 4831 3387 4838 3439
rect 4642 3377 4838 3387
rect 315 3158 1280 3168
rect 315 3157 1074 3158
rect 315 3123 340 3157
rect 374 3123 1074 3157
rect 315 3106 1074 3123
rect 1126 3106 1138 3158
rect 1190 3106 1202 3158
rect 1254 3106 1280 3158
rect 315 3098 1280 3106
rect 2108 3158 2312 3168
rect 2108 3106 2117 3158
rect 2169 3106 2181 3158
rect 2233 3106 2245 3158
rect 2297 3106 2312 3158
rect 2108 3098 2312 3106
rect 2914 3158 3110 3168
rect 2914 3106 2921 3158
rect 2973 3106 2985 3158
rect 3037 3106 3049 3158
rect 3101 3106 3110 3158
rect 2914 3098 3110 3106
rect 4008 3158 4248 3168
rect 4008 3106 4034 3158
rect 4086 3106 4098 3158
rect 4150 3106 4162 3158
rect 4214 3106 4248 3158
rect 4008 3098 4248 3106
rect 315 3085 1098 3098
rect 315 3051 340 3085
rect 374 3051 1098 3085
rect 315 3013 1098 3051
rect 315 2979 340 3013
rect 374 2979 1098 3013
rect 315 2941 1098 2979
rect 315 2907 340 2941
rect 374 2907 1098 2941
rect 315 2869 1098 2907
rect 315 2835 340 2869
rect 374 2835 1098 2869
rect 315 2797 1098 2835
rect 315 2763 340 2797
rect 374 2763 1098 2797
rect 315 2731 1098 2763
rect 315 2725 530 2731
rect 315 2691 340 2725
rect 374 2697 530 2725
rect 564 2697 788 2731
rect 822 2697 1046 2731
rect 1080 2697 1098 2731
rect 374 2691 1098 2697
rect 315 2659 1098 2691
rect 1234 2660 1280 3098
rect 1672 2879 1868 2889
rect 1672 2827 1681 2879
rect 1733 2827 1745 2879
rect 1797 2827 1809 2879
rect 1861 2827 1868 2879
rect 1672 2819 1868 2827
rect 1750 2689 1796 2819
rect 2266 2660 2312 3098
rect 2460 3020 2656 3028
rect 2460 2968 2469 3020
rect 2521 2968 2533 3020
rect 2585 2968 2597 3020
rect 2649 2968 2656 3020
rect 2460 2958 2656 2968
rect 2460 2689 2506 2958
rect 2976 2660 3022 3098
rect 3417 3020 3613 3028
rect 3417 2968 3424 3020
rect 3476 2968 3488 3020
rect 3540 2968 3552 3020
rect 3604 2968 3613 3020
rect 3417 2958 3613 2968
rect 3492 2689 3538 2958
rect 4008 2661 4054 3098
rect 4202 2661 4248 3098
rect 5234 3168 5280 3486
rect 5427 3483 6132 3517
rect 6166 3483 6191 3517
rect 5427 3445 6191 3483
rect 5427 3411 6132 3445
rect 6166 3411 6191 3445
rect 5427 3373 6191 3411
rect 5427 3339 6132 3373
rect 6166 3339 6191 3373
rect 5427 3301 6191 3339
rect 5427 3267 6132 3301
rect 6166 3267 6191 3301
rect 5427 3229 6191 3267
rect 5427 3195 6132 3229
rect 6166 3195 6191 3229
rect 5427 3168 6191 3195
rect 5234 3158 6191 3168
rect 5234 3106 5262 3158
rect 5314 3106 5326 3158
rect 5378 3106 5390 3158
rect 5442 3157 6191 3158
rect 5442 3123 6132 3157
rect 6166 3123 6191 3157
rect 5442 3106 6191 3123
rect 5234 3098 6191 3106
rect 4642 2879 4838 2889
rect 4642 2827 4651 2879
rect 4703 2827 4715 2879
rect 4767 2827 4779 2879
rect 4831 2827 4838 2879
rect 4642 2819 4838 2827
rect 4718 2689 4764 2819
rect 5234 2661 5280 3098
rect 5427 3085 6191 3098
rect 5427 3051 6132 3085
rect 6166 3051 6191 3085
rect 5427 3013 6191 3051
rect 5427 2979 6132 3013
rect 6166 2979 6191 3013
rect 5427 2941 6191 2979
rect 5427 2907 6132 2941
rect 6166 2907 6191 2941
rect 5427 2869 6191 2907
rect 5427 2835 6132 2869
rect 6166 2835 6191 2869
rect 5427 2797 6191 2835
rect 5427 2763 6132 2797
rect 6166 2763 6191 2797
rect 5427 2731 6191 2763
rect 5427 2697 5433 2731
rect 5467 2697 5691 2731
rect 5725 2697 5949 2731
rect 5983 2725 6191 2731
rect 5983 2697 6132 2725
rect 5427 2691 6132 2697
rect 6166 2691 6191 2725
rect 315 2653 530 2659
rect 315 2619 340 2653
rect 374 2625 530 2653
rect 564 2625 788 2659
rect 822 2625 1046 2659
rect 1080 2625 1098 2659
rect 374 2619 1098 2625
rect 315 2581 1098 2619
rect 315 2547 340 2581
rect 374 2547 1098 2581
rect 5427 2659 6191 2691
rect 5427 2625 5433 2659
rect 5467 2625 5691 2659
rect 5725 2625 5949 2659
rect 5983 2653 6191 2659
rect 5983 2625 6132 2653
rect 5427 2619 6132 2625
rect 6166 2619 6191 2653
rect 5427 2581 6191 2619
rect 315 2531 1098 2547
rect 315 2509 623 2531
rect 315 2475 340 2509
rect 374 2497 623 2509
rect 657 2497 695 2531
rect 729 2497 881 2531
rect 915 2497 953 2531
rect 987 2497 1098 2531
rect 374 2475 1098 2497
rect 315 2437 1098 2475
rect 315 2403 340 2437
rect 374 2403 1098 2437
rect 1290 2478 1740 2550
rect 1290 2426 1421 2478
rect 1473 2426 1485 2478
rect 1537 2426 1549 2478
rect 1601 2426 1740 2478
rect 1290 2418 1740 2426
rect 1806 2478 2256 2550
rect 1806 2426 1937 2478
rect 1989 2426 2001 2478
rect 2053 2426 2065 2478
rect 2117 2426 2256 2478
rect 1806 2418 2256 2426
rect 2516 2478 2966 2550
rect 2516 2426 2647 2478
rect 2699 2426 2711 2478
rect 2763 2426 2775 2478
rect 2827 2426 2966 2478
rect 2516 2418 2966 2426
rect 3032 2478 3482 2550
rect 3032 2426 3163 2478
rect 3215 2426 3227 2478
rect 3279 2426 3291 2478
rect 3343 2426 3482 2478
rect 3032 2418 3482 2426
rect 3548 2478 3998 2550
rect 3548 2426 3679 2478
rect 3731 2426 3743 2478
rect 3795 2426 3807 2478
rect 3859 2426 3998 2478
rect 3548 2418 3998 2426
rect 4258 2478 4708 2550
rect 4258 2426 4389 2478
rect 4441 2426 4453 2478
rect 4505 2426 4517 2478
rect 4569 2426 4708 2478
rect 4258 2418 4708 2426
rect 4774 2478 5224 2550
rect 4774 2426 4905 2478
rect 4957 2426 4969 2478
rect 5021 2426 5033 2478
rect 5085 2426 5224 2478
rect 4774 2418 5224 2426
rect 5427 2547 6132 2581
rect 6166 2547 6191 2581
rect 5427 2531 6191 2547
rect 5427 2497 5526 2531
rect 5560 2497 5598 2531
rect 5632 2497 5784 2531
rect 5818 2497 5856 2531
rect 5890 2509 6191 2531
rect 5890 2497 6132 2509
rect 5427 2475 6132 2497
rect 6166 2475 6191 2509
rect 5427 2437 6191 2475
rect 315 2365 1098 2403
rect 315 2331 340 2365
rect 374 2331 1098 2365
rect 5427 2403 6132 2437
rect 6166 2403 6191 2437
rect 5427 2365 6191 2403
rect 315 2293 1098 2331
rect 315 2259 340 2293
rect 374 2259 1098 2293
rect 315 2250 1098 2259
rect 315 2221 623 2250
rect 315 2187 340 2221
rect 374 2216 623 2221
rect 657 2216 695 2250
rect 729 2216 881 2250
rect 915 2216 953 2250
rect 987 2216 1098 2250
rect 374 2187 1098 2216
rect 1290 2330 1740 2338
rect 1290 2278 1421 2330
rect 1473 2278 1485 2330
rect 1537 2278 1549 2330
rect 1601 2278 1740 2330
rect 1290 2206 1740 2278
rect 1806 2330 2256 2338
rect 1806 2278 1937 2330
rect 1989 2278 2001 2330
rect 2053 2278 2065 2330
rect 2117 2278 2256 2330
rect 1806 2206 2256 2278
rect 2516 2330 2966 2338
rect 2516 2278 2647 2330
rect 2699 2278 2711 2330
rect 2763 2278 2775 2330
rect 2827 2278 2966 2330
rect 2516 2206 2966 2278
rect 3032 2330 3482 2338
rect 3032 2278 3163 2330
rect 3215 2278 3227 2330
rect 3279 2278 3291 2330
rect 3343 2278 3482 2330
rect 3032 2206 3482 2278
rect 3548 2330 3998 2338
rect 3548 2278 3679 2330
rect 3731 2278 3743 2330
rect 3795 2278 3807 2330
rect 3859 2278 3998 2330
rect 3548 2206 3998 2278
rect 4258 2330 4708 2338
rect 4258 2278 4389 2330
rect 4441 2278 4453 2330
rect 4505 2278 4517 2330
rect 4569 2278 4708 2330
rect 4258 2206 4708 2278
rect 4774 2330 5224 2338
rect 4774 2278 4905 2330
rect 4957 2278 4969 2330
rect 5021 2278 5033 2330
rect 5085 2278 5224 2330
rect 4774 2206 5224 2278
rect 5427 2331 6132 2365
rect 6166 2331 6191 2365
rect 5427 2293 6191 2331
rect 5427 2259 6132 2293
rect 6166 2259 6191 2293
rect 5427 2250 6191 2259
rect 5427 2216 5526 2250
rect 5560 2216 5598 2250
rect 5632 2216 5784 2250
rect 5818 2216 5856 2250
rect 5890 2221 6191 2250
rect 5890 2216 6132 2221
rect 315 2149 1098 2187
rect 315 2115 340 2149
rect 374 2122 1098 2149
rect 374 2115 530 2122
rect 315 2088 530 2115
rect 564 2088 788 2122
rect 822 2088 1046 2122
rect 1080 2088 1098 2122
rect 315 2077 1098 2088
rect 315 2043 340 2077
rect 374 2050 1098 2077
rect 5427 2187 6132 2216
rect 6166 2187 6191 2221
rect 5427 2149 6191 2187
rect 5427 2122 6132 2149
rect 5427 2088 5433 2122
rect 5467 2088 5691 2122
rect 5725 2088 5949 2122
rect 5983 2115 6132 2122
rect 6166 2115 6191 2149
rect 5983 2088 6191 2115
rect 5427 2077 6191 2088
rect 374 2043 530 2050
rect 315 2016 530 2043
rect 564 2016 788 2050
rect 822 2016 1046 2050
rect 1080 2016 1098 2050
rect 315 1928 1098 2016
rect 315 1894 340 1928
rect 374 1894 1098 1928
rect 315 1856 1098 1894
rect 315 1822 340 1856
rect 374 1822 1098 1856
rect 315 1784 1098 1822
rect 315 1750 340 1784
rect 374 1750 1098 1784
rect 315 1712 1098 1750
rect 315 1678 340 1712
rect 374 1678 1098 1712
rect 315 1660 1098 1678
rect 1234 1660 1280 1978
rect 1750 1939 1796 2069
rect 1672 1931 1868 1939
rect 1672 1879 1681 1931
rect 1733 1879 1745 1931
rect 1797 1879 1809 1931
rect 1861 1879 1868 1931
rect 1672 1869 1868 1879
rect 2266 1660 2312 1978
rect 2460 1799 2506 2069
rect 2460 1791 2656 1799
rect 2460 1739 2469 1791
rect 2521 1739 2533 1791
rect 2585 1739 2597 1791
rect 2649 1739 2656 1791
rect 2460 1729 2656 1739
rect 2976 1660 3022 1978
rect 3492 1799 3538 2069
rect 3417 1791 3613 1799
rect 3417 1739 3424 1791
rect 3476 1739 3488 1791
rect 3540 1739 3552 1791
rect 3604 1739 3613 1791
rect 3417 1729 3613 1739
rect 4008 1660 4054 1978
rect 4202 1660 4248 1978
rect 4718 1939 4764 2069
rect 5427 2050 6132 2077
rect 5427 2016 5433 2050
rect 5467 2016 5691 2050
rect 5725 2016 5949 2050
rect 5983 2043 6132 2050
rect 6166 2043 6191 2077
rect 5983 2016 6191 2043
rect 4642 1931 4838 1939
rect 4642 1879 4651 1931
rect 4703 1879 4715 1931
rect 4767 1879 4779 1931
rect 4831 1879 4838 1931
rect 4642 1869 4838 1879
rect 315 1650 1280 1660
rect 315 1640 1074 1650
rect 315 1606 340 1640
rect 374 1606 1074 1640
rect 315 1598 1074 1606
rect 1126 1598 1138 1650
rect 1190 1598 1202 1650
rect 1254 1598 1280 1650
rect 315 1590 1280 1598
rect 2108 1650 2312 1660
rect 2108 1598 2117 1650
rect 2169 1598 2181 1650
rect 2233 1598 2245 1650
rect 2297 1598 2312 1650
rect 2108 1590 2312 1598
rect 2914 1650 3110 1660
rect 2914 1598 2921 1650
rect 2973 1598 2985 1650
rect 3037 1598 3049 1650
rect 3101 1598 3110 1650
rect 2914 1590 3110 1598
rect 4008 1650 4248 1660
rect 4008 1598 4034 1650
rect 4086 1598 4098 1650
rect 4150 1598 4162 1650
rect 4214 1598 4248 1650
rect 4008 1590 4248 1598
rect 315 1568 1098 1590
rect 315 1534 340 1568
rect 374 1534 1098 1568
rect 315 1496 1098 1534
rect 315 1462 340 1496
rect 374 1462 1098 1496
rect 315 1424 1098 1462
rect 315 1390 340 1424
rect 374 1390 1098 1424
rect 315 1362 1098 1390
rect 315 1352 530 1362
rect 315 1318 340 1352
rect 374 1328 530 1352
rect 564 1328 788 1362
rect 822 1328 1046 1362
rect 1080 1328 1098 1362
rect 374 1318 1098 1328
rect 315 1290 1098 1318
rect 1234 1292 1280 1590
rect 1672 1510 1868 1520
rect 1672 1458 1681 1510
rect 1733 1458 1745 1510
rect 1797 1458 1809 1510
rect 1861 1458 1868 1510
rect 1672 1450 1868 1458
rect 1750 1320 1796 1450
rect 2266 1292 2312 1590
rect 2460 1510 2665 1520
rect 2460 1458 2478 1510
rect 2530 1458 2542 1510
rect 2594 1458 2606 1510
rect 2658 1458 2665 1510
rect 2460 1450 2665 1458
rect 2460 1320 2506 1450
rect 2976 1292 3022 1590
rect 3417 1510 3613 1520
rect 3417 1458 3424 1510
rect 3476 1458 3488 1510
rect 3540 1458 3552 1510
rect 3604 1458 3613 1510
rect 3417 1450 3613 1458
rect 3492 1320 3538 1450
rect 4008 1292 4054 1590
rect 4202 1292 4248 1590
rect 5234 1660 5280 1978
rect 5427 1928 6191 2016
rect 5427 1894 6132 1928
rect 6166 1894 6191 1928
rect 5427 1856 6191 1894
rect 5427 1822 6132 1856
rect 6166 1822 6191 1856
rect 5427 1784 6191 1822
rect 5427 1750 6132 1784
rect 6166 1750 6191 1784
rect 5427 1712 6191 1750
rect 5427 1678 6132 1712
rect 6166 1678 6191 1712
rect 5427 1660 6191 1678
rect 5234 1650 6191 1660
rect 5234 1598 5262 1650
rect 5314 1598 5326 1650
rect 5378 1598 5390 1650
rect 5442 1640 6191 1650
rect 5442 1606 6132 1640
rect 6166 1606 6191 1640
rect 5442 1598 6191 1606
rect 5234 1590 6191 1598
rect 4642 1510 4838 1520
rect 4642 1458 4651 1510
rect 4703 1458 4715 1510
rect 4767 1458 4779 1510
rect 4831 1458 4838 1510
rect 4642 1450 4838 1458
rect 4718 1320 4764 1450
rect 5234 1292 5280 1590
rect 5427 1568 6191 1590
rect 5427 1534 6132 1568
rect 6166 1534 6191 1568
rect 5427 1496 6191 1534
rect 5427 1462 6132 1496
rect 6166 1462 6191 1496
rect 5427 1424 6191 1462
rect 5427 1390 6132 1424
rect 6166 1390 6191 1424
rect 5427 1362 6191 1390
rect 5427 1328 5433 1362
rect 5467 1328 5691 1362
rect 5725 1328 5949 1362
rect 5983 1352 6191 1362
rect 5983 1328 6132 1352
rect 5427 1318 6132 1328
rect 6166 1318 6191 1352
rect 315 1280 530 1290
rect 315 1246 340 1280
rect 374 1256 530 1280
rect 564 1256 788 1290
rect 822 1256 1046 1290
rect 1080 1256 1098 1290
rect 374 1246 1098 1256
rect 315 1208 1098 1246
rect 315 1174 340 1208
rect 374 1174 1098 1208
rect 5427 1290 6191 1318
rect 5427 1256 5433 1290
rect 5467 1256 5691 1290
rect 5725 1256 5949 1290
rect 5983 1280 6191 1290
rect 5983 1256 6132 1280
rect 5427 1246 6132 1256
rect 6166 1246 6191 1280
rect 5427 1208 6191 1246
rect 315 1162 1098 1174
rect 315 1136 623 1162
rect 315 1102 340 1136
rect 374 1128 623 1136
rect 657 1128 695 1162
rect 729 1128 881 1162
rect 915 1128 953 1162
rect 987 1128 1098 1162
rect 374 1102 1098 1128
rect 315 1064 1098 1102
rect 315 1030 340 1064
rect 374 1030 1098 1064
rect 1290 1111 1740 1183
rect 1290 1059 1421 1111
rect 1473 1059 1485 1111
rect 1537 1059 1549 1111
rect 1601 1059 1740 1111
rect 1290 1051 1740 1059
rect 1806 1111 2256 1183
rect 1806 1059 1937 1111
rect 1989 1059 2001 1111
rect 2053 1059 2065 1111
rect 2117 1059 2256 1111
rect 1806 1051 2256 1059
rect 2516 1111 2966 1183
rect 2516 1059 2647 1111
rect 2699 1059 2711 1111
rect 2763 1059 2775 1111
rect 2827 1059 2966 1111
rect 2516 1051 2966 1059
rect 3032 1111 3482 1183
rect 3032 1059 3163 1111
rect 3215 1059 3227 1111
rect 3279 1059 3291 1111
rect 3343 1059 3482 1111
rect 3032 1051 3482 1059
rect 3548 1111 3998 1183
rect 3548 1059 3679 1111
rect 3731 1059 3743 1111
rect 3795 1059 3807 1111
rect 3859 1059 3998 1111
rect 3548 1051 3998 1059
rect 4258 1111 4708 1183
rect 4258 1059 4389 1111
rect 4441 1059 4453 1111
rect 4505 1059 4517 1111
rect 4569 1059 4708 1111
rect 4258 1051 4708 1059
rect 4774 1111 5224 1183
rect 4774 1059 4905 1111
rect 4957 1059 4969 1111
rect 5021 1059 5033 1111
rect 5085 1059 5224 1111
rect 4774 1051 5224 1059
rect 5427 1174 6132 1208
rect 6166 1174 6191 1208
rect 5427 1162 6191 1174
rect 5427 1128 5526 1162
rect 5560 1128 5598 1162
rect 5632 1128 5784 1162
rect 5818 1128 5856 1162
rect 5890 1136 6191 1162
rect 5890 1128 6132 1136
rect 5427 1102 6132 1128
rect 6166 1102 6191 1136
rect 5427 1064 6191 1102
rect 315 992 1098 1030
rect 315 958 340 992
rect 374 958 1098 992
rect 5427 1030 6132 1064
rect 6166 1030 6191 1064
rect 5427 992 6191 1030
rect 315 920 1098 958
rect 315 886 340 920
rect 374 886 1098 920
rect 315 881 1098 886
rect 315 848 623 881
rect 315 814 340 848
rect 374 847 623 848
rect 657 847 695 881
rect 729 847 881 881
rect 915 847 953 881
rect 987 847 1098 881
rect 374 814 1098 847
rect 1290 963 1740 971
rect 1290 911 1421 963
rect 1473 911 1485 963
rect 1537 911 1549 963
rect 1601 911 1740 963
rect 1290 839 1740 911
rect 1806 963 2256 971
rect 1806 911 1937 963
rect 1989 911 2001 963
rect 2053 911 2065 963
rect 2117 911 2256 963
rect 1806 839 2256 911
rect 2516 963 2966 971
rect 2516 911 2647 963
rect 2699 911 2711 963
rect 2763 911 2775 963
rect 2827 911 2966 963
rect 2516 839 2966 911
rect 3032 963 3482 971
rect 3032 911 3163 963
rect 3215 911 3227 963
rect 3279 911 3291 963
rect 3343 911 3482 963
rect 3032 839 3482 911
rect 3548 963 3998 971
rect 3548 911 3679 963
rect 3731 911 3743 963
rect 3795 911 3807 963
rect 3859 911 3998 963
rect 3548 839 3998 911
rect 4258 963 4708 971
rect 4258 911 4389 963
rect 4441 911 4453 963
rect 4505 911 4517 963
rect 4569 911 4708 963
rect 4258 839 4708 911
rect 4774 963 5224 971
rect 4774 911 4905 963
rect 4957 911 4969 963
rect 5021 911 5033 963
rect 5085 911 5224 963
rect 4774 839 5224 911
rect 5427 958 6132 992
rect 6166 958 6191 992
rect 5427 920 6191 958
rect 5427 886 6132 920
rect 6166 886 6191 920
rect 5427 881 6191 886
rect 5427 847 5526 881
rect 5560 847 5598 881
rect 5632 847 5784 881
rect 5818 847 5856 881
rect 5890 848 6191 881
rect 5890 847 6132 848
rect 315 776 1098 814
rect 315 742 340 776
rect 374 753 1098 776
rect 374 742 530 753
rect 315 719 530 742
rect 564 719 788 753
rect 822 719 1046 753
rect 1080 719 1098 753
rect 5427 814 6132 847
rect 6166 814 6191 848
rect 5427 776 6191 814
rect 5427 753 6132 776
rect 315 704 1098 719
rect 315 670 340 704
rect 374 681 1098 704
rect 374 670 530 681
rect 315 647 530 670
rect 564 647 788 681
rect 822 647 1046 681
rect 1080 647 1098 681
rect 315 632 1098 647
rect 315 598 340 632
rect 374 598 1098 632
rect 315 570 1098 598
rect 1234 570 1280 740
rect 315 560 1280 570
rect 315 526 340 560
rect 374 526 1074 560
rect 315 508 1074 526
rect 1126 508 1138 560
rect 1190 508 1202 560
rect 1254 508 1280 560
rect 315 500 1280 508
rect 315 488 1098 500
rect 315 454 340 488
rect 374 454 1098 488
rect 315 416 1098 454
rect 315 382 340 416
rect 374 382 1098 416
rect 315 344 1098 382
rect 315 310 340 344
rect 374 310 1098 344
rect 315 272 1098 310
rect 315 238 340 272
rect 374 267 1098 272
rect 374 238 530 267
rect 315 233 530 238
rect 564 233 788 267
rect 822 233 1046 267
rect 1080 233 1098 267
rect 315 200 1098 233
rect 1234 226 1280 500
rect 1750 433 1796 736
rect 2266 570 2312 740
rect 2112 560 2312 570
rect 2112 508 2121 560
rect 2173 508 2185 560
rect 2237 508 2249 560
rect 2301 508 2312 560
rect 2112 500 2312 508
rect 1672 423 1868 433
rect 1672 371 1681 423
rect 1733 371 1745 423
rect 1797 371 1809 423
rect 1861 371 1868 423
rect 1672 363 1868 371
rect 1750 222 1796 363
rect 2266 226 2312 500
rect 2460 433 2506 740
rect 2976 570 3022 715
rect 2914 560 3110 570
rect 2914 508 2921 560
rect 2973 508 2985 560
rect 3037 508 3049 560
rect 3101 508 3110 560
rect 2914 500 3110 508
rect 2460 423 2665 433
rect 2460 371 2478 423
rect 2530 371 2542 423
rect 2594 371 2606 423
rect 2658 371 2665 423
rect 2460 363 2665 371
rect 2460 226 2506 363
rect 2976 202 3022 500
rect 3492 433 3538 715
rect 4008 570 4054 740
rect 4202 570 4248 740
rect 4008 560 4248 570
rect 4008 508 4034 560
rect 4086 508 4098 560
rect 4150 508 4162 560
rect 4214 508 4248 560
rect 4008 500 4248 508
rect 3417 423 3613 433
rect 3417 371 3424 423
rect 3476 371 3488 423
rect 3540 371 3552 423
rect 3604 371 3613 423
rect 3417 363 3613 371
rect 3492 202 3538 363
rect 4008 226 4054 500
rect 4202 226 4248 500
rect 4718 433 4764 736
rect 5234 570 5280 740
rect 5427 719 5433 753
rect 5467 719 5691 753
rect 5725 719 5949 753
rect 5983 742 6132 753
rect 6166 742 6191 776
rect 5983 719 6191 742
rect 5427 704 6191 719
rect 5427 681 6132 704
rect 5427 647 5433 681
rect 5467 647 5691 681
rect 5725 647 5949 681
rect 5983 670 6132 681
rect 6166 670 6191 704
rect 5983 647 6191 670
rect 5427 632 6191 647
rect 5427 598 6132 632
rect 6166 598 6191 632
rect 5427 570 6191 598
rect 5234 560 6191 570
rect 5234 508 5262 560
rect 5314 508 5326 560
rect 5378 508 5390 560
rect 5442 526 6132 560
rect 6166 526 6191 560
rect 5442 508 6191 526
rect 5234 500 6191 508
rect 4642 423 4838 433
rect 4642 371 4651 423
rect 4703 371 4715 423
rect 4767 371 4779 423
rect 4831 371 4838 423
rect 4642 363 4838 371
rect 4718 222 4764 363
rect 5234 226 5280 500
rect 5427 488 6191 500
rect 5427 454 6132 488
rect 6166 454 6191 488
rect 5427 416 6191 454
rect 5427 382 6132 416
rect 6166 382 6191 416
rect 5427 344 6191 382
rect 5427 310 6132 344
rect 6166 310 6191 344
rect 5427 272 6191 310
rect 5427 267 6132 272
rect 5427 233 5433 267
rect 5467 233 5691 267
rect 5725 233 5949 267
rect 5983 238 6132 267
rect 6166 238 6191 272
rect 5983 233 6191 238
rect 315 166 340 200
rect 374 195 1098 200
rect 374 166 530 195
rect 315 161 530 166
rect 564 161 788 195
rect 822 161 1046 195
rect 1080 161 1098 195
rect 315 128 1098 161
rect 315 94 340 128
rect 374 94 1098 128
rect 315 67 1098 94
rect 5427 200 6191 233
rect 5427 195 6132 200
rect 5427 161 5433 195
rect 5467 161 5691 195
rect 5725 161 5949 195
rect 5983 166 6132 195
rect 6166 166 6191 200
rect 5983 161 6191 166
rect 5427 128 6191 161
rect 5427 94 6132 128
rect 6166 94 6191 128
rect 315 56 623 67
rect 315 22 340 56
rect 374 33 623 56
rect 657 33 695 67
rect 729 33 881 67
rect 915 33 953 67
rect 987 33 1098 67
rect 374 22 1098 33
rect 315 -16 1098 22
rect 315 -50 340 -16
rect 374 -50 1098 -16
rect 1290 17 1740 89
rect 1290 -35 1421 17
rect 1473 -35 1485 17
rect 1537 -35 1549 17
rect 1601 -35 1740 17
rect 1290 -43 1740 -35
rect 1806 17 2256 89
rect 1806 -35 1937 17
rect 1989 -35 2001 17
rect 2053 -35 2065 17
rect 2117 -35 2256 17
rect 1806 -43 2256 -35
rect 2516 17 2966 89
rect 2516 -35 2647 17
rect 2699 -35 2711 17
rect 2763 -35 2775 17
rect 2827 -35 2966 17
rect 2516 -43 2966 -35
rect 3032 17 3482 89
rect 3032 -35 3163 17
rect 3215 -35 3227 17
rect 3279 -35 3291 17
rect 3343 -35 3482 17
rect 3032 -43 3482 -35
rect 3548 17 3998 89
rect 3548 -35 3679 17
rect 3731 -35 3743 17
rect 3795 -35 3807 17
rect 3859 -35 3998 17
rect 3548 -43 3998 -35
rect 4258 17 4708 89
rect 4258 -35 4389 17
rect 4441 -35 4453 17
rect 4505 -35 4517 17
rect 4569 -35 4708 17
rect 4258 -43 4708 -35
rect 4774 17 5224 89
rect 4774 -35 4905 17
rect 4957 -35 4969 17
rect 5021 -35 5033 17
rect 5085 -35 5224 17
rect 4774 -43 5224 -35
rect 5427 67 6191 94
rect 5427 33 5526 67
rect 5560 33 5598 67
rect 5632 33 5784 67
rect 5818 33 5856 67
rect 5890 56 6191 67
rect 5890 33 6132 56
rect 5427 22 6132 33
rect 6166 22 6191 56
rect 5427 -16 6191 22
rect 315 -88 1098 -50
rect 315 -122 340 -88
rect 374 -122 1098 -88
rect 315 -160 1098 -122
rect 5427 -50 6132 -16
rect 6166 -50 6191 -16
rect 5427 -88 6191 -50
rect 5427 -122 6132 -88
rect 6166 -122 6191 -88
rect 315 -194 340 -160
rect 374 -194 1098 -160
rect 315 -214 1098 -194
rect 315 -232 623 -214
rect 315 -266 340 -232
rect 374 -248 623 -232
rect 657 -248 695 -214
rect 729 -248 881 -214
rect 915 -248 953 -214
rect 987 -248 1098 -214
rect 374 -266 1098 -248
rect 1290 -132 1740 -124
rect 1290 -184 1421 -132
rect 1473 -184 1485 -132
rect 1537 -184 1549 -132
rect 1601 -184 1740 -132
rect 1290 -256 1740 -184
rect 1806 -132 2256 -124
rect 1806 -184 1937 -132
rect 1989 -184 2001 -132
rect 2053 -184 2065 -132
rect 2117 -184 2256 -132
rect 1806 -256 2256 -184
rect 2516 -132 2966 -124
rect 2516 -184 2647 -132
rect 2699 -184 2711 -132
rect 2763 -184 2775 -132
rect 2827 -184 2966 -132
rect 2516 -256 2966 -184
rect 3032 -132 3482 -124
rect 3032 -184 3163 -132
rect 3215 -184 3227 -132
rect 3279 -184 3291 -132
rect 3343 -184 3482 -132
rect 3032 -256 3482 -184
rect 3548 -132 3998 -124
rect 3548 -184 3679 -132
rect 3731 -184 3743 -132
rect 3795 -184 3807 -132
rect 3859 -184 3998 -132
rect 3548 -256 3998 -184
rect 4258 -132 4708 -124
rect 4258 -184 4389 -132
rect 4441 -184 4453 -132
rect 4505 -184 4517 -132
rect 4569 -184 4708 -132
rect 4258 -256 4708 -184
rect 4774 -132 5224 -124
rect 4774 -184 4905 -132
rect 4957 -184 4969 -132
rect 5021 -184 5033 -132
rect 5085 -184 5224 -132
rect 4774 -256 5224 -184
rect 5427 -160 6191 -122
rect 5427 -194 6132 -160
rect 6166 -194 6191 -160
rect 5427 -214 6191 -194
rect 5427 -248 5526 -214
rect 5560 -248 5598 -214
rect 5632 -248 5784 -214
rect 5818 -248 5856 -214
rect 5890 -232 6191 -214
rect 5890 -248 6132 -232
rect 315 -304 1098 -266
rect 315 -338 340 -304
rect 374 -338 1098 -304
rect 315 -342 1098 -338
rect 315 -376 530 -342
rect 564 -376 788 -342
rect 822 -376 1046 -342
rect 1080 -376 1098 -342
rect 5427 -266 6132 -248
rect 6166 -266 6191 -232
rect 5427 -304 6191 -266
rect 5427 -338 6132 -304
rect 6166 -338 6191 -304
rect 5427 -342 6191 -338
rect 315 -410 340 -376
rect 374 -410 1098 -376
rect 315 -414 1098 -410
rect 315 -448 530 -414
rect 564 -448 788 -414
rect 822 -448 1046 -414
rect 1080 -448 1098 -414
rect 315 -482 340 -448
rect 374 -482 1098 -448
rect 315 -520 1098 -482
rect 315 -554 340 -520
rect 374 -522 1098 -520
rect 1234 -522 1280 -355
rect 374 -532 1280 -522
rect 374 -554 1074 -532
rect 315 -584 1074 -554
rect 1126 -584 1138 -532
rect 1190 -584 1202 -532
rect 1254 -584 1280 -532
rect 315 -592 1280 -584
rect 315 -626 340 -592
rect 374 -626 1098 -592
rect 315 -664 1098 -626
rect 315 -698 340 -664
rect 374 -698 1098 -664
rect 315 -736 1098 -698
rect 315 -770 340 -736
rect 374 -770 1098 -736
rect 315 -808 1098 -770
rect 315 -842 340 -808
rect 374 -819 1098 -808
rect 374 -842 530 -819
rect 315 -853 530 -842
rect 564 -853 788 -819
rect 822 -853 1046 -819
rect 1080 -853 1098 -819
rect 315 -880 1098 -853
rect 1234 -869 1280 -592
rect 1750 -662 1796 -355
rect 2266 -523 2312 -355
rect 2110 -533 2312 -523
rect 2110 -585 2119 -533
rect 2171 -585 2183 -533
rect 2235 -585 2247 -533
rect 2299 -585 2312 -533
rect 2110 -593 2312 -585
rect 1672 -672 1868 -662
rect 1672 -724 1681 -672
rect 1733 -724 1745 -672
rect 1797 -724 1809 -672
rect 1861 -724 1868 -672
rect 1672 -732 1868 -724
rect 1750 -869 1796 -732
rect 2266 -869 2312 -593
rect 2460 -662 2506 -355
rect 2976 -523 3022 -376
rect 2914 -533 3110 -523
rect 2914 -585 2921 -533
rect 2973 -585 2985 -533
rect 3037 -585 3049 -533
rect 3101 -585 3110 -533
rect 2914 -593 3110 -585
rect 2460 -672 2665 -662
rect 2460 -724 2478 -672
rect 2530 -724 2542 -672
rect 2594 -724 2606 -672
rect 2658 -724 2665 -672
rect 2460 -732 2665 -724
rect 2460 -869 2506 -732
rect 315 -914 340 -880
rect 374 -891 1098 -880
rect 2976 -889 3022 -593
rect 3492 -662 3538 -376
rect 4008 -523 4054 -355
rect 4202 -523 4248 -355
rect 4008 -533 4248 -523
rect 4008 -585 4034 -533
rect 4086 -585 4098 -533
rect 4150 -585 4162 -533
rect 4214 -585 4248 -533
rect 4008 -593 4248 -585
rect 3417 -672 3613 -662
rect 3417 -724 3424 -672
rect 3476 -724 3488 -672
rect 3540 -724 3552 -672
rect 3604 -724 3613 -672
rect 3417 -732 3613 -724
rect 3492 -889 3538 -732
rect 4008 -869 4054 -593
rect 4202 -869 4248 -593
rect 4718 -662 4764 -355
rect 5234 -523 5280 -355
rect 5427 -376 5433 -342
rect 5467 -376 5691 -342
rect 5725 -376 5949 -342
rect 5983 -376 6191 -342
rect 5427 -410 6132 -376
rect 6166 -410 6191 -376
rect 5427 -414 6191 -410
rect 5427 -448 5433 -414
rect 5467 -448 5691 -414
rect 5725 -448 5949 -414
rect 5983 -448 6191 -414
rect 5427 -482 6132 -448
rect 6166 -482 6191 -448
rect 5427 -520 6191 -482
rect 5427 -523 6132 -520
rect 5234 -533 6132 -523
rect 5234 -585 5262 -533
rect 5314 -585 5326 -533
rect 5378 -585 5390 -533
rect 5442 -554 6132 -533
rect 6166 -554 6191 -520
rect 5442 -585 6191 -554
rect 5234 -592 6191 -585
rect 5234 -593 6132 -592
rect 4642 -672 4838 -662
rect 4642 -724 4651 -672
rect 4703 -724 4715 -672
rect 4767 -724 4779 -672
rect 4831 -724 4838 -672
rect 4642 -732 4838 -724
rect 4718 -869 4764 -732
rect 5234 -869 5280 -593
rect 5427 -626 6132 -593
rect 6166 -626 6191 -592
rect 5427 -664 6191 -626
rect 5427 -698 6132 -664
rect 6166 -698 6191 -664
rect 5427 -736 6191 -698
rect 5427 -770 6132 -736
rect 6166 -770 6191 -736
rect 5427 -808 6191 -770
rect 5427 -819 6132 -808
rect 5427 -853 5433 -819
rect 5467 -853 5691 -819
rect 5725 -853 5949 -819
rect 5983 -842 6132 -819
rect 6166 -842 6191 -808
rect 5983 -853 6191 -842
rect 5427 -880 6191 -853
rect 374 -914 530 -891
rect 315 -925 530 -914
rect 564 -925 788 -891
rect 822 -925 1046 -891
rect 1080 -925 1098 -891
rect 315 -952 1098 -925
rect 315 -986 340 -952
rect 374 -986 1098 -952
rect 315 -1019 1098 -986
rect 5427 -891 6132 -880
rect 5427 -925 5433 -891
rect 5467 -925 5691 -891
rect 5725 -925 5949 -891
rect 5983 -914 6132 -891
rect 6166 -914 6191 -880
rect 5983 -925 6191 -914
rect 5427 -952 6191 -925
rect 5427 -986 6132 -952
rect 6166 -986 6191 -952
rect 315 -1024 623 -1019
rect 315 -1058 340 -1024
rect 374 -1053 623 -1024
rect 657 -1053 695 -1019
rect 729 -1053 881 -1019
rect 915 -1053 953 -1019
rect 987 -1053 1098 -1019
rect 374 -1058 1098 -1053
rect 315 -1096 1098 -1058
rect 315 -1130 340 -1096
rect 374 -1130 1098 -1096
rect 315 -1168 1098 -1130
rect 1290 -1075 1740 -1003
rect 1290 -1127 1421 -1075
rect 1473 -1127 1485 -1075
rect 1537 -1127 1549 -1075
rect 1601 -1127 1740 -1075
rect 1290 -1135 1740 -1127
rect 1806 -1075 2256 -1003
rect 1806 -1127 1937 -1075
rect 1989 -1127 2001 -1075
rect 2053 -1127 2065 -1075
rect 2117 -1127 2256 -1075
rect 1806 -1135 2256 -1127
rect 2516 -1075 2966 -1003
rect 2516 -1127 2647 -1075
rect 2699 -1127 2711 -1075
rect 2763 -1127 2775 -1075
rect 2827 -1127 2966 -1075
rect 2516 -1135 2966 -1127
rect 3032 -1075 3482 -1003
rect 3032 -1127 3163 -1075
rect 3215 -1127 3227 -1075
rect 3279 -1127 3291 -1075
rect 3343 -1127 3482 -1075
rect 3032 -1135 3482 -1127
rect 3548 -1075 3998 -1003
rect 3548 -1127 3679 -1075
rect 3731 -1127 3743 -1075
rect 3795 -1127 3807 -1075
rect 3859 -1127 3998 -1075
rect 3548 -1135 3998 -1127
rect 4258 -1075 4708 -1003
rect 4258 -1127 4389 -1075
rect 4441 -1127 4453 -1075
rect 4505 -1127 4517 -1075
rect 4569 -1127 4708 -1075
rect 4258 -1135 4708 -1127
rect 4774 -1075 5224 -1003
rect 4774 -1127 4905 -1075
rect 4957 -1127 4969 -1075
rect 5021 -1127 5033 -1075
rect 5085 -1127 5224 -1075
rect 4774 -1135 5224 -1127
rect 5427 -1019 6191 -986
rect 5427 -1053 5526 -1019
rect 5560 -1053 5598 -1019
rect 5632 -1053 5784 -1019
rect 5818 -1053 5856 -1019
rect 5890 -1024 6191 -1019
rect 5890 -1053 6132 -1024
rect 5427 -1058 6132 -1053
rect 6166 -1058 6191 -1024
rect 5427 -1096 6191 -1058
rect 5427 -1130 6132 -1096
rect 6166 -1130 6191 -1096
rect 315 -1202 340 -1168
rect 374 -1202 1098 -1168
rect 315 -1240 1098 -1202
rect 5427 -1168 6191 -1130
rect 5427 -1202 6132 -1168
rect 6166 -1202 6191 -1168
rect 315 -1274 340 -1240
rect 374 -1274 1098 -1240
rect 315 -1300 1098 -1274
rect 315 -1312 623 -1300
rect 315 -1346 340 -1312
rect 374 -1334 623 -1312
rect 657 -1334 695 -1300
rect 729 -1334 881 -1300
rect 915 -1334 953 -1300
rect 987 -1334 1098 -1300
rect 374 -1346 1098 -1334
rect 1290 -1213 1740 -1205
rect 1290 -1265 1421 -1213
rect 1473 -1265 1485 -1213
rect 1537 -1265 1549 -1213
rect 1601 -1265 1740 -1213
rect 1290 -1337 1740 -1265
rect 1806 -1213 2256 -1205
rect 1806 -1265 1937 -1213
rect 1989 -1265 2001 -1213
rect 2053 -1265 2065 -1213
rect 2117 -1265 2256 -1213
rect 1806 -1337 2256 -1265
rect 2516 -1213 2966 -1205
rect 2516 -1265 2647 -1213
rect 2699 -1265 2711 -1213
rect 2763 -1265 2775 -1213
rect 2827 -1265 2966 -1213
rect 2516 -1337 2966 -1265
rect 3032 -1213 3482 -1205
rect 3032 -1265 3163 -1213
rect 3215 -1265 3227 -1213
rect 3279 -1265 3291 -1213
rect 3343 -1265 3482 -1213
rect 3032 -1337 3482 -1265
rect 3548 -1213 3998 -1205
rect 3548 -1265 3679 -1213
rect 3731 -1265 3743 -1213
rect 3795 -1265 3807 -1213
rect 3859 -1265 3998 -1213
rect 3548 -1337 3998 -1265
rect 4258 -1213 4708 -1205
rect 4258 -1265 4389 -1213
rect 4441 -1265 4453 -1213
rect 4505 -1265 4517 -1213
rect 4569 -1265 4708 -1213
rect 4258 -1337 4708 -1265
rect 4774 -1213 5224 -1205
rect 4774 -1265 4905 -1213
rect 4957 -1265 4969 -1213
rect 5021 -1265 5033 -1213
rect 5085 -1265 5224 -1213
rect 4774 -1337 5224 -1265
rect 5427 -1240 6191 -1202
rect 5427 -1274 6132 -1240
rect 6166 -1274 6191 -1240
rect 5427 -1300 6191 -1274
rect 5427 -1334 5526 -1300
rect 5560 -1334 5598 -1300
rect 5632 -1334 5784 -1300
rect 5818 -1334 5856 -1300
rect 5890 -1312 6191 -1300
rect 5890 -1334 6132 -1312
rect 315 -1384 1098 -1346
rect 315 -1418 340 -1384
rect 374 -1418 1098 -1384
rect 315 -1428 1098 -1418
rect 315 -1456 530 -1428
rect 315 -1490 340 -1456
rect 374 -1462 530 -1456
rect 564 -1462 788 -1428
rect 822 -1462 1046 -1428
rect 1080 -1462 1098 -1428
rect 374 -1490 1098 -1462
rect 5427 -1346 6132 -1334
rect 6166 -1346 6191 -1312
rect 5427 -1384 6191 -1346
rect 5427 -1418 6132 -1384
rect 6166 -1418 6191 -1384
rect 5427 -1428 6191 -1418
rect 5427 -1462 5433 -1428
rect 5467 -1462 5691 -1428
rect 5725 -1462 5949 -1428
rect 5983 -1456 6191 -1428
rect 5983 -1462 6132 -1456
rect 315 -1500 1098 -1490
rect 315 -1528 530 -1500
rect 315 -1562 340 -1528
rect 374 -1534 530 -1528
rect 564 -1534 788 -1500
rect 822 -1534 1046 -1500
rect 1080 -1534 1098 -1500
rect 374 -1562 1098 -1534
rect 315 -1600 1098 -1562
rect 315 -1634 340 -1600
rect 374 -1634 1098 -1600
rect 315 -1672 1098 -1634
rect 315 -1706 340 -1672
rect 374 -1706 1098 -1672
rect 315 -1744 1098 -1706
rect 315 -1778 340 -1744
rect 374 -1778 1098 -1744
rect 315 -1816 1098 -1778
rect 315 -1850 340 -1816
rect 374 -1850 1098 -1816
rect 315 -1888 1098 -1850
rect 315 -1922 340 -1888
rect 374 -1889 1098 -1888
rect 1234 -1889 1280 -1571
rect 1750 -1610 1796 -1480
rect 1672 -1618 1868 -1610
rect 1672 -1670 1681 -1618
rect 1733 -1670 1745 -1618
rect 1797 -1670 1809 -1618
rect 1861 -1670 1868 -1618
rect 1672 -1680 1868 -1670
rect 2266 -1889 2312 -1571
rect 2460 -1750 2506 -1480
rect 2460 -1758 2656 -1750
rect 2460 -1810 2469 -1758
rect 2521 -1810 2533 -1758
rect 2585 -1810 2597 -1758
rect 2649 -1810 2656 -1758
rect 2460 -1820 2656 -1810
rect 2976 -1889 3022 -1571
rect 3492 -1750 3538 -1480
rect 3417 -1758 3613 -1750
rect 3417 -1810 3424 -1758
rect 3476 -1810 3488 -1758
rect 3540 -1810 3552 -1758
rect 3604 -1810 3613 -1758
rect 3417 -1820 3613 -1810
rect 4008 -1889 4054 -1571
rect 4202 -1889 4248 -1571
rect 4718 -1610 4764 -1480
rect 5427 -1490 6132 -1462
rect 6166 -1490 6191 -1456
rect 5427 -1500 6191 -1490
rect 5427 -1534 5433 -1500
rect 5467 -1534 5691 -1500
rect 5725 -1534 5949 -1500
rect 5983 -1528 6191 -1500
rect 5983 -1534 6132 -1528
rect 5427 -1562 6132 -1534
rect 6166 -1562 6191 -1528
rect 4642 -1618 4838 -1610
rect 4642 -1670 4651 -1618
rect 4703 -1670 4715 -1618
rect 4767 -1670 4779 -1618
rect 4831 -1670 4838 -1618
rect 4642 -1680 4838 -1670
rect 374 -1899 1280 -1889
rect 374 -1922 1074 -1899
rect 315 -1951 1074 -1922
rect 1126 -1951 1138 -1899
rect 1190 -1951 1202 -1899
rect 1254 -1951 1280 -1899
rect 315 -1959 1280 -1951
rect 2108 -1899 2312 -1889
rect 2108 -1951 2117 -1899
rect 2169 -1951 2181 -1899
rect 2233 -1951 2245 -1899
rect 2297 -1951 2312 -1899
rect 2108 -1959 2312 -1951
rect 2914 -1899 3110 -1889
rect 2914 -1951 2921 -1899
rect 2973 -1951 2985 -1899
rect 3037 -1951 3049 -1899
rect 3101 -1951 3110 -1899
rect 2914 -1959 3110 -1951
rect 4008 -1899 4248 -1889
rect 4008 -1951 4034 -1899
rect 4086 -1951 4098 -1899
rect 4150 -1951 4162 -1899
rect 4214 -1951 4248 -1899
rect 4008 -1959 4248 -1951
rect 315 -1960 1098 -1959
rect 315 -1994 340 -1960
rect 374 -1994 1098 -1960
rect 315 -2032 1098 -1994
rect 315 -2066 340 -2032
rect 374 -2066 1098 -2032
rect 315 -2104 1098 -2066
rect 315 -2138 340 -2104
rect 374 -2138 1098 -2104
rect 315 -2176 1098 -2138
rect 315 -2210 340 -2176
rect 374 -2210 1098 -2176
rect 315 -2248 1098 -2210
rect 315 -2282 340 -2248
rect 374 -2282 1098 -2248
rect 315 -2320 1098 -2282
rect 315 -2354 340 -2320
rect 374 -2323 1098 -2320
rect 374 -2354 530 -2323
rect 315 -2357 530 -2354
rect 564 -2357 788 -2323
rect 822 -2357 1046 -2323
rect 1080 -2357 1098 -2323
rect 315 -2392 1098 -2357
rect 315 -2426 340 -2392
rect 374 -2395 1098 -2392
rect 374 -2426 530 -2395
rect 315 -2429 530 -2426
rect 564 -2429 788 -2395
rect 822 -2429 1046 -2395
rect 1080 -2429 1098 -2395
rect 1234 -2397 1280 -1959
rect 1672 -2178 1868 -2168
rect 1672 -2230 1681 -2178
rect 1733 -2230 1745 -2178
rect 1797 -2230 1809 -2178
rect 1861 -2230 1868 -2178
rect 1672 -2238 1868 -2230
rect 1750 -2368 1796 -2238
rect 2266 -2397 2312 -1959
rect 2460 -2037 2656 -2029
rect 2460 -2089 2469 -2037
rect 2521 -2089 2533 -2037
rect 2585 -2089 2597 -2037
rect 2649 -2089 2656 -2037
rect 2460 -2099 2656 -2089
rect 2460 -2368 2506 -2099
rect 2976 -2397 3022 -1959
rect 3417 -2037 3613 -2029
rect 3417 -2089 3424 -2037
rect 3476 -2089 3488 -2037
rect 3540 -2089 3552 -2037
rect 3604 -2089 3613 -2037
rect 3417 -2099 3613 -2089
rect 3492 -2368 3538 -2099
rect 4008 -2396 4054 -1959
rect 4202 -2396 4248 -1959
rect 5234 -1889 5280 -1571
rect 5427 -1600 6191 -1562
rect 5427 -1634 6132 -1600
rect 6166 -1634 6191 -1600
rect 5427 -1672 6191 -1634
rect 5427 -1706 6132 -1672
rect 6166 -1706 6191 -1672
rect 5427 -1744 6191 -1706
rect 5427 -1778 6132 -1744
rect 6166 -1778 6191 -1744
rect 5427 -1816 6191 -1778
rect 5427 -1850 6132 -1816
rect 6166 -1850 6191 -1816
rect 5427 -1888 6191 -1850
rect 5427 -1889 6132 -1888
rect 5234 -1899 6132 -1889
rect 5234 -1951 5262 -1899
rect 5314 -1951 5326 -1899
rect 5378 -1951 5390 -1899
rect 5442 -1922 6132 -1899
rect 6166 -1922 6191 -1888
rect 5442 -1951 6191 -1922
rect 5234 -1959 6191 -1951
rect 4642 -2178 4838 -2168
rect 4642 -2230 4651 -2178
rect 4703 -2230 4715 -2178
rect 4767 -2230 4779 -2178
rect 4831 -2230 4838 -2178
rect 4642 -2238 4838 -2230
rect 4718 -2368 4764 -2238
rect 5234 -2396 5280 -1959
rect 5427 -1960 6191 -1959
rect 5427 -1994 6132 -1960
rect 6166 -1994 6191 -1960
rect 5427 -2032 6191 -1994
rect 5427 -2066 6132 -2032
rect 6166 -2066 6191 -2032
rect 5427 -2104 6191 -2066
rect 5427 -2138 6132 -2104
rect 6166 -2138 6191 -2104
rect 5427 -2176 6191 -2138
rect 5427 -2210 6132 -2176
rect 6166 -2210 6191 -2176
rect 5427 -2248 6191 -2210
rect 5427 -2282 6132 -2248
rect 6166 -2282 6191 -2248
rect 5427 -2320 6191 -2282
rect 5427 -2323 6132 -2320
rect 5427 -2357 5433 -2323
rect 5467 -2357 5691 -2323
rect 5725 -2357 5949 -2323
rect 5983 -2354 6132 -2323
rect 6166 -2354 6191 -2320
rect 5983 -2357 6191 -2354
rect 5427 -2392 6191 -2357
rect 5427 -2395 6132 -2392
rect 315 -2464 1098 -2429
rect 315 -2498 340 -2464
rect 374 -2498 1098 -2464
rect 315 -2523 1098 -2498
rect 5427 -2429 5433 -2395
rect 5467 -2429 5691 -2395
rect 5725 -2429 5949 -2395
rect 5983 -2426 6132 -2395
rect 6166 -2426 6191 -2392
rect 5983 -2429 6191 -2426
rect 5427 -2464 6191 -2429
rect 5427 -2498 6132 -2464
rect 6166 -2498 6191 -2464
rect 315 -2536 623 -2523
rect 315 -2570 340 -2536
rect 374 -2557 623 -2536
rect 657 -2557 695 -2523
rect 729 -2557 881 -2523
rect 915 -2557 953 -2523
rect 987 -2557 1098 -2523
rect 374 -2570 1098 -2557
rect 315 -2608 1098 -2570
rect 315 -2642 340 -2608
rect 374 -2642 1098 -2608
rect 1290 -2579 1740 -2507
rect 1290 -2631 1421 -2579
rect 1473 -2631 1485 -2579
rect 1537 -2631 1549 -2579
rect 1601 -2631 1740 -2579
rect 1290 -2639 1740 -2631
rect 1806 -2579 2256 -2507
rect 1806 -2631 1937 -2579
rect 1989 -2631 2001 -2579
rect 2053 -2631 2065 -2579
rect 2117 -2631 2256 -2579
rect 1806 -2639 2256 -2631
rect 2516 -2579 2966 -2507
rect 2516 -2631 2647 -2579
rect 2699 -2631 2711 -2579
rect 2763 -2631 2775 -2579
rect 2827 -2631 2966 -2579
rect 2516 -2639 2966 -2631
rect 3032 -2579 3482 -2507
rect 3032 -2631 3163 -2579
rect 3215 -2631 3227 -2579
rect 3279 -2631 3291 -2579
rect 3343 -2631 3482 -2579
rect 3032 -2639 3482 -2631
rect 3548 -2579 3998 -2507
rect 3548 -2631 3679 -2579
rect 3731 -2631 3743 -2579
rect 3795 -2631 3807 -2579
rect 3859 -2631 3998 -2579
rect 3548 -2639 3998 -2631
rect 4258 -2579 4708 -2507
rect 4258 -2631 4389 -2579
rect 4441 -2631 4453 -2579
rect 4505 -2631 4517 -2579
rect 4569 -2631 4708 -2579
rect 4258 -2639 4708 -2631
rect 4774 -2579 5224 -2507
rect 4774 -2631 4905 -2579
rect 4957 -2631 4969 -2579
rect 5021 -2631 5033 -2579
rect 5085 -2631 5224 -2579
rect 4774 -2639 5224 -2631
rect 5427 -2523 6191 -2498
rect 5427 -2557 5526 -2523
rect 5560 -2557 5598 -2523
rect 5632 -2557 5784 -2523
rect 5818 -2557 5856 -2523
rect 5890 -2536 6191 -2523
rect 5890 -2557 6132 -2536
rect 5427 -2570 6132 -2557
rect 6166 -2570 6191 -2536
rect 5427 -2608 6191 -2570
rect 315 -2680 1098 -2642
rect 315 -2714 340 -2680
rect 374 -2714 1098 -2680
rect 5427 -2642 6132 -2608
rect 6166 -2642 6191 -2608
rect 5427 -2680 6191 -2642
rect 315 -2752 1098 -2714
rect 315 -2786 340 -2752
rect 374 -2786 1098 -2752
rect 315 -2804 1098 -2786
rect 315 -2824 623 -2804
rect 315 -2858 340 -2824
rect 374 -2838 623 -2824
rect 657 -2838 695 -2804
rect 729 -2838 881 -2804
rect 915 -2838 953 -2804
rect 987 -2838 1098 -2804
rect 374 -2858 1098 -2838
rect 1290 -2717 1740 -2709
rect 1290 -2769 1421 -2717
rect 1473 -2769 1485 -2717
rect 1537 -2769 1549 -2717
rect 1601 -2769 1740 -2717
rect 1290 -2841 1740 -2769
rect 1806 -2717 2256 -2709
rect 1806 -2769 1937 -2717
rect 1989 -2769 2001 -2717
rect 2053 -2769 2065 -2717
rect 2117 -2769 2256 -2717
rect 1806 -2841 2256 -2769
rect 2516 -2717 2966 -2709
rect 2516 -2769 2647 -2717
rect 2699 -2769 2711 -2717
rect 2763 -2769 2775 -2717
rect 2827 -2769 2966 -2717
rect 2516 -2841 2966 -2769
rect 3032 -2717 3482 -2709
rect 3032 -2769 3163 -2717
rect 3215 -2769 3227 -2717
rect 3279 -2769 3291 -2717
rect 3343 -2769 3482 -2717
rect 3032 -2841 3482 -2769
rect 3548 -2717 3998 -2709
rect 3548 -2769 3679 -2717
rect 3731 -2769 3743 -2717
rect 3795 -2769 3807 -2717
rect 3859 -2769 3998 -2717
rect 3548 -2841 3998 -2769
rect 4258 -2717 4708 -2709
rect 4258 -2769 4389 -2717
rect 4441 -2769 4453 -2717
rect 4505 -2769 4517 -2717
rect 4569 -2769 4708 -2717
rect 4258 -2841 4708 -2769
rect 4774 -2717 5224 -2709
rect 4774 -2769 4905 -2717
rect 4957 -2769 4969 -2717
rect 5021 -2769 5033 -2717
rect 5085 -2769 5224 -2717
rect 4774 -2841 5224 -2769
rect 5427 -2714 6132 -2680
rect 6166 -2714 6191 -2680
rect 5427 -2752 6191 -2714
rect 5427 -2786 6132 -2752
rect 6166 -2786 6191 -2752
rect 5427 -2804 6191 -2786
rect 5427 -2838 5526 -2804
rect 5560 -2838 5598 -2804
rect 5632 -2838 5784 -2804
rect 5818 -2838 5856 -2804
rect 5890 -2824 6191 -2804
rect 5890 -2838 6132 -2824
rect 315 -2896 1098 -2858
rect 315 -2930 340 -2896
rect 374 -2930 1098 -2896
rect 315 -2932 1098 -2930
rect 315 -2966 530 -2932
rect 564 -2966 788 -2932
rect 822 -2966 1046 -2932
rect 1080 -2966 1098 -2932
rect 315 -2968 1098 -2966
rect 315 -3002 340 -2968
rect 374 -3002 1098 -2968
rect 5427 -2858 6132 -2838
rect 6166 -2858 6191 -2824
rect 5427 -2896 6191 -2858
rect 5427 -2930 6132 -2896
rect 6166 -2930 6191 -2896
rect 5427 -2932 6191 -2930
rect 5427 -2966 5433 -2932
rect 5467 -2966 5691 -2932
rect 5725 -2966 5949 -2932
rect 5983 -2966 6191 -2932
rect 5427 -2968 6191 -2966
rect 315 -3004 1098 -3002
rect 315 -3038 530 -3004
rect 564 -3038 788 -3004
rect 822 -3038 1046 -3004
rect 1080 -3038 1098 -3004
rect 315 -3040 1098 -3038
rect 315 -3074 340 -3040
rect 374 -3074 1098 -3040
rect 315 -3112 1098 -3074
rect 315 -3146 340 -3112
rect 374 -3146 1098 -3112
rect 315 -3184 1098 -3146
rect 315 -3218 340 -3184
rect 374 -3218 1098 -3184
rect 315 -3256 1098 -3218
rect 315 -3290 340 -3256
rect 374 -3290 1098 -3256
rect 315 -3328 1098 -3290
rect 315 -3362 340 -3328
rect 374 -3362 1098 -3328
rect 315 -3393 1098 -3362
rect 1234 -3393 1280 -3075
rect 1750 -3114 1796 -2984
rect 1672 -3122 1868 -3114
rect 1672 -3174 1681 -3122
rect 1733 -3174 1745 -3122
rect 1797 -3174 1809 -3122
rect 1861 -3174 1868 -3122
rect 1672 -3184 1868 -3174
rect 2266 -3393 2312 -3075
rect 2460 -3254 2506 -2984
rect 2460 -3262 2656 -3254
rect 2460 -3314 2469 -3262
rect 2521 -3314 2533 -3262
rect 2585 -3314 2597 -3262
rect 2649 -3314 2656 -3262
rect 2460 -3324 2656 -3314
rect 2976 -3393 3022 -3075
rect 3492 -3254 3538 -2984
rect 3417 -3262 3613 -3254
rect 3417 -3314 3424 -3262
rect 3476 -3314 3488 -3262
rect 3540 -3314 3552 -3262
rect 3604 -3314 3613 -3262
rect 3417 -3324 3613 -3314
rect 4008 -3393 4054 -3075
rect 4202 -3393 4248 -3075
rect 4718 -3114 4764 -2984
rect 5427 -3002 6132 -2968
rect 6166 -3002 6191 -2968
rect 5427 -3004 6191 -3002
rect 5427 -3038 5433 -3004
rect 5467 -3038 5691 -3004
rect 5725 -3038 5949 -3004
rect 5983 -3038 6191 -3004
rect 5427 -3040 6191 -3038
rect 5427 -3074 6132 -3040
rect 6166 -3074 6191 -3040
rect 4642 -3122 4838 -3114
rect 4642 -3174 4651 -3122
rect 4703 -3174 4715 -3122
rect 4767 -3174 4779 -3122
rect 4831 -3174 4838 -3122
rect 4642 -3184 4838 -3174
rect 315 -3400 1280 -3393
rect 315 -3434 340 -3400
rect 374 -3403 1280 -3400
rect 374 -3434 1074 -3403
rect 315 -3455 1074 -3434
rect 1126 -3455 1138 -3403
rect 1190 -3455 1202 -3403
rect 1254 -3455 1280 -3403
rect 315 -3463 1280 -3455
rect 2108 -3403 2312 -3393
rect 2108 -3455 2117 -3403
rect 2169 -3455 2181 -3403
rect 2233 -3455 2245 -3403
rect 2297 -3455 2312 -3403
rect 2108 -3463 2312 -3455
rect 2914 -3403 3110 -3393
rect 2914 -3455 2921 -3403
rect 2973 -3455 2985 -3403
rect 3037 -3455 3049 -3403
rect 3101 -3455 3110 -3403
rect 2914 -3463 3110 -3455
rect 4008 -3403 4248 -3393
rect 4008 -3455 4034 -3403
rect 4086 -3455 4098 -3403
rect 4150 -3455 4162 -3403
rect 4214 -3455 4248 -3403
rect 4008 -3463 4248 -3455
rect 315 -3472 1098 -3463
rect 315 -3506 340 -3472
rect 374 -3506 1098 -3472
rect 315 -3544 1098 -3506
rect 315 -3578 340 -3544
rect 374 -3578 1098 -3544
rect 315 -3616 1098 -3578
rect 315 -3650 340 -3616
rect 374 -3650 1098 -3616
rect 315 -3688 1098 -3650
rect 315 -3722 340 -3688
rect 374 -3722 1098 -3688
rect 315 -3760 1098 -3722
rect 315 -3794 340 -3760
rect 374 -3794 1098 -3760
rect 315 -3827 1098 -3794
rect 315 -3832 530 -3827
rect 315 -3866 340 -3832
rect 374 -3861 530 -3832
rect 564 -3861 788 -3827
rect 822 -3861 1046 -3827
rect 1080 -3861 1098 -3827
rect 374 -3866 1098 -3861
rect 315 -3899 1098 -3866
rect 315 -3904 530 -3899
rect 315 -3938 340 -3904
rect 374 -3933 530 -3904
rect 564 -3933 788 -3899
rect 822 -3933 1046 -3899
rect 1080 -3933 1098 -3899
rect 1234 -3901 1280 -3463
rect 1672 -3682 1868 -3672
rect 1672 -3734 1681 -3682
rect 1733 -3734 1745 -3682
rect 1797 -3734 1809 -3682
rect 1861 -3734 1868 -3682
rect 1672 -3742 1868 -3734
rect 1750 -3872 1796 -3742
rect 2266 -3901 2312 -3463
rect 2460 -3541 2656 -3533
rect 2460 -3593 2469 -3541
rect 2521 -3593 2533 -3541
rect 2585 -3593 2597 -3541
rect 2649 -3593 2656 -3541
rect 2460 -3603 2656 -3593
rect 2460 -3872 2506 -3603
rect 2976 -3901 3022 -3463
rect 3417 -3541 3613 -3533
rect 3417 -3593 3424 -3541
rect 3476 -3593 3488 -3541
rect 3540 -3593 3552 -3541
rect 3604 -3593 3613 -3541
rect 3417 -3603 3613 -3593
rect 3492 -3872 3538 -3603
rect 4008 -3900 4054 -3463
rect 4202 -3900 4248 -3463
rect 5234 -3393 5280 -3075
rect 5427 -3112 6191 -3074
rect 5427 -3146 6132 -3112
rect 6166 -3146 6191 -3112
rect 5427 -3184 6191 -3146
rect 5427 -3218 6132 -3184
rect 6166 -3218 6191 -3184
rect 5427 -3256 6191 -3218
rect 5427 -3290 6132 -3256
rect 6166 -3290 6191 -3256
rect 5427 -3328 6191 -3290
rect 5427 -3362 6132 -3328
rect 6166 -3362 6191 -3328
rect 5427 -3393 6191 -3362
rect 5234 -3400 6191 -3393
rect 5234 -3403 6132 -3400
rect 5234 -3455 5262 -3403
rect 5314 -3455 5326 -3403
rect 5378 -3455 5390 -3403
rect 5442 -3434 6132 -3403
rect 6166 -3434 6191 -3400
rect 5442 -3455 6191 -3434
rect 5234 -3463 6191 -3455
rect 4642 -3682 4838 -3672
rect 4642 -3734 4651 -3682
rect 4703 -3734 4715 -3682
rect 4767 -3734 4779 -3682
rect 4831 -3734 4838 -3682
rect 4642 -3742 4838 -3734
rect 4718 -3872 4764 -3742
rect 5234 -3900 5280 -3463
rect 5427 -3472 6191 -3463
rect 5427 -3506 6132 -3472
rect 6166 -3506 6191 -3472
rect 5427 -3544 6191 -3506
rect 5427 -3578 6132 -3544
rect 6166 -3578 6191 -3544
rect 5427 -3616 6191 -3578
rect 5427 -3650 6132 -3616
rect 6166 -3650 6191 -3616
rect 5427 -3688 6191 -3650
rect 5427 -3722 6132 -3688
rect 6166 -3722 6191 -3688
rect 5427 -3760 6191 -3722
rect 5427 -3794 6132 -3760
rect 6166 -3794 6191 -3760
rect 5427 -3827 6191 -3794
rect 5427 -3861 5433 -3827
rect 5467 -3861 5691 -3827
rect 5725 -3861 5949 -3827
rect 5983 -3832 6191 -3827
rect 5983 -3861 6132 -3832
rect 5427 -3866 6132 -3861
rect 6166 -3866 6191 -3832
rect 5427 -3899 6191 -3866
rect 374 -3938 1098 -3933
rect 315 -3976 1098 -3938
rect 315 -4010 340 -3976
rect 374 -4010 1098 -3976
rect 315 -4027 1098 -4010
rect 5427 -3933 5433 -3899
rect 5467 -3933 5691 -3899
rect 5725 -3933 5949 -3899
rect 5983 -3904 6191 -3899
rect 5983 -3933 6132 -3904
rect 5427 -3938 6132 -3933
rect 6166 -3938 6191 -3904
rect 5427 -3976 6191 -3938
rect 5427 -4010 6132 -3976
rect 6166 -4010 6191 -3976
rect 315 -4048 623 -4027
rect 315 -4082 340 -4048
rect 374 -4061 623 -4048
rect 657 -4061 695 -4027
rect 729 -4061 881 -4027
rect 915 -4061 953 -4027
rect 987 -4061 1098 -4027
rect 374 -4082 1098 -4061
rect 315 -4120 1098 -4082
rect 315 -4154 340 -4120
rect 374 -4154 1098 -4120
rect 1290 -4083 1740 -4011
rect 1290 -4135 1421 -4083
rect 1473 -4135 1485 -4083
rect 1537 -4135 1549 -4083
rect 1601 -4135 1740 -4083
rect 1290 -4143 1740 -4135
rect 1806 -4083 2256 -4011
rect 1806 -4135 1937 -4083
rect 1989 -4135 2001 -4083
rect 2053 -4135 2065 -4083
rect 2117 -4135 2256 -4083
rect 1806 -4143 2256 -4135
rect 2516 -4083 2966 -4011
rect 2516 -4135 2647 -4083
rect 2699 -4135 2711 -4083
rect 2763 -4135 2775 -4083
rect 2827 -4135 2966 -4083
rect 2516 -4143 2966 -4135
rect 3032 -4083 3482 -4011
rect 3032 -4135 3163 -4083
rect 3215 -4135 3227 -4083
rect 3279 -4135 3291 -4083
rect 3343 -4135 3482 -4083
rect 3032 -4143 3482 -4135
rect 3548 -4083 3998 -4011
rect 3548 -4135 3679 -4083
rect 3731 -4135 3743 -4083
rect 3795 -4135 3807 -4083
rect 3859 -4135 3998 -4083
rect 3548 -4143 3998 -4135
rect 4258 -4083 4708 -4011
rect 4258 -4135 4389 -4083
rect 4441 -4135 4453 -4083
rect 4505 -4135 4517 -4083
rect 4569 -4135 4708 -4083
rect 4258 -4143 4708 -4135
rect 4774 -4083 5224 -4011
rect 4774 -4135 4905 -4083
rect 4957 -4135 4969 -4083
rect 5021 -4135 5033 -4083
rect 5085 -4135 5224 -4083
rect 4774 -4143 5224 -4135
rect 5427 -4027 6191 -4010
rect 5427 -4061 5526 -4027
rect 5560 -4061 5598 -4027
rect 5632 -4061 5784 -4027
rect 5818 -4061 5856 -4027
rect 5890 -4048 6191 -4027
rect 5890 -4061 6132 -4048
rect 5427 -4082 6132 -4061
rect 6166 -4082 6191 -4048
rect 5427 -4120 6191 -4082
rect 315 -4192 1098 -4154
rect 315 -4226 340 -4192
rect 374 -4226 1098 -4192
rect 5427 -4154 6132 -4120
rect 6166 -4154 6191 -4120
rect 5427 -4192 6191 -4154
rect 315 -4264 1098 -4226
rect 315 -4298 340 -4264
rect 374 -4298 1098 -4264
rect 315 -4308 1098 -4298
rect 315 -4336 623 -4308
rect 315 -4370 340 -4336
rect 374 -4342 623 -4336
rect 657 -4342 695 -4308
rect 729 -4342 881 -4308
rect 915 -4342 953 -4308
rect 987 -4342 1098 -4308
rect 374 -4370 1098 -4342
rect 1290 -4221 1740 -4213
rect 1290 -4273 1421 -4221
rect 1473 -4273 1485 -4221
rect 1537 -4273 1549 -4221
rect 1601 -4273 1740 -4221
rect 1290 -4345 1740 -4273
rect 1806 -4221 2256 -4213
rect 1806 -4273 1937 -4221
rect 1989 -4273 2001 -4221
rect 2053 -4273 2065 -4221
rect 2117 -4273 2256 -4221
rect 1806 -4345 2256 -4273
rect 2516 -4221 2966 -4213
rect 2516 -4273 2647 -4221
rect 2699 -4273 2711 -4221
rect 2763 -4273 2775 -4221
rect 2827 -4273 2966 -4221
rect 2516 -4345 2966 -4273
rect 3032 -4221 3482 -4213
rect 3032 -4273 3163 -4221
rect 3215 -4273 3227 -4221
rect 3279 -4273 3291 -4221
rect 3343 -4273 3482 -4221
rect 3032 -4345 3482 -4273
rect 3548 -4221 3998 -4213
rect 3548 -4273 3679 -4221
rect 3731 -4273 3743 -4221
rect 3795 -4273 3807 -4221
rect 3859 -4273 3998 -4221
rect 3548 -4345 3998 -4273
rect 4258 -4221 4708 -4213
rect 4258 -4273 4389 -4221
rect 4441 -4273 4453 -4221
rect 4505 -4273 4517 -4221
rect 4569 -4273 4708 -4221
rect 4258 -4345 4708 -4273
rect 4774 -4221 5224 -4213
rect 4774 -4273 4905 -4221
rect 4957 -4273 4969 -4221
rect 5021 -4273 5033 -4221
rect 5085 -4273 5224 -4221
rect 4774 -4345 5224 -4273
rect 5427 -4226 6132 -4192
rect 6166 -4226 6191 -4192
rect 5427 -4264 6191 -4226
rect 5427 -4298 6132 -4264
rect 6166 -4298 6191 -4264
rect 5427 -4308 6191 -4298
rect 5427 -4342 5526 -4308
rect 5560 -4342 5598 -4308
rect 5632 -4342 5784 -4308
rect 5818 -4342 5856 -4308
rect 5890 -4336 6191 -4308
rect 5890 -4342 6132 -4336
rect 315 -4408 1098 -4370
rect 315 -4442 340 -4408
rect 374 -4436 1098 -4408
rect 374 -4442 530 -4436
rect 315 -4470 530 -4442
rect 564 -4470 788 -4436
rect 822 -4470 1046 -4436
rect 1080 -4470 1098 -4436
rect 315 -4480 1098 -4470
rect 315 -4514 340 -4480
rect 374 -4508 1098 -4480
rect 5427 -4370 6132 -4342
rect 6166 -4370 6191 -4336
rect 5427 -4408 6191 -4370
rect 5427 -4436 6132 -4408
rect 5427 -4470 5433 -4436
rect 5467 -4470 5691 -4436
rect 5725 -4470 5949 -4436
rect 5983 -4442 6132 -4436
rect 6166 -4442 6191 -4408
rect 5983 -4470 6191 -4442
rect 5427 -4480 6191 -4470
rect 374 -4514 530 -4508
rect 315 -4542 530 -4514
rect 564 -4542 788 -4508
rect 822 -4542 1046 -4508
rect 1080 -4542 1098 -4508
rect 315 -4552 1098 -4542
rect 315 -4586 340 -4552
rect 374 -4586 1098 -4552
rect 315 -4624 1098 -4586
rect 315 -4658 340 -4624
rect 374 -4658 1098 -4624
rect 315 -4696 1098 -4658
rect 315 -4730 340 -4696
rect 374 -4730 1098 -4696
rect 315 -4768 1098 -4730
rect 315 -4802 340 -4768
rect 374 -4802 1098 -4768
rect 315 -4840 1098 -4802
rect 315 -4874 340 -4840
rect 374 -4874 1098 -4840
rect 315 -4897 1098 -4874
rect 1234 -4897 1280 -4579
rect 1750 -4618 1796 -4488
rect 1672 -4626 1868 -4618
rect 1672 -4678 1681 -4626
rect 1733 -4678 1745 -4626
rect 1797 -4678 1809 -4626
rect 1861 -4678 1868 -4626
rect 1672 -4688 1868 -4678
rect 2266 -4897 2312 -4579
rect 2460 -4758 2506 -4488
rect 2460 -4766 2656 -4758
rect 2460 -4818 2469 -4766
rect 2521 -4818 2533 -4766
rect 2585 -4818 2597 -4766
rect 2649 -4818 2656 -4766
rect 2460 -4828 2656 -4818
rect 2976 -4897 3022 -4579
rect 3492 -4758 3538 -4488
rect 3417 -4766 3613 -4758
rect 3417 -4818 3424 -4766
rect 3476 -4818 3488 -4766
rect 3540 -4818 3552 -4766
rect 3604 -4818 3613 -4766
rect 3417 -4828 3613 -4818
rect 4008 -4897 4054 -4579
rect 4202 -4897 4248 -4579
rect 4718 -4618 4764 -4488
rect 5427 -4508 6132 -4480
rect 5427 -4542 5433 -4508
rect 5467 -4542 5691 -4508
rect 5725 -4542 5949 -4508
rect 5983 -4514 6132 -4508
rect 6166 -4514 6191 -4480
rect 5983 -4542 6191 -4514
rect 5427 -4552 6191 -4542
rect 4642 -4626 4838 -4618
rect 4642 -4678 4651 -4626
rect 4703 -4678 4715 -4626
rect 4767 -4678 4779 -4626
rect 4831 -4678 4838 -4626
rect 4642 -4688 4838 -4678
rect 5234 -4897 5280 -4579
rect 5427 -4586 6132 -4552
rect 6166 -4586 6191 -4552
rect 5427 -4624 6191 -4586
rect 5427 -4658 6132 -4624
rect 6166 -4658 6191 -4624
rect 5427 -4696 6191 -4658
rect 5427 -4730 6132 -4696
rect 6166 -4730 6191 -4696
rect 5427 -4768 6191 -4730
rect 5427 -4802 6132 -4768
rect 6166 -4802 6191 -4768
rect 5427 -4840 6191 -4802
rect 5427 -4874 6132 -4840
rect 6166 -4874 6191 -4840
rect 5427 -4897 6191 -4874
rect 315 -4907 6191 -4897
rect 315 -4912 1074 -4907
rect 315 -4946 340 -4912
rect 374 -4946 1074 -4912
rect 315 -4959 1074 -4946
rect 1126 -4959 1138 -4907
rect 1190 -4959 1202 -4907
rect 1254 -4959 2117 -4907
rect 2169 -4959 2181 -4907
rect 2233 -4959 2245 -4907
rect 2297 -4959 2921 -4907
rect 2973 -4959 2985 -4907
rect 3037 -4959 3049 -4907
rect 3101 -4959 4034 -4907
rect 4086 -4959 4098 -4907
rect 4150 -4959 4162 -4907
rect 4214 -4959 5262 -4907
rect 5314 -4959 5326 -4907
rect 5378 -4959 5390 -4907
rect 5442 -4912 6191 -4907
rect 5442 -4946 6132 -4912
rect 6166 -4946 6191 -4912
rect 5442 -4959 6191 -4946
rect 315 -4984 6191 -4959
rect 315 -5018 340 -4984
rect 374 -5018 6132 -4984
rect 6166 -5018 6191 -4984
rect 315 -5056 6191 -5018
rect 315 -5090 340 -5056
rect 374 -5090 6132 -5056
rect 6166 -5090 6191 -5056
rect 315 -5128 6191 -5090
rect 315 -5162 340 -5128
rect 374 -5162 6132 -5128
rect 6166 -5162 6191 -5128
rect 315 -5183 6191 -5162
rect 315 -5200 530 -5183
rect 315 -5234 340 -5200
rect 374 -5217 530 -5200
rect 564 -5217 788 -5183
rect 822 -5217 1046 -5183
rect 1080 -5217 1240 -5183
rect 1274 -5217 1498 -5183
rect 1532 -5217 1756 -5183
rect 1790 -5217 2014 -5183
rect 2048 -5217 2272 -5183
rect 2306 -5217 2466 -5183
rect 2500 -5217 2724 -5183
rect 2758 -5217 2982 -5183
rect 3016 -5217 3240 -5183
rect 3274 -5217 3498 -5183
rect 3532 -5217 3756 -5183
rect 3790 -5217 4014 -5183
rect 4048 -5217 4208 -5183
rect 4242 -5217 4466 -5183
rect 4500 -5217 4724 -5183
rect 4758 -5217 4982 -5183
rect 5016 -5217 5240 -5183
rect 5274 -5217 5433 -5183
rect 5467 -5217 5691 -5183
rect 5725 -5217 5949 -5183
rect 5983 -5200 6191 -5183
rect 5983 -5217 6132 -5200
rect 374 -5234 6132 -5217
rect 6166 -5234 6191 -5200
rect 315 -5255 6191 -5234
rect 315 -5272 530 -5255
rect 315 -5306 340 -5272
rect 374 -5289 530 -5272
rect 564 -5289 788 -5255
rect 822 -5289 1046 -5255
rect 1080 -5289 1240 -5255
rect 1274 -5289 1498 -5255
rect 1532 -5289 1756 -5255
rect 1790 -5289 2014 -5255
rect 2048 -5289 2272 -5255
rect 2306 -5289 2466 -5255
rect 2500 -5289 2724 -5255
rect 2758 -5289 2982 -5255
rect 3016 -5289 3240 -5255
rect 3274 -5289 3498 -5255
rect 3532 -5289 3756 -5255
rect 3790 -5289 4014 -5255
rect 4048 -5289 4208 -5255
rect 4242 -5289 4466 -5255
rect 4500 -5289 4724 -5255
rect 4758 -5289 4982 -5255
rect 5016 -5289 5240 -5255
rect 5274 -5289 5433 -5255
rect 5467 -5289 5691 -5255
rect 5725 -5289 5949 -5255
rect 5983 -5272 6191 -5255
rect 5983 -5289 6132 -5272
rect 374 -5306 6132 -5289
rect 6166 -5306 6191 -5272
rect 315 -5344 6191 -5306
rect 315 -5378 340 -5344
rect 374 -5378 6132 -5344
rect 6166 -5378 6191 -5344
rect 315 -5383 6191 -5378
rect 315 -5417 623 -5383
rect 657 -5417 695 -5383
rect 729 -5417 881 -5383
rect 915 -5417 953 -5383
rect 987 -5417 1333 -5383
rect 1367 -5417 1405 -5383
rect 1439 -5417 1591 -5383
rect 1625 -5417 1663 -5383
rect 1697 -5417 1849 -5383
rect 1883 -5417 1921 -5383
rect 1955 -5417 2107 -5383
rect 2141 -5417 2179 -5383
rect 2213 -5417 2559 -5383
rect 2593 -5417 2631 -5383
rect 2665 -5417 2817 -5383
rect 2851 -5417 2889 -5383
rect 2923 -5417 3075 -5383
rect 3109 -5417 3147 -5383
rect 3181 -5417 3333 -5383
rect 3367 -5417 3405 -5383
rect 3439 -5417 3591 -5383
rect 3625 -5417 3663 -5383
rect 3697 -5417 3849 -5383
rect 3883 -5417 3921 -5383
rect 3955 -5417 4301 -5383
rect 4335 -5417 4373 -5383
rect 4407 -5417 4559 -5383
rect 4593 -5417 4631 -5383
rect 4665 -5417 4817 -5383
rect 4851 -5417 4889 -5383
rect 4923 -5417 5075 -5383
rect 5109 -5417 5147 -5383
rect 5181 -5417 5526 -5383
rect 5560 -5417 5598 -5383
rect 5632 -5417 5784 -5383
rect 5818 -5417 5856 -5383
rect 5890 -5417 6191 -5383
rect 315 -5506 6191 -5417
rect 315 -5540 487 -5506
rect 521 -5540 559 -5506
rect 593 -5540 631 -5506
rect 665 -5540 703 -5506
rect 737 -5540 775 -5506
rect 809 -5540 847 -5506
rect 881 -5540 919 -5506
rect 953 -5540 991 -5506
rect 1025 -5540 1063 -5506
rect 1097 -5540 1135 -5506
rect 1169 -5540 1207 -5506
rect 1241 -5540 1279 -5506
rect 1313 -5540 1351 -5506
rect 1385 -5540 1423 -5506
rect 1457 -5540 1495 -5506
rect 1529 -5540 1567 -5506
rect 1601 -5540 1639 -5506
rect 1673 -5540 1711 -5506
rect 1745 -5540 1783 -5506
rect 1817 -5540 1855 -5506
rect 1889 -5540 1927 -5506
rect 1961 -5540 1999 -5506
rect 2033 -5540 2071 -5506
rect 2105 -5540 2143 -5506
rect 2177 -5540 2215 -5506
rect 2249 -5540 2287 -5506
rect 2321 -5540 2359 -5506
rect 2393 -5540 2431 -5506
rect 2465 -5540 2503 -5506
rect 2537 -5540 2575 -5506
rect 2609 -5540 2647 -5506
rect 2681 -5540 2719 -5506
rect 2753 -5540 2791 -5506
rect 2825 -5540 2863 -5506
rect 2897 -5540 2935 -5506
rect 2969 -5540 3007 -5506
rect 3041 -5540 3079 -5506
rect 3113 -5540 3151 -5506
rect 3185 -5540 3223 -5506
rect 3257 -5540 3295 -5506
rect 3329 -5540 3367 -5506
rect 3401 -5540 3439 -5506
rect 3473 -5540 3511 -5506
rect 3545 -5540 3583 -5506
rect 3617 -5540 3655 -5506
rect 3689 -5540 3727 -5506
rect 3761 -5540 3799 -5506
rect 3833 -5540 3871 -5506
rect 3905 -5540 3943 -5506
rect 3977 -5540 4015 -5506
rect 4049 -5540 4087 -5506
rect 4121 -5540 4159 -5506
rect 4193 -5540 4231 -5506
rect 4265 -5540 4303 -5506
rect 4337 -5540 4375 -5506
rect 4409 -5540 4447 -5506
rect 4481 -5540 4519 -5506
rect 4553 -5540 4591 -5506
rect 4625 -5540 4663 -5506
rect 4697 -5540 4735 -5506
rect 4769 -5540 4807 -5506
rect 4841 -5540 4879 -5506
rect 4913 -5540 4951 -5506
rect 4985 -5540 5023 -5506
rect 5057 -5540 5095 -5506
rect 5129 -5540 5167 -5506
rect 5201 -5540 5239 -5506
rect 5273 -5540 5311 -5506
rect 5345 -5540 5383 -5506
rect 5417 -5540 5455 -5506
rect 5489 -5540 5527 -5506
rect 5561 -5540 5599 -5506
rect 5633 -5540 5671 -5506
rect 5705 -5540 5743 -5506
rect 5777 -5540 5815 -5506
rect 5849 -5540 5887 -5506
rect 5921 -5540 5959 -5506
rect 5993 -5540 6191 -5506
rect 315 -5565 6191 -5540
<< via1 >>
rect 1421 5296 1473 5348
rect 1485 5296 1537 5348
rect 1549 5296 1601 5348
rect 1937 5296 1989 5348
rect 2001 5296 2053 5348
rect 2065 5296 2117 5348
rect 2647 5296 2699 5348
rect 2711 5296 2763 5348
rect 2775 5296 2827 5348
rect 3163 5296 3215 5348
rect 3227 5296 3279 5348
rect 3291 5296 3343 5348
rect 3679 5296 3731 5348
rect 3743 5296 3795 5348
rect 3807 5296 3859 5348
rect 4389 5296 4441 5348
rect 4453 5296 4505 5348
rect 4517 5296 4569 5348
rect 4905 5296 4957 5348
rect 4969 5296 5021 5348
rect 5033 5296 5085 5348
rect 1681 4891 1733 4943
rect 1745 4891 1797 4943
rect 1809 4891 1861 4943
rect 2469 4751 2521 4803
rect 2533 4751 2585 4803
rect 2597 4751 2649 4803
rect 3424 4751 3476 4803
rect 3488 4751 3540 4803
rect 3552 4751 3604 4803
rect 4651 4891 4703 4943
rect 4715 4891 4767 4943
rect 4779 4891 4831 4943
rect 1074 4610 1126 4662
rect 1138 4610 1190 4662
rect 1202 4610 1254 4662
rect 2117 4610 2169 4662
rect 2181 4610 2233 4662
rect 2245 4610 2297 4662
rect 2921 4610 2973 4662
rect 2985 4610 3037 4662
rect 3049 4610 3101 4662
rect 4034 4610 4086 4662
rect 4098 4610 4150 4662
rect 4162 4610 4214 4662
rect 1681 4331 1733 4383
rect 1745 4331 1797 4383
rect 1809 4331 1861 4383
rect 2469 4472 2521 4524
rect 2533 4472 2585 4524
rect 2597 4472 2649 4524
rect 3424 4472 3476 4524
rect 3488 4472 3540 4524
rect 3552 4472 3604 4524
rect 5262 4610 5314 4662
rect 5326 4610 5378 4662
rect 5390 4610 5442 4662
rect 4651 4331 4703 4383
rect 4715 4331 4767 4383
rect 4779 4331 4831 4383
rect 1421 3930 1473 3982
rect 1485 3930 1537 3982
rect 1549 3930 1601 3982
rect 1937 3930 1989 3982
rect 2001 3930 2053 3982
rect 2065 3930 2117 3982
rect 2647 3930 2699 3982
rect 2711 3930 2763 3982
rect 2775 3930 2827 3982
rect 3163 3930 3215 3982
rect 3227 3930 3279 3982
rect 3291 3930 3343 3982
rect 3679 3930 3731 3982
rect 3743 3930 3795 3982
rect 3807 3930 3859 3982
rect 4389 3930 4441 3982
rect 4453 3930 4505 3982
rect 4517 3930 4569 3982
rect 4905 3930 4957 3982
rect 4969 3930 5021 3982
rect 5033 3930 5085 3982
rect 1421 3792 1473 3844
rect 1485 3792 1537 3844
rect 1549 3792 1601 3844
rect 1937 3792 1989 3844
rect 2001 3792 2053 3844
rect 2065 3792 2117 3844
rect 2647 3792 2699 3844
rect 2711 3792 2763 3844
rect 2775 3792 2827 3844
rect 3163 3792 3215 3844
rect 3227 3792 3279 3844
rect 3291 3792 3343 3844
rect 3679 3792 3731 3844
rect 3743 3792 3795 3844
rect 3807 3792 3859 3844
rect 4389 3792 4441 3844
rect 4453 3792 4505 3844
rect 4517 3792 4569 3844
rect 4905 3792 4957 3844
rect 4969 3792 5021 3844
rect 5033 3792 5085 3844
rect 1681 3387 1733 3439
rect 1745 3387 1797 3439
rect 1809 3387 1861 3439
rect 2469 3247 2521 3299
rect 2533 3247 2585 3299
rect 2597 3247 2649 3299
rect 3424 3247 3476 3299
rect 3488 3247 3540 3299
rect 3552 3247 3604 3299
rect 4651 3387 4703 3439
rect 4715 3387 4767 3439
rect 4779 3387 4831 3439
rect 1074 3106 1126 3158
rect 1138 3106 1190 3158
rect 1202 3106 1254 3158
rect 2117 3106 2169 3158
rect 2181 3106 2233 3158
rect 2245 3106 2297 3158
rect 2921 3106 2973 3158
rect 2985 3106 3037 3158
rect 3049 3106 3101 3158
rect 4034 3106 4086 3158
rect 4098 3106 4150 3158
rect 4162 3106 4214 3158
rect 1681 2827 1733 2879
rect 1745 2827 1797 2879
rect 1809 2827 1861 2879
rect 2469 2968 2521 3020
rect 2533 2968 2585 3020
rect 2597 2968 2649 3020
rect 3424 2968 3476 3020
rect 3488 2968 3540 3020
rect 3552 2968 3604 3020
rect 5262 3106 5314 3158
rect 5326 3106 5378 3158
rect 5390 3106 5442 3158
rect 4651 2827 4703 2879
rect 4715 2827 4767 2879
rect 4779 2827 4831 2879
rect 1421 2426 1473 2478
rect 1485 2426 1537 2478
rect 1549 2426 1601 2478
rect 1937 2426 1989 2478
rect 2001 2426 2053 2478
rect 2065 2426 2117 2478
rect 2647 2426 2699 2478
rect 2711 2426 2763 2478
rect 2775 2426 2827 2478
rect 3163 2426 3215 2478
rect 3227 2426 3279 2478
rect 3291 2426 3343 2478
rect 3679 2426 3731 2478
rect 3743 2426 3795 2478
rect 3807 2426 3859 2478
rect 4389 2426 4441 2478
rect 4453 2426 4505 2478
rect 4517 2426 4569 2478
rect 4905 2426 4957 2478
rect 4969 2426 5021 2478
rect 5033 2426 5085 2478
rect 1421 2278 1473 2330
rect 1485 2278 1537 2330
rect 1549 2278 1601 2330
rect 1937 2278 1989 2330
rect 2001 2278 2053 2330
rect 2065 2278 2117 2330
rect 2647 2278 2699 2330
rect 2711 2278 2763 2330
rect 2775 2278 2827 2330
rect 3163 2278 3215 2330
rect 3227 2278 3279 2330
rect 3291 2278 3343 2330
rect 3679 2278 3731 2330
rect 3743 2278 3795 2330
rect 3807 2278 3859 2330
rect 4389 2278 4441 2330
rect 4453 2278 4505 2330
rect 4517 2278 4569 2330
rect 4905 2278 4957 2330
rect 4969 2278 5021 2330
rect 5033 2278 5085 2330
rect 1681 1879 1733 1931
rect 1745 1879 1797 1931
rect 1809 1879 1861 1931
rect 2469 1739 2521 1791
rect 2533 1739 2585 1791
rect 2597 1739 2649 1791
rect 3424 1739 3476 1791
rect 3488 1739 3540 1791
rect 3552 1739 3604 1791
rect 4651 1879 4703 1931
rect 4715 1879 4767 1931
rect 4779 1879 4831 1931
rect 1074 1598 1126 1650
rect 1138 1598 1190 1650
rect 1202 1598 1254 1650
rect 2117 1598 2169 1650
rect 2181 1598 2233 1650
rect 2245 1598 2297 1650
rect 2921 1598 2973 1650
rect 2985 1598 3037 1650
rect 3049 1598 3101 1650
rect 4034 1598 4086 1650
rect 4098 1598 4150 1650
rect 4162 1598 4214 1650
rect 1681 1458 1733 1510
rect 1745 1458 1797 1510
rect 1809 1458 1861 1510
rect 2478 1458 2530 1510
rect 2542 1458 2594 1510
rect 2606 1458 2658 1510
rect 3424 1458 3476 1510
rect 3488 1458 3540 1510
rect 3552 1458 3604 1510
rect 5262 1598 5314 1650
rect 5326 1598 5378 1650
rect 5390 1598 5442 1650
rect 4651 1458 4703 1510
rect 4715 1458 4767 1510
rect 4779 1458 4831 1510
rect 1421 1059 1473 1111
rect 1485 1059 1537 1111
rect 1549 1059 1601 1111
rect 1937 1059 1989 1111
rect 2001 1059 2053 1111
rect 2065 1059 2117 1111
rect 2647 1059 2699 1111
rect 2711 1059 2763 1111
rect 2775 1059 2827 1111
rect 3163 1059 3215 1111
rect 3227 1059 3279 1111
rect 3291 1059 3343 1111
rect 3679 1059 3731 1111
rect 3743 1059 3795 1111
rect 3807 1059 3859 1111
rect 4389 1059 4441 1111
rect 4453 1059 4505 1111
rect 4517 1059 4569 1111
rect 4905 1059 4957 1111
rect 4969 1059 5021 1111
rect 5033 1059 5085 1111
rect 1421 911 1473 963
rect 1485 911 1537 963
rect 1549 911 1601 963
rect 1937 911 1989 963
rect 2001 911 2053 963
rect 2065 911 2117 963
rect 2647 911 2699 963
rect 2711 911 2763 963
rect 2775 911 2827 963
rect 3163 911 3215 963
rect 3227 911 3279 963
rect 3291 911 3343 963
rect 3679 911 3731 963
rect 3743 911 3795 963
rect 3807 911 3859 963
rect 4389 911 4441 963
rect 4453 911 4505 963
rect 4517 911 4569 963
rect 4905 911 4957 963
rect 4969 911 5021 963
rect 5033 911 5085 963
rect 1074 508 1126 560
rect 1138 508 1190 560
rect 1202 508 1254 560
rect 2121 508 2173 560
rect 2185 508 2237 560
rect 2249 508 2301 560
rect 1681 371 1733 423
rect 1745 371 1797 423
rect 1809 371 1861 423
rect 2921 508 2973 560
rect 2985 508 3037 560
rect 3049 508 3101 560
rect 2478 371 2530 423
rect 2542 371 2594 423
rect 2606 371 2658 423
rect 4034 508 4086 560
rect 4098 508 4150 560
rect 4162 508 4214 560
rect 3424 371 3476 423
rect 3488 371 3540 423
rect 3552 371 3604 423
rect 5262 508 5314 560
rect 5326 508 5378 560
rect 5390 508 5442 560
rect 4651 371 4703 423
rect 4715 371 4767 423
rect 4779 371 4831 423
rect 1421 -35 1473 17
rect 1485 -35 1537 17
rect 1549 -35 1601 17
rect 1937 -35 1989 17
rect 2001 -35 2053 17
rect 2065 -35 2117 17
rect 2647 -35 2699 17
rect 2711 -35 2763 17
rect 2775 -35 2827 17
rect 3163 -35 3215 17
rect 3227 -35 3279 17
rect 3291 -35 3343 17
rect 3679 -35 3731 17
rect 3743 -35 3795 17
rect 3807 -35 3859 17
rect 4389 -35 4441 17
rect 4453 -35 4505 17
rect 4517 -35 4569 17
rect 4905 -35 4957 17
rect 4969 -35 5021 17
rect 5033 -35 5085 17
rect 1421 -184 1473 -132
rect 1485 -184 1537 -132
rect 1549 -184 1601 -132
rect 1937 -184 1989 -132
rect 2001 -184 2053 -132
rect 2065 -184 2117 -132
rect 2647 -184 2699 -132
rect 2711 -184 2763 -132
rect 2775 -184 2827 -132
rect 3163 -184 3215 -132
rect 3227 -184 3279 -132
rect 3291 -184 3343 -132
rect 3679 -184 3731 -132
rect 3743 -184 3795 -132
rect 3807 -184 3859 -132
rect 4389 -184 4441 -132
rect 4453 -184 4505 -132
rect 4517 -184 4569 -132
rect 4905 -184 4957 -132
rect 4969 -184 5021 -132
rect 5033 -184 5085 -132
rect 1074 -584 1126 -532
rect 1138 -584 1190 -532
rect 1202 -584 1254 -532
rect 2119 -585 2171 -533
rect 2183 -585 2235 -533
rect 2247 -585 2299 -533
rect 1681 -724 1733 -672
rect 1745 -724 1797 -672
rect 1809 -724 1861 -672
rect 2921 -585 2973 -533
rect 2985 -585 3037 -533
rect 3049 -585 3101 -533
rect 2478 -724 2530 -672
rect 2542 -724 2594 -672
rect 2606 -724 2658 -672
rect 4034 -585 4086 -533
rect 4098 -585 4150 -533
rect 4162 -585 4214 -533
rect 3424 -724 3476 -672
rect 3488 -724 3540 -672
rect 3552 -724 3604 -672
rect 5262 -585 5314 -533
rect 5326 -585 5378 -533
rect 5390 -585 5442 -533
rect 4651 -724 4703 -672
rect 4715 -724 4767 -672
rect 4779 -724 4831 -672
rect 1421 -1127 1473 -1075
rect 1485 -1127 1537 -1075
rect 1549 -1127 1601 -1075
rect 1937 -1127 1989 -1075
rect 2001 -1127 2053 -1075
rect 2065 -1127 2117 -1075
rect 2647 -1127 2699 -1075
rect 2711 -1127 2763 -1075
rect 2775 -1127 2827 -1075
rect 3163 -1127 3215 -1075
rect 3227 -1127 3279 -1075
rect 3291 -1127 3343 -1075
rect 3679 -1127 3731 -1075
rect 3743 -1127 3795 -1075
rect 3807 -1127 3859 -1075
rect 4389 -1127 4441 -1075
rect 4453 -1127 4505 -1075
rect 4517 -1127 4569 -1075
rect 4905 -1127 4957 -1075
rect 4969 -1127 5021 -1075
rect 5033 -1127 5085 -1075
rect 1421 -1265 1473 -1213
rect 1485 -1265 1537 -1213
rect 1549 -1265 1601 -1213
rect 1937 -1265 1989 -1213
rect 2001 -1265 2053 -1213
rect 2065 -1265 2117 -1213
rect 2647 -1265 2699 -1213
rect 2711 -1265 2763 -1213
rect 2775 -1265 2827 -1213
rect 3163 -1265 3215 -1213
rect 3227 -1265 3279 -1213
rect 3291 -1265 3343 -1213
rect 3679 -1265 3731 -1213
rect 3743 -1265 3795 -1213
rect 3807 -1265 3859 -1213
rect 4389 -1265 4441 -1213
rect 4453 -1265 4505 -1213
rect 4517 -1265 4569 -1213
rect 4905 -1265 4957 -1213
rect 4969 -1265 5021 -1213
rect 5033 -1265 5085 -1213
rect 1681 -1670 1733 -1618
rect 1745 -1670 1797 -1618
rect 1809 -1670 1861 -1618
rect 2469 -1810 2521 -1758
rect 2533 -1810 2585 -1758
rect 2597 -1810 2649 -1758
rect 3424 -1810 3476 -1758
rect 3488 -1810 3540 -1758
rect 3552 -1810 3604 -1758
rect 4651 -1670 4703 -1618
rect 4715 -1670 4767 -1618
rect 4779 -1670 4831 -1618
rect 1074 -1951 1126 -1899
rect 1138 -1951 1190 -1899
rect 1202 -1951 1254 -1899
rect 2117 -1951 2169 -1899
rect 2181 -1951 2233 -1899
rect 2245 -1951 2297 -1899
rect 2921 -1951 2973 -1899
rect 2985 -1951 3037 -1899
rect 3049 -1951 3101 -1899
rect 4034 -1951 4086 -1899
rect 4098 -1951 4150 -1899
rect 4162 -1951 4214 -1899
rect 1681 -2230 1733 -2178
rect 1745 -2230 1797 -2178
rect 1809 -2230 1861 -2178
rect 2469 -2089 2521 -2037
rect 2533 -2089 2585 -2037
rect 2597 -2089 2649 -2037
rect 3424 -2089 3476 -2037
rect 3488 -2089 3540 -2037
rect 3552 -2089 3604 -2037
rect 5262 -1951 5314 -1899
rect 5326 -1951 5378 -1899
rect 5390 -1951 5442 -1899
rect 4651 -2230 4703 -2178
rect 4715 -2230 4767 -2178
rect 4779 -2230 4831 -2178
rect 1421 -2631 1473 -2579
rect 1485 -2631 1537 -2579
rect 1549 -2631 1601 -2579
rect 1937 -2631 1989 -2579
rect 2001 -2631 2053 -2579
rect 2065 -2631 2117 -2579
rect 2647 -2631 2699 -2579
rect 2711 -2631 2763 -2579
rect 2775 -2631 2827 -2579
rect 3163 -2631 3215 -2579
rect 3227 -2631 3279 -2579
rect 3291 -2631 3343 -2579
rect 3679 -2631 3731 -2579
rect 3743 -2631 3795 -2579
rect 3807 -2631 3859 -2579
rect 4389 -2631 4441 -2579
rect 4453 -2631 4505 -2579
rect 4517 -2631 4569 -2579
rect 4905 -2631 4957 -2579
rect 4969 -2631 5021 -2579
rect 5033 -2631 5085 -2579
rect 1421 -2769 1473 -2717
rect 1485 -2769 1537 -2717
rect 1549 -2769 1601 -2717
rect 1937 -2769 1989 -2717
rect 2001 -2769 2053 -2717
rect 2065 -2769 2117 -2717
rect 2647 -2769 2699 -2717
rect 2711 -2769 2763 -2717
rect 2775 -2769 2827 -2717
rect 3163 -2769 3215 -2717
rect 3227 -2769 3279 -2717
rect 3291 -2769 3343 -2717
rect 3679 -2769 3731 -2717
rect 3743 -2769 3795 -2717
rect 3807 -2769 3859 -2717
rect 4389 -2769 4441 -2717
rect 4453 -2769 4505 -2717
rect 4517 -2769 4569 -2717
rect 4905 -2769 4957 -2717
rect 4969 -2769 5021 -2717
rect 5033 -2769 5085 -2717
rect 1681 -3174 1733 -3122
rect 1745 -3174 1797 -3122
rect 1809 -3174 1861 -3122
rect 2469 -3314 2521 -3262
rect 2533 -3314 2585 -3262
rect 2597 -3314 2649 -3262
rect 3424 -3314 3476 -3262
rect 3488 -3314 3540 -3262
rect 3552 -3314 3604 -3262
rect 4651 -3174 4703 -3122
rect 4715 -3174 4767 -3122
rect 4779 -3174 4831 -3122
rect 1074 -3455 1126 -3403
rect 1138 -3455 1190 -3403
rect 1202 -3455 1254 -3403
rect 2117 -3455 2169 -3403
rect 2181 -3455 2233 -3403
rect 2245 -3455 2297 -3403
rect 2921 -3455 2973 -3403
rect 2985 -3455 3037 -3403
rect 3049 -3455 3101 -3403
rect 4034 -3455 4086 -3403
rect 4098 -3455 4150 -3403
rect 4162 -3455 4214 -3403
rect 1681 -3734 1733 -3682
rect 1745 -3734 1797 -3682
rect 1809 -3734 1861 -3682
rect 2469 -3593 2521 -3541
rect 2533 -3593 2585 -3541
rect 2597 -3593 2649 -3541
rect 3424 -3593 3476 -3541
rect 3488 -3593 3540 -3541
rect 3552 -3593 3604 -3541
rect 5262 -3455 5314 -3403
rect 5326 -3455 5378 -3403
rect 5390 -3455 5442 -3403
rect 4651 -3734 4703 -3682
rect 4715 -3734 4767 -3682
rect 4779 -3734 4831 -3682
rect 1421 -4135 1473 -4083
rect 1485 -4135 1537 -4083
rect 1549 -4135 1601 -4083
rect 1937 -4135 1989 -4083
rect 2001 -4135 2053 -4083
rect 2065 -4135 2117 -4083
rect 2647 -4135 2699 -4083
rect 2711 -4135 2763 -4083
rect 2775 -4135 2827 -4083
rect 3163 -4135 3215 -4083
rect 3227 -4135 3279 -4083
rect 3291 -4135 3343 -4083
rect 3679 -4135 3731 -4083
rect 3743 -4135 3795 -4083
rect 3807 -4135 3859 -4083
rect 4389 -4135 4441 -4083
rect 4453 -4135 4505 -4083
rect 4517 -4135 4569 -4083
rect 4905 -4135 4957 -4083
rect 4969 -4135 5021 -4083
rect 5033 -4135 5085 -4083
rect 1421 -4273 1473 -4221
rect 1485 -4273 1537 -4221
rect 1549 -4273 1601 -4221
rect 1937 -4273 1989 -4221
rect 2001 -4273 2053 -4221
rect 2065 -4273 2117 -4221
rect 2647 -4273 2699 -4221
rect 2711 -4273 2763 -4221
rect 2775 -4273 2827 -4221
rect 3163 -4273 3215 -4221
rect 3227 -4273 3279 -4221
rect 3291 -4273 3343 -4221
rect 3679 -4273 3731 -4221
rect 3743 -4273 3795 -4221
rect 3807 -4273 3859 -4221
rect 4389 -4273 4441 -4221
rect 4453 -4273 4505 -4221
rect 4517 -4273 4569 -4221
rect 4905 -4273 4957 -4221
rect 4969 -4273 5021 -4221
rect 5033 -4273 5085 -4221
rect 1681 -4678 1733 -4626
rect 1745 -4678 1797 -4626
rect 1809 -4678 1861 -4626
rect 2469 -4818 2521 -4766
rect 2533 -4818 2585 -4766
rect 2597 -4818 2649 -4766
rect 3424 -4818 3476 -4766
rect 3488 -4818 3540 -4766
rect 3552 -4818 3604 -4766
rect 4651 -4678 4703 -4626
rect 4715 -4678 4767 -4626
rect 4779 -4678 4831 -4626
rect 1074 -4959 1126 -4907
rect 1138 -4959 1190 -4907
rect 1202 -4959 1254 -4907
rect 2117 -4959 2169 -4907
rect 2181 -4959 2233 -4907
rect 2245 -4959 2297 -4907
rect 2921 -4959 2973 -4907
rect 2985 -4959 3037 -4907
rect 3049 -4959 3101 -4907
rect 4034 -4959 4086 -4907
rect 4098 -4959 4150 -4907
rect 4162 -4959 4214 -4907
rect 5262 -4959 5314 -4907
rect 5326 -4959 5378 -4907
rect 5390 -4959 5442 -4907
<< metal2 >>
rect 505 5348 6057 5356
rect 505 5296 1421 5348
rect 1473 5296 1485 5348
rect 1537 5296 1549 5348
rect 1601 5296 1937 5348
rect 1989 5296 2001 5348
rect 2053 5296 2065 5348
rect 2117 5334 2647 5348
rect 2117 5296 2281 5334
rect 505 5286 2281 5296
rect 2241 5278 2281 5286
rect 2337 5278 2361 5334
rect 2417 5278 2441 5334
rect 2497 5296 2647 5334
rect 2699 5296 2711 5348
rect 2763 5296 2775 5348
rect 2827 5296 3163 5348
rect 3215 5296 3227 5348
rect 3279 5296 3291 5348
rect 3343 5296 3679 5348
rect 3731 5296 3743 5348
rect 3795 5296 3807 5348
rect 3859 5296 4389 5348
rect 4441 5296 4453 5348
rect 4505 5296 4517 5348
rect 4569 5296 4905 5348
rect 4957 5296 4969 5348
rect 5021 5296 5033 5348
rect 5085 5296 6057 5348
rect 2497 5286 6057 5296
rect 2497 5278 2541 5286
rect 2241 5256 2541 5278
rect 5204 4959 5504 4981
rect 5204 4951 5244 4959
rect 505 4943 5244 4951
rect 505 4891 1681 4943
rect 1733 4891 1745 4943
rect 1797 4891 1809 4943
rect 1861 4891 4651 4943
rect 4703 4891 4715 4943
rect 4767 4891 4779 4943
rect 4831 4903 5244 4943
rect 5300 4903 5324 4959
rect 5380 4903 5404 4959
rect 5460 4951 5504 4959
rect 5460 4903 6057 4951
rect 4831 4891 6057 4903
rect 505 4881 6057 4891
rect 3986 4811 4286 4824
rect 505 4803 6057 4811
rect 505 4751 2469 4803
rect 2521 4751 2533 4803
rect 2585 4751 2597 4803
rect 2649 4751 3424 4803
rect 3476 4751 3488 4803
rect 3540 4751 3552 4803
rect 3604 4802 6057 4803
rect 3604 4751 4026 4802
rect 505 4746 4026 4751
rect 4082 4746 4106 4802
rect 4162 4746 4186 4802
rect 4242 4746 6057 4802
rect 505 4741 6057 4746
rect 3986 4724 4286 4741
rect 1001 4680 1301 4702
rect 1001 4672 1041 4680
rect 505 4624 1041 4672
rect 1097 4662 1121 4680
rect 1177 4662 1201 4680
rect 1257 4672 1301 4680
rect 1257 4662 6057 4672
rect 1190 4624 1201 4662
rect 1257 4624 2117 4662
rect 505 4610 1074 4624
rect 1126 4610 1138 4624
rect 1190 4610 1202 4624
rect 1254 4610 2117 4624
rect 2169 4610 2181 4662
rect 2233 4610 2245 4662
rect 2297 4610 2921 4662
rect 2973 4610 2985 4662
rect 3037 4610 3049 4662
rect 3101 4610 4034 4662
rect 4086 4610 4098 4662
rect 4150 4610 4162 4662
rect 4214 4610 5262 4662
rect 5314 4610 5326 4662
rect 5378 4610 5390 4662
rect 5442 4610 6057 4662
rect 505 4602 6057 4610
rect 5204 4532 5504 4545
rect 505 4524 6057 4532
rect 505 4472 2469 4524
rect 2521 4472 2533 4524
rect 2585 4472 2597 4524
rect 2649 4472 3424 4524
rect 3476 4472 3488 4524
rect 3540 4472 3552 4524
rect 3604 4523 6057 4524
rect 3604 4472 5244 4523
rect 505 4467 5244 4472
rect 5300 4467 5324 4523
rect 5380 4467 5404 4523
rect 5460 4467 6057 4523
rect 505 4462 6057 4467
rect 5204 4445 5504 4462
rect 505 4383 6057 4393
rect 505 4331 1681 4383
rect 1733 4331 1745 4383
rect 1797 4331 1809 4383
rect 1861 4371 4651 4383
rect 1861 4331 4026 4371
rect 505 4323 4026 4331
rect 3986 4315 4026 4323
rect 4082 4315 4106 4371
rect 4162 4315 4186 4371
rect 4242 4331 4651 4371
rect 4703 4331 4715 4383
rect 4767 4331 4779 4383
rect 4831 4331 6057 4383
rect 4242 4323 6057 4331
rect 4242 4315 4286 4323
rect 3986 4293 4286 4315
rect 2241 4000 2541 4022
rect 2241 3992 2281 4000
rect 505 3982 2281 3992
rect 505 3930 1421 3982
rect 1473 3930 1485 3982
rect 1537 3930 1549 3982
rect 1601 3930 1937 3982
rect 1989 3930 2001 3982
rect 2053 3930 2065 3982
rect 2117 3944 2281 3982
rect 2337 3944 2361 4000
rect 2417 3944 2441 4000
rect 2497 3992 2541 4000
rect 2497 3982 6057 3992
rect 2497 3944 2647 3982
rect 2117 3930 2647 3944
rect 2699 3930 2711 3982
rect 2763 3930 2775 3982
rect 2827 3930 3163 3982
rect 3215 3930 3227 3982
rect 3279 3930 3291 3982
rect 3343 3930 3679 3982
rect 3731 3930 3743 3982
rect 3795 3930 3807 3982
rect 3859 3930 4389 3982
rect 4441 3930 4453 3982
rect 4505 3930 4517 3982
rect 4569 3930 4905 3982
rect 4957 3930 4969 3982
rect 5021 3930 5033 3982
rect 5085 3930 6057 3982
rect 505 3922 6057 3930
rect 505 3844 6057 3852
rect 505 3792 1421 3844
rect 1473 3792 1485 3844
rect 1537 3792 1549 3844
rect 1601 3792 1937 3844
rect 1989 3792 2001 3844
rect 2053 3792 2065 3844
rect 2117 3830 2647 3844
rect 2117 3792 2281 3830
rect 505 3782 2281 3792
rect 2241 3774 2281 3782
rect 2337 3774 2361 3830
rect 2417 3774 2441 3830
rect 2497 3792 2647 3830
rect 2699 3792 2711 3844
rect 2763 3792 2775 3844
rect 2827 3792 3163 3844
rect 3215 3792 3227 3844
rect 3279 3792 3291 3844
rect 3343 3792 3679 3844
rect 3731 3792 3743 3844
rect 3795 3792 3807 3844
rect 3859 3792 4389 3844
rect 4441 3792 4453 3844
rect 4505 3792 4517 3844
rect 4569 3792 4905 3844
rect 4957 3792 4969 3844
rect 5021 3792 5033 3844
rect 5085 3792 6057 3844
rect 2497 3782 6057 3792
rect 2497 3774 2541 3782
rect 2241 3752 2541 3774
rect 5204 3455 5504 3477
rect 5204 3447 5244 3455
rect 505 3439 5244 3447
rect 505 3387 1681 3439
rect 1733 3387 1745 3439
rect 1797 3387 1809 3439
rect 1861 3387 4651 3439
rect 4703 3387 4715 3439
rect 4767 3387 4779 3439
rect 4831 3399 5244 3439
rect 5300 3399 5324 3455
rect 5380 3399 5404 3455
rect 5460 3447 5504 3455
rect 5460 3399 6057 3447
rect 4831 3387 6057 3399
rect 505 3377 6057 3387
rect 3986 3307 4286 3320
rect 505 3299 6057 3307
rect 505 3247 2469 3299
rect 2521 3247 2533 3299
rect 2585 3247 2597 3299
rect 2649 3247 3424 3299
rect 3476 3247 3488 3299
rect 3540 3247 3552 3299
rect 3604 3298 6057 3299
rect 3604 3247 4026 3298
rect 505 3242 4026 3247
rect 4082 3242 4106 3298
rect 4162 3242 4186 3298
rect 4242 3242 6057 3298
rect 505 3237 6057 3242
rect 3986 3220 4286 3237
rect 1001 3176 1301 3198
rect 1001 3168 1041 3176
rect 505 3120 1041 3168
rect 1097 3158 1121 3176
rect 1177 3158 1201 3176
rect 1257 3168 1301 3176
rect 1257 3158 6057 3168
rect 1190 3120 1201 3158
rect 1257 3120 2117 3158
rect 505 3106 1074 3120
rect 1126 3106 1138 3120
rect 1190 3106 1202 3120
rect 1254 3106 2117 3120
rect 2169 3106 2181 3158
rect 2233 3106 2245 3158
rect 2297 3106 2921 3158
rect 2973 3106 2985 3158
rect 3037 3106 3049 3158
rect 3101 3106 4034 3158
rect 4086 3106 4098 3158
rect 4150 3106 4162 3158
rect 4214 3106 5262 3158
rect 5314 3106 5326 3158
rect 5378 3106 5390 3158
rect 5442 3106 6057 3158
rect 505 3098 6057 3106
rect 5204 3028 5504 3041
rect 505 3020 6057 3028
rect 505 2968 2469 3020
rect 2521 2968 2533 3020
rect 2585 2968 2597 3020
rect 2649 2968 3424 3020
rect 3476 2968 3488 3020
rect 3540 2968 3552 3020
rect 3604 3019 6057 3020
rect 3604 2968 5244 3019
rect 505 2963 5244 2968
rect 5300 2963 5324 3019
rect 5380 2963 5404 3019
rect 5460 2963 6057 3019
rect 505 2958 6057 2963
rect 5204 2941 5504 2958
rect 505 2879 6057 2889
rect 505 2827 1681 2879
rect 1733 2827 1745 2879
rect 1797 2827 1809 2879
rect 1861 2867 4651 2879
rect 1861 2827 4026 2867
rect 505 2819 4026 2827
rect 3986 2811 4026 2819
rect 4082 2811 4106 2867
rect 4162 2811 4186 2867
rect 4242 2827 4651 2867
rect 4703 2827 4715 2879
rect 4767 2827 4779 2879
rect 4831 2827 6057 2879
rect 4242 2819 6057 2827
rect 4242 2811 4286 2819
rect 3986 2789 4286 2811
rect 2241 2496 2541 2518
rect 2241 2488 2281 2496
rect 505 2478 2281 2488
rect 505 2426 1421 2478
rect 1473 2426 1485 2478
rect 1537 2426 1549 2478
rect 1601 2426 1937 2478
rect 1989 2426 2001 2478
rect 2053 2426 2065 2478
rect 2117 2440 2281 2478
rect 2337 2440 2361 2496
rect 2417 2440 2441 2496
rect 2497 2488 2541 2496
rect 2497 2478 6057 2488
rect 2497 2440 2647 2478
rect 2117 2426 2647 2440
rect 2699 2426 2711 2478
rect 2763 2426 2775 2478
rect 2827 2426 3163 2478
rect 3215 2426 3227 2478
rect 3279 2426 3291 2478
rect 3343 2426 3679 2478
rect 3731 2426 3743 2478
rect 3795 2426 3807 2478
rect 3859 2426 4389 2478
rect 4441 2426 4453 2478
rect 4505 2426 4517 2478
rect 4569 2426 4905 2478
rect 4957 2426 4969 2478
rect 5021 2426 5033 2478
rect 5085 2426 6057 2478
rect 505 2418 6057 2426
rect 505 2330 6057 2338
rect 505 2278 1421 2330
rect 1473 2278 1485 2330
rect 1537 2278 1549 2330
rect 1601 2278 1937 2330
rect 1989 2278 2001 2330
rect 2053 2278 2065 2330
rect 2117 2316 2647 2330
rect 2117 2278 2281 2316
rect 505 2268 2281 2278
rect 2241 2260 2281 2268
rect 2337 2260 2361 2316
rect 2417 2260 2441 2316
rect 2497 2278 2647 2316
rect 2699 2278 2711 2330
rect 2763 2278 2775 2330
rect 2827 2278 3163 2330
rect 3215 2278 3227 2330
rect 3279 2278 3291 2330
rect 3343 2278 3679 2330
rect 3731 2278 3743 2330
rect 3795 2278 3807 2330
rect 3859 2278 4389 2330
rect 4441 2278 4453 2330
rect 4505 2278 4517 2330
rect 4569 2278 4905 2330
rect 4957 2278 4969 2330
rect 5021 2278 5033 2330
rect 5085 2278 6057 2330
rect 2497 2268 6057 2278
rect 2497 2260 2541 2268
rect 2241 2238 2541 2260
rect 5204 1947 5504 1969
rect 5204 1939 5244 1947
rect 505 1931 5244 1939
rect 505 1879 1681 1931
rect 1733 1879 1745 1931
rect 1797 1879 1809 1931
rect 1861 1879 4651 1931
rect 4703 1879 4715 1931
rect 4767 1879 4779 1931
rect 4831 1891 5244 1931
rect 5300 1891 5324 1947
rect 5380 1891 5404 1947
rect 5460 1939 5504 1947
rect 5460 1891 6057 1939
rect 4831 1879 6057 1891
rect 505 1869 6057 1879
rect 3986 1807 4286 1829
rect 3986 1799 4026 1807
rect 505 1791 4026 1799
rect 505 1739 2469 1791
rect 2521 1739 2533 1791
rect 2585 1739 2597 1791
rect 2649 1739 3424 1791
rect 3476 1739 3488 1791
rect 3540 1739 3552 1791
rect 3604 1751 4026 1791
rect 4082 1751 4106 1807
rect 4162 1751 4186 1807
rect 4242 1799 4286 1807
rect 4242 1751 6057 1799
rect 3604 1739 6057 1751
rect 505 1729 6057 1739
rect 1001 1668 1301 1690
rect 1001 1660 1041 1668
rect 505 1612 1041 1660
rect 1097 1650 1121 1668
rect 1177 1650 1201 1668
rect 1257 1660 1301 1668
rect 1257 1650 6057 1660
rect 1190 1612 1201 1650
rect 1257 1612 2117 1650
rect 505 1598 1074 1612
rect 1126 1598 1138 1612
rect 1190 1598 1202 1612
rect 1254 1598 2117 1612
rect 2169 1598 2181 1650
rect 2233 1598 2245 1650
rect 2297 1598 2921 1650
rect 2973 1598 2985 1650
rect 3037 1598 3049 1650
rect 3101 1598 4034 1650
rect 4086 1598 4098 1650
rect 4150 1598 4162 1650
rect 4214 1598 5262 1650
rect 5314 1598 5326 1650
rect 5378 1598 5390 1650
rect 5442 1598 6057 1650
rect 505 1590 6057 1598
rect 505 1510 6057 1520
rect 505 1458 1681 1510
rect 1733 1458 1745 1510
rect 1797 1458 1809 1510
rect 1861 1498 2478 1510
rect 1861 1458 2281 1498
rect 505 1450 2281 1458
rect 2241 1442 2281 1450
rect 2337 1442 2361 1498
rect 2417 1442 2441 1498
rect 2530 1458 2542 1510
rect 2594 1458 2606 1510
rect 2658 1458 3424 1510
rect 3476 1458 3488 1510
rect 3540 1458 3552 1510
rect 3604 1458 4651 1510
rect 4703 1458 4715 1510
rect 4767 1458 4779 1510
rect 4831 1458 6057 1510
rect 2497 1450 6057 1458
rect 2497 1442 2541 1450
rect 2241 1420 2541 1442
rect 2241 1129 2541 1151
rect 2241 1121 2281 1129
rect 505 1111 2281 1121
rect 505 1059 1421 1111
rect 1473 1059 1485 1111
rect 1537 1059 1549 1111
rect 1601 1059 1937 1111
rect 1989 1059 2001 1111
rect 2053 1059 2065 1111
rect 2117 1073 2281 1111
rect 2337 1073 2361 1129
rect 2417 1073 2441 1129
rect 2497 1121 2541 1129
rect 2497 1111 6057 1121
rect 2497 1073 2647 1111
rect 2117 1059 2647 1073
rect 2699 1059 2711 1111
rect 2763 1059 2775 1111
rect 2827 1059 3163 1111
rect 3215 1059 3227 1111
rect 3279 1059 3291 1111
rect 3343 1059 3679 1111
rect 3731 1059 3743 1111
rect 3795 1059 3807 1111
rect 3859 1059 4389 1111
rect 4441 1059 4453 1111
rect 4505 1059 4517 1111
rect 4569 1059 4905 1111
rect 4957 1059 4969 1111
rect 5021 1059 5033 1111
rect 5085 1059 6057 1111
rect 505 1051 6057 1059
rect 505 963 6057 971
rect 505 911 1421 963
rect 1473 911 1485 963
rect 1537 911 1549 963
rect 1601 911 1937 963
rect 1989 911 2001 963
rect 2053 911 2065 963
rect 2117 949 2647 963
rect 2117 911 2281 949
rect 505 901 2281 911
rect 2241 893 2281 901
rect 2337 893 2361 949
rect 2417 893 2441 949
rect 2497 911 2647 949
rect 2699 911 2711 963
rect 2763 911 2775 963
rect 2827 911 3163 963
rect 3215 911 3227 963
rect 3279 911 3291 963
rect 3343 911 3679 963
rect 3731 911 3743 963
rect 3795 911 3807 963
rect 3859 911 4389 963
rect 4441 911 4453 963
rect 4505 911 4517 963
rect 4569 911 4905 963
rect 4957 911 4969 963
rect 5021 911 5033 963
rect 5085 911 6057 963
rect 2497 901 6057 911
rect 2497 893 2541 901
rect 2241 871 2541 893
rect 1001 578 1301 600
rect 1001 570 1041 578
rect 505 522 1041 570
rect 1097 560 1121 578
rect 1177 560 1201 578
rect 1257 570 1301 578
rect 2688 570 6057 571
rect 1257 560 6057 570
rect 1190 522 1201 560
rect 1257 522 2121 560
rect 505 508 1074 522
rect 1126 508 1138 522
rect 1190 508 1202 522
rect 1254 508 2121 522
rect 2173 508 2185 560
rect 2237 508 2249 560
rect 2301 508 2921 560
rect 2973 508 2985 560
rect 3037 508 3049 560
rect 3101 508 4034 560
rect 4086 508 4098 560
rect 4150 508 4162 560
rect 4214 508 5262 560
rect 5314 508 5326 560
rect 5378 508 5390 560
rect 5442 508 6057 560
rect 505 501 6057 508
rect 505 500 2771 501
rect 2241 432 2541 433
rect 2688 432 6057 433
rect 505 423 6057 432
rect 505 371 1681 423
rect 1733 371 1745 423
rect 1797 371 1809 423
rect 1861 411 2478 423
rect 1861 371 2281 411
rect 505 362 2281 371
rect 2241 355 2281 362
rect 2337 355 2361 411
rect 2417 355 2441 411
rect 2530 371 2542 423
rect 2594 371 2606 423
rect 2658 371 3424 423
rect 3476 371 3488 423
rect 3540 371 3552 423
rect 3604 371 4651 423
rect 4703 371 4715 423
rect 4767 371 4779 423
rect 4831 371 6057 423
rect 2497 363 6057 371
rect 2497 362 2771 363
rect 2497 355 2541 362
rect 2241 333 2541 355
rect 2241 35 2541 57
rect 2241 27 2281 35
rect 505 17 2281 27
rect 505 -35 1421 17
rect 1473 -35 1485 17
rect 1537 -35 1549 17
rect 1601 -35 1937 17
rect 1989 -35 2001 17
rect 2053 -35 2065 17
rect 2117 -21 2281 17
rect 2337 -21 2361 35
rect 2417 -21 2441 35
rect 2497 27 2541 35
rect 2497 17 6057 27
rect 2497 -21 2647 17
rect 2117 -35 2647 -21
rect 2699 -35 2711 17
rect 2763 -35 2775 17
rect 2827 -35 3163 17
rect 3215 -35 3227 17
rect 3279 -35 3291 17
rect 3343 -35 3679 17
rect 3731 -35 3743 17
rect 3795 -35 3807 17
rect 3859 -35 4389 17
rect 4441 -35 4453 17
rect 4505 -35 4517 17
rect 4569 -35 4905 17
rect 4957 -35 4969 17
rect 5021 -35 5033 17
rect 5085 -35 6057 17
rect 505 -43 6057 -35
rect 505 -132 6057 -124
rect 505 -184 1421 -132
rect 1473 -184 1485 -132
rect 1537 -184 1549 -132
rect 1601 -184 1937 -132
rect 1989 -184 2001 -132
rect 2053 -184 2065 -132
rect 2117 -146 2647 -132
rect 2117 -184 2281 -146
rect 505 -194 2281 -184
rect 2241 -202 2281 -194
rect 2337 -202 2361 -146
rect 2417 -202 2441 -146
rect 2497 -184 2647 -146
rect 2699 -184 2711 -132
rect 2763 -184 2775 -132
rect 2827 -184 3163 -132
rect 3215 -184 3227 -132
rect 3279 -184 3291 -132
rect 3343 -184 3679 -132
rect 3731 -184 3743 -132
rect 3795 -184 3807 -132
rect 3859 -184 4389 -132
rect 4441 -184 4453 -132
rect 4505 -184 4517 -132
rect 4569 -184 4905 -132
rect 4957 -184 4969 -132
rect 5021 -184 5033 -132
rect 5085 -184 6057 -132
rect 2497 -194 6057 -184
rect 2497 -202 2541 -194
rect 2241 -224 2541 -202
rect 1001 -514 1301 -492
rect 1001 -522 1041 -514
rect 505 -570 1041 -522
rect 1097 -532 1121 -514
rect 1177 -532 1201 -514
rect 1257 -522 1301 -514
rect 1190 -570 1201 -532
rect 1257 -533 6057 -522
rect 1257 -570 2119 -533
rect 505 -584 1074 -570
rect 1126 -584 1138 -570
rect 1190 -584 1202 -570
rect 1254 -584 2119 -570
rect 505 -585 2119 -584
rect 2171 -585 2183 -533
rect 2235 -585 2247 -533
rect 2299 -585 2921 -533
rect 2973 -585 2985 -533
rect 3037 -585 3049 -533
rect 3101 -585 4034 -533
rect 4086 -585 4098 -533
rect 4150 -585 4162 -533
rect 4214 -585 5262 -533
rect 5314 -585 5326 -533
rect 5378 -585 5390 -533
rect 5442 -585 6057 -533
rect 505 -592 6057 -585
rect 2290 -593 2574 -592
rect 2914 -593 3110 -592
rect 5253 -593 5449 -592
rect 505 -672 6057 -662
rect 505 -724 1681 -672
rect 1733 -724 1745 -672
rect 1797 -724 1809 -672
rect 1861 -684 2478 -672
rect 1861 -724 2281 -684
rect 505 -732 2281 -724
rect 2241 -740 2281 -732
rect 2337 -740 2361 -684
rect 2417 -740 2441 -684
rect 2530 -724 2542 -672
rect 2594 -724 2606 -672
rect 2658 -724 3424 -672
rect 3476 -724 3488 -672
rect 3540 -724 3552 -672
rect 3604 -724 4651 -672
rect 4703 -724 4715 -672
rect 4767 -724 4779 -672
rect 4831 -724 6057 -672
rect 2497 -732 6057 -724
rect 2497 -740 2541 -732
rect 2241 -762 2541 -740
rect 2241 -1057 2541 -1035
rect 2241 -1065 2281 -1057
rect 505 -1075 2281 -1065
rect 505 -1127 1421 -1075
rect 1473 -1127 1485 -1075
rect 1537 -1127 1549 -1075
rect 1601 -1127 1937 -1075
rect 1989 -1127 2001 -1075
rect 2053 -1127 2065 -1075
rect 2117 -1113 2281 -1075
rect 2337 -1113 2361 -1057
rect 2417 -1113 2441 -1057
rect 2497 -1065 2541 -1057
rect 2497 -1075 6057 -1065
rect 2497 -1113 2647 -1075
rect 2117 -1127 2647 -1113
rect 2699 -1127 2711 -1075
rect 2763 -1127 2775 -1075
rect 2827 -1127 3163 -1075
rect 3215 -1127 3227 -1075
rect 3279 -1127 3291 -1075
rect 3343 -1127 3679 -1075
rect 3731 -1127 3743 -1075
rect 3795 -1127 3807 -1075
rect 3859 -1127 4389 -1075
rect 4441 -1127 4453 -1075
rect 4505 -1127 4517 -1075
rect 4569 -1127 4905 -1075
rect 4957 -1127 4969 -1075
rect 5021 -1127 5033 -1075
rect 5085 -1127 6057 -1075
rect 505 -1135 6057 -1127
rect 505 -1213 6057 -1205
rect 505 -1265 1421 -1213
rect 1473 -1265 1485 -1213
rect 1537 -1265 1549 -1213
rect 1601 -1265 1937 -1213
rect 1989 -1265 2001 -1213
rect 2053 -1265 2065 -1213
rect 2117 -1227 2647 -1213
rect 2117 -1265 2281 -1227
rect 505 -1275 2281 -1265
rect 2241 -1283 2281 -1275
rect 2337 -1283 2361 -1227
rect 2417 -1283 2441 -1227
rect 2497 -1265 2647 -1227
rect 2699 -1265 2711 -1213
rect 2763 -1265 2775 -1213
rect 2827 -1265 3163 -1213
rect 3215 -1265 3227 -1213
rect 3279 -1265 3291 -1213
rect 3343 -1265 3679 -1213
rect 3731 -1265 3743 -1213
rect 3795 -1265 3807 -1213
rect 3859 -1265 4389 -1213
rect 4441 -1265 4453 -1213
rect 4505 -1265 4517 -1213
rect 4569 -1265 4905 -1213
rect 4957 -1265 4969 -1213
rect 5021 -1265 5033 -1213
rect 5085 -1265 6057 -1213
rect 2497 -1275 6057 -1265
rect 2497 -1283 2541 -1275
rect 2241 -1305 2541 -1283
rect 3986 -1602 4286 -1580
rect 3986 -1610 4026 -1602
rect 505 -1618 4026 -1610
rect 505 -1670 1681 -1618
rect 1733 -1670 1745 -1618
rect 1797 -1670 1809 -1618
rect 1861 -1658 4026 -1618
rect 4082 -1658 4106 -1602
rect 4162 -1658 4186 -1602
rect 4242 -1610 4286 -1602
rect 4242 -1618 6057 -1610
rect 4242 -1658 4651 -1618
rect 1861 -1670 4651 -1658
rect 4703 -1670 4715 -1618
rect 4767 -1670 4779 -1618
rect 4831 -1670 6057 -1618
rect 505 -1680 6057 -1670
rect 5204 -1750 5504 -1728
rect 505 -1758 5244 -1750
rect 505 -1810 2469 -1758
rect 2521 -1810 2533 -1758
rect 2585 -1810 2597 -1758
rect 2649 -1810 3424 -1758
rect 3476 -1810 3488 -1758
rect 3540 -1810 3552 -1758
rect 3604 -1806 5244 -1758
rect 5300 -1806 5324 -1750
rect 5380 -1806 5404 -1750
rect 5460 -1806 6057 -1750
rect 3604 -1810 6057 -1806
rect 505 -1820 6057 -1810
rect 5204 -1828 5504 -1820
rect 1001 -1881 1301 -1859
rect 1001 -1889 1041 -1881
rect 505 -1937 1041 -1889
rect 1097 -1899 1121 -1881
rect 1177 -1899 1201 -1881
rect 1257 -1889 1301 -1881
rect 1257 -1899 6057 -1889
rect 1190 -1937 1201 -1899
rect 1257 -1937 2117 -1899
rect 505 -1951 1074 -1937
rect 1126 -1951 1138 -1937
rect 1190 -1951 1202 -1937
rect 1254 -1951 2117 -1937
rect 2169 -1951 2181 -1899
rect 2233 -1951 2245 -1899
rect 2297 -1951 2921 -1899
rect 2973 -1951 2985 -1899
rect 3037 -1951 3049 -1899
rect 3101 -1951 4034 -1899
rect 4086 -1951 4098 -1899
rect 4150 -1951 4162 -1899
rect 4214 -1951 5262 -1899
rect 5314 -1951 5326 -1899
rect 5378 -1951 5390 -1899
rect 5442 -1951 6057 -1899
rect 505 -1959 6057 -1951
rect 3986 -2029 4286 -2016
rect 505 -2037 6057 -2029
rect 505 -2089 2469 -2037
rect 2521 -2089 2533 -2037
rect 2585 -2089 2597 -2037
rect 2649 -2089 3424 -2037
rect 3476 -2089 3488 -2037
rect 3540 -2089 3552 -2037
rect 3604 -2038 6057 -2037
rect 3604 -2089 4026 -2038
rect 505 -2094 4026 -2089
rect 4082 -2094 4106 -2038
rect 4162 -2094 4186 -2038
rect 4242 -2094 6057 -2038
rect 505 -2099 6057 -2094
rect 3986 -2116 4286 -2099
rect 505 -2178 6057 -2168
rect 505 -2230 1681 -2178
rect 1733 -2230 1745 -2178
rect 1797 -2230 1809 -2178
rect 1861 -2230 4651 -2178
rect 4703 -2230 4715 -2178
rect 4767 -2230 4779 -2178
rect 4831 -2190 6057 -2178
rect 4831 -2230 5244 -2190
rect 505 -2238 5244 -2230
rect 5204 -2246 5244 -2238
rect 5300 -2246 5324 -2190
rect 5380 -2246 5404 -2190
rect 5460 -2238 6057 -2190
rect 5460 -2246 5504 -2238
rect 5204 -2268 5504 -2246
rect 2241 -2561 2541 -2539
rect 2241 -2569 2281 -2561
rect 505 -2579 2281 -2569
rect 505 -2631 1421 -2579
rect 1473 -2631 1485 -2579
rect 1537 -2631 1549 -2579
rect 1601 -2631 1937 -2579
rect 1989 -2631 2001 -2579
rect 2053 -2631 2065 -2579
rect 2117 -2617 2281 -2579
rect 2337 -2617 2361 -2561
rect 2417 -2617 2441 -2561
rect 2497 -2569 2541 -2561
rect 2497 -2579 6057 -2569
rect 2497 -2617 2647 -2579
rect 2117 -2631 2647 -2617
rect 2699 -2631 2711 -2579
rect 2763 -2631 2775 -2579
rect 2827 -2631 3163 -2579
rect 3215 -2631 3227 -2579
rect 3279 -2631 3291 -2579
rect 3343 -2631 3679 -2579
rect 3731 -2631 3743 -2579
rect 3795 -2631 3807 -2579
rect 3859 -2631 4389 -2579
rect 4441 -2631 4453 -2579
rect 4505 -2631 4517 -2579
rect 4569 -2631 4905 -2579
rect 4957 -2631 4969 -2579
rect 5021 -2631 5033 -2579
rect 5085 -2631 6057 -2579
rect 505 -2639 6057 -2631
rect 505 -2717 6057 -2709
rect 505 -2769 1421 -2717
rect 1473 -2769 1485 -2717
rect 1537 -2769 1549 -2717
rect 1601 -2769 1937 -2717
rect 1989 -2769 2001 -2717
rect 2053 -2769 2065 -2717
rect 2117 -2731 2647 -2717
rect 2117 -2769 2281 -2731
rect 505 -2779 2281 -2769
rect 2241 -2787 2281 -2779
rect 2337 -2787 2361 -2731
rect 2417 -2787 2441 -2731
rect 2497 -2769 2647 -2731
rect 2699 -2769 2711 -2717
rect 2763 -2769 2775 -2717
rect 2827 -2769 3163 -2717
rect 3215 -2769 3227 -2717
rect 3279 -2769 3291 -2717
rect 3343 -2769 3679 -2717
rect 3731 -2769 3743 -2717
rect 3795 -2769 3807 -2717
rect 3859 -2769 4389 -2717
rect 4441 -2769 4453 -2717
rect 4505 -2769 4517 -2717
rect 4569 -2769 4905 -2717
rect 4957 -2769 4969 -2717
rect 5021 -2769 5033 -2717
rect 5085 -2769 6057 -2717
rect 2497 -2779 6057 -2769
rect 2497 -2787 2541 -2779
rect 2241 -2809 2541 -2787
rect 3986 -3106 4286 -3084
rect 3986 -3114 4026 -3106
rect 505 -3122 4026 -3114
rect 505 -3174 1681 -3122
rect 1733 -3174 1745 -3122
rect 1797 -3174 1809 -3122
rect 1861 -3162 4026 -3122
rect 4082 -3162 4106 -3106
rect 4162 -3162 4186 -3106
rect 4242 -3114 4286 -3106
rect 4242 -3122 6057 -3114
rect 4242 -3162 4651 -3122
rect 1861 -3174 4651 -3162
rect 4703 -3174 4715 -3122
rect 4767 -3174 4779 -3122
rect 4831 -3174 6057 -3122
rect 505 -3184 6057 -3174
rect 5204 -3246 5504 -3224
rect 5204 -3254 5244 -3246
rect 505 -3262 5244 -3254
rect 505 -3314 2469 -3262
rect 2521 -3314 2533 -3262
rect 2585 -3314 2597 -3262
rect 2649 -3314 3424 -3262
rect 3476 -3314 3488 -3262
rect 3540 -3314 3552 -3262
rect 3604 -3302 5244 -3262
rect 5300 -3302 5324 -3246
rect 5380 -3302 5404 -3246
rect 5460 -3254 5504 -3246
rect 5460 -3302 6057 -3254
rect 3604 -3314 6057 -3302
rect 505 -3324 6057 -3314
rect 1001 -3385 1301 -3363
rect 1001 -3393 1041 -3385
rect 505 -3441 1041 -3393
rect 1097 -3403 1121 -3385
rect 1177 -3403 1201 -3385
rect 1257 -3393 1301 -3385
rect 1257 -3403 6057 -3393
rect 1190 -3441 1201 -3403
rect 1257 -3441 2117 -3403
rect 505 -3455 1074 -3441
rect 1126 -3455 1138 -3441
rect 1190 -3455 1202 -3441
rect 1254 -3455 2117 -3441
rect 2169 -3455 2181 -3403
rect 2233 -3455 2245 -3403
rect 2297 -3455 2921 -3403
rect 2973 -3455 2985 -3403
rect 3037 -3455 3049 -3403
rect 3101 -3455 4034 -3403
rect 4086 -3455 4098 -3403
rect 4150 -3455 4162 -3403
rect 4214 -3455 5262 -3403
rect 5314 -3455 5326 -3403
rect 5378 -3455 5390 -3403
rect 5442 -3455 6057 -3403
rect 505 -3463 6057 -3455
rect 3986 -3533 4286 -3520
rect 505 -3541 6057 -3533
rect 505 -3593 2469 -3541
rect 2521 -3593 2533 -3541
rect 2585 -3593 2597 -3541
rect 2649 -3593 3424 -3541
rect 3476 -3593 3488 -3541
rect 3540 -3593 3552 -3541
rect 3604 -3542 6057 -3541
rect 3604 -3593 4026 -3542
rect 505 -3598 4026 -3593
rect 4082 -3598 4106 -3542
rect 4162 -3598 4186 -3542
rect 4242 -3598 6057 -3542
rect 505 -3603 6057 -3598
rect 3986 -3620 4286 -3603
rect 505 -3682 6057 -3672
rect 505 -3734 1681 -3682
rect 1733 -3734 1745 -3682
rect 1797 -3734 1809 -3682
rect 1861 -3734 4651 -3682
rect 4703 -3734 4715 -3682
rect 4767 -3734 4779 -3682
rect 4831 -3694 6057 -3682
rect 4831 -3734 5244 -3694
rect 505 -3742 5244 -3734
rect 5204 -3750 5244 -3742
rect 5300 -3750 5324 -3694
rect 5380 -3750 5404 -3694
rect 5460 -3742 6057 -3694
rect 5460 -3750 5504 -3742
rect 5204 -3772 5504 -3750
rect 2241 -4065 2541 -4043
rect 2241 -4073 2281 -4065
rect 505 -4083 2281 -4073
rect 505 -4135 1421 -4083
rect 1473 -4135 1485 -4083
rect 1537 -4135 1549 -4083
rect 1601 -4135 1937 -4083
rect 1989 -4135 2001 -4083
rect 2053 -4135 2065 -4083
rect 2117 -4121 2281 -4083
rect 2337 -4121 2361 -4065
rect 2417 -4121 2441 -4065
rect 2497 -4073 2541 -4065
rect 2497 -4083 6057 -4073
rect 2497 -4121 2647 -4083
rect 2117 -4135 2647 -4121
rect 2699 -4135 2711 -4083
rect 2763 -4135 2775 -4083
rect 2827 -4135 3163 -4083
rect 3215 -4135 3227 -4083
rect 3279 -4135 3291 -4083
rect 3343 -4135 3679 -4083
rect 3731 -4135 3743 -4083
rect 3795 -4135 3807 -4083
rect 3859 -4135 4389 -4083
rect 4441 -4135 4453 -4083
rect 4505 -4135 4517 -4083
rect 4569 -4135 4905 -4083
rect 4957 -4135 4969 -4083
rect 5021 -4135 5033 -4083
rect 5085 -4135 6057 -4083
rect 505 -4143 6057 -4135
rect 505 -4221 6057 -4213
rect 505 -4273 1421 -4221
rect 1473 -4273 1485 -4221
rect 1537 -4273 1549 -4221
rect 1601 -4273 1937 -4221
rect 1989 -4273 2001 -4221
rect 2053 -4273 2065 -4221
rect 2117 -4235 2647 -4221
rect 2117 -4273 2281 -4235
rect 505 -4283 2281 -4273
rect 2241 -4291 2281 -4283
rect 2337 -4291 2361 -4235
rect 2417 -4291 2441 -4235
rect 2497 -4273 2647 -4235
rect 2699 -4273 2711 -4221
rect 2763 -4273 2775 -4221
rect 2827 -4273 3163 -4221
rect 3215 -4273 3227 -4221
rect 3279 -4273 3291 -4221
rect 3343 -4273 3679 -4221
rect 3731 -4273 3743 -4221
rect 3795 -4273 3807 -4221
rect 3859 -4273 4389 -4221
rect 4441 -4273 4453 -4221
rect 4505 -4273 4517 -4221
rect 4569 -4273 4905 -4221
rect 4957 -4273 4969 -4221
rect 5021 -4273 5033 -4221
rect 5085 -4273 6057 -4221
rect 2497 -4283 6057 -4273
rect 2497 -4291 2541 -4283
rect 2241 -4313 2541 -4291
rect 3986 -4610 4286 -4588
rect 3986 -4618 4026 -4610
rect 505 -4626 4026 -4618
rect 505 -4678 1681 -4626
rect 1733 -4678 1745 -4626
rect 1797 -4678 1809 -4626
rect 1861 -4666 4026 -4626
rect 4082 -4666 4106 -4610
rect 4162 -4666 4186 -4610
rect 4242 -4618 4286 -4610
rect 4242 -4626 6057 -4618
rect 4242 -4666 4651 -4626
rect 1861 -4678 4651 -4666
rect 4703 -4678 4715 -4626
rect 4767 -4678 4779 -4626
rect 4831 -4678 6057 -4626
rect 505 -4688 6057 -4678
rect 5204 -4758 5504 -4745
rect 505 -4766 6057 -4758
rect 505 -4818 2469 -4766
rect 2521 -4818 2533 -4766
rect 2585 -4818 2597 -4766
rect 2649 -4818 3424 -4766
rect 3476 -4818 3488 -4766
rect 3540 -4818 3552 -4766
rect 3604 -4767 6057 -4766
rect 3604 -4818 5244 -4767
rect 505 -4823 5244 -4818
rect 5300 -4823 5324 -4767
rect 5380 -4823 5404 -4767
rect 5460 -4823 6057 -4767
rect 505 -4828 6057 -4823
rect 5204 -4845 5504 -4828
rect 1001 -4889 1301 -4867
rect 1001 -4897 1041 -4889
rect 505 -4945 1041 -4897
rect 1097 -4907 1121 -4889
rect 1177 -4907 1201 -4889
rect 1257 -4897 1301 -4889
rect 1257 -4907 6057 -4897
rect 1190 -4945 1201 -4907
rect 1257 -4945 2117 -4907
rect 505 -4959 1074 -4945
rect 1126 -4959 1138 -4945
rect 1190 -4959 1202 -4945
rect 1254 -4959 2117 -4945
rect 2169 -4959 2181 -4907
rect 2233 -4959 2245 -4907
rect 2297 -4959 2921 -4907
rect 2973 -4959 2985 -4907
rect 3037 -4959 3049 -4907
rect 3101 -4959 4034 -4907
rect 4086 -4959 4098 -4907
rect 4150 -4959 4162 -4907
rect 4214 -4959 5262 -4907
rect 5314 -4959 5326 -4907
rect 5378 -4959 5390 -4907
rect 5442 -4959 6057 -4907
rect 505 -4967 6057 -4959
<< via2 >>
rect 2281 5278 2337 5334
rect 2361 5278 2417 5334
rect 2441 5278 2497 5334
rect 5244 4903 5300 4959
rect 5324 4903 5380 4959
rect 5404 4903 5460 4959
rect 4026 4746 4082 4802
rect 4106 4746 4162 4802
rect 4186 4746 4242 4802
rect 1041 4662 1097 4680
rect 1121 4662 1177 4680
rect 1201 4662 1257 4680
rect 1041 4624 1074 4662
rect 1074 4624 1097 4662
rect 1121 4624 1126 4662
rect 1126 4624 1138 4662
rect 1138 4624 1177 4662
rect 1201 4624 1202 4662
rect 1202 4624 1254 4662
rect 1254 4624 1257 4662
rect 5244 4467 5300 4523
rect 5324 4467 5380 4523
rect 5404 4467 5460 4523
rect 4026 4315 4082 4371
rect 4106 4315 4162 4371
rect 4186 4315 4242 4371
rect 2281 3944 2337 4000
rect 2361 3944 2417 4000
rect 2441 3944 2497 4000
rect 2281 3774 2337 3830
rect 2361 3774 2417 3830
rect 2441 3774 2497 3830
rect 5244 3399 5300 3455
rect 5324 3399 5380 3455
rect 5404 3399 5460 3455
rect 4026 3242 4082 3298
rect 4106 3242 4162 3298
rect 4186 3242 4242 3298
rect 1041 3158 1097 3176
rect 1121 3158 1177 3176
rect 1201 3158 1257 3176
rect 1041 3120 1074 3158
rect 1074 3120 1097 3158
rect 1121 3120 1126 3158
rect 1126 3120 1138 3158
rect 1138 3120 1177 3158
rect 1201 3120 1202 3158
rect 1202 3120 1254 3158
rect 1254 3120 1257 3158
rect 5244 2963 5300 3019
rect 5324 2963 5380 3019
rect 5404 2963 5460 3019
rect 4026 2811 4082 2867
rect 4106 2811 4162 2867
rect 4186 2811 4242 2867
rect 2281 2440 2337 2496
rect 2361 2440 2417 2496
rect 2441 2440 2497 2496
rect 2281 2260 2337 2316
rect 2361 2260 2417 2316
rect 2441 2260 2497 2316
rect 5244 1891 5300 1947
rect 5324 1891 5380 1947
rect 5404 1891 5460 1947
rect 4026 1751 4082 1807
rect 4106 1751 4162 1807
rect 4186 1751 4242 1807
rect 1041 1650 1097 1668
rect 1121 1650 1177 1668
rect 1201 1650 1257 1668
rect 1041 1612 1074 1650
rect 1074 1612 1097 1650
rect 1121 1612 1126 1650
rect 1126 1612 1138 1650
rect 1138 1612 1177 1650
rect 1201 1612 1202 1650
rect 1202 1612 1254 1650
rect 1254 1612 1257 1650
rect 2281 1442 2337 1498
rect 2361 1442 2417 1498
rect 2441 1458 2478 1498
rect 2478 1458 2497 1498
rect 2441 1442 2497 1458
rect 2281 1073 2337 1129
rect 2361 1073 2417 1129
rect 2441 1073 2497 1129
rect 2281 893 2337 949
rect 2361 893 2417 949
rect 2441 893 2497 949
rect 1041 560 1097 578
rect 1121 560 1177 578
rect 1201 560 1257 578
rect 1041 522 1074 560
rect 1074 522 1097 560
rect 1121 522 1126 560
rect 1126 522 1138 560
rect 1138 522 1177 560
rect 1201 522 1202 560
rect 1202 522 1254 560
rect 1254 522 1257 560
rect 2281 355 2337 411
rect 2361 355 2417 411
rect 2441 371 2478 411
rect 2478 371 2497 411
rect 2441 355 2497 371
rect 2281 -21 2337 35
rect 2361 -21 2417 35
rect 2441 -21 2497 35
rect 2281 -202 2337 -146
rect 2361 -202 2417 -146
rect 2441 -202 2497 -146
rect 1041 -532 1097 -514
rect 1121 -532 1177 -514
rect 1201 -532 1257 -514
rect 1041 -570 1074 -532
rect 1074 -570 1097 -532
rect 1121 -570 1126 -532
rect 1126 -570 1138 -532
rect 1138 -570 1177 -532
rect 1201 -570 1202 -532
rect 1202 -570 1254 -532
rect 1254 -570 1257 -532
rect 2281 -740 2337 -684
rect 2361 -740 2417 -684
rect 2441 -724 2478 -684
rect 2478 -724 2497 -684
rect 2441 -740 2497 -724
rect 2281 -1113 2337 -1057
rect 2361 -1113 2417 -1057
rect 2441 -1113 2497 -1057
rect 2281 -1283 2337 -1227
rect 2361 -1283 2417 -1227
rect 2441 -1283 2497 -1227
rect 4026 -1658 4082 -1602
rect 4106 -1658 4162 -1602
rect 4186 -1658 4242 -1602
rect 5244 -1806 5300 -1750
rect 5324 -1806 5380 -1750
rect 5404 -1806 5460 -1750
rect 1041 -1899 1097 -1881
rect 1121 -1899 1177 -1881
rect 1201 -1899 1257 -1881
rect 1041 -1937 1074 -1899
rect 1074 -1937 1097 -1899
rect 1121 -1937 1126 -1899
rect 1126 -1937 1138 -1899
rect 1138 -1937 1177 -1899
rect 1201 -1937 1202 -1899
rect 1202 -1937 1254 -1899
rect 1254 -1937 1257 -1899
rect 4026 -2094 4082 -2038
rect 4106 -2094 4162 -2038
rect 4186 -2094 4242 -2038
rect 5244 -2246 5300 -2190
rect 5324 -2246 5380 -2190
rect 5404 -2246 5460 -2190
rect 2281 -2617 2337 -2561
rect 2361 -2617 2417 -2561
rect 2441 -2617 2497 -2561
rect 2281 -2787 2337 -2731
rect 2361 -2787 2417 -2731
rect 2441 -2787 2497 -2731
rect 4026 -3162 4082 -3106
rect 4106 -3162 4162 -3106
rect 4186 -3162 4242 -3106
rect 5244 -3302 5300 -3246
rect 5324 -3302 5380 -3246
rect 5404 -3302 5460 -3246
rect 1041 -3403 1097 -3385
rect 1121 -3403 1177 -3385
rect 1201 -3403 1257 -3385
rect 1041 -3441 1074 -3403
rect 1074 -3441 1097 -3403
rect 1121 -3441 1126 -3403
rect 1126 -3441 1138 -3403
rect 1138 -3441 1177 -3403
rect 1201 -3441 1202 -3403
rect 1202 -3441 1254 -3403
rect 1254 -3441 1257 -3403
rect 4026 -3598 4082 -3542
rect 4106 -3598 4162 -3542
rect 4186 -3598 4242 -3542
rect 5244 -3750 5300 -3694
rect 5324 -3750 5380 -3694
rect 5404 -3750 5460 -3694
rect 2281 -4121 2337 -4065
rect 2361 -4121 2417 -4065
rect 2441 -4121 2497 -4065
rect 2281 -4291 2337 -4235
rect 2361 -4291 2417 -4235
rect 2441 -4291 2497 -4235
rect 4026 -4666 4082 -4610
rect 4106 -4666 4162 -4610
rect 4186 -4666 4242 -4610
rect 5244 -4823 5300 -4767
rect 5324 -4823 5380 -4767
rect 5404 -4823 5460 -4767
rect 1041 -4907 1097 -4889
rect 1121 -4907 1177 -4889
rect 1201 -4907 1257 -4889
rect 1041 -4945 1074 -4907
rect 1074 -4945 1097 -4907
rect 1121 -4945 1126 -4907
rect 1126 -4945 1138 -4907
rect 1138 -4945 1177 -4907
rect 1201 -4945 1202 -4907
rect 1202 -4945 1254 -4907
rect 1254 -4945 1257 -4907
<< metal3 >>
rect 2241 5334 2541 5463
rect 2241 5278 2281 5334
rect 2337 5278 2361 5334
rect 2417 5278 2441 5334
rect 2497 5278 2541 5334
rect 1001 4680 1301 4710
rect 1001 4624 1041 4680
rect 1097 4624 1121 4680
rect 1177 4624 1201 4680
rect 1257 4624 1301 4680
rect 1001 3176 1301 4624
rect 1001 3120 1041 3176
rect 1097 3120 1121 3176
rect 1177 3120 1201 3176
rect 1257 3120 1301 3176
rect 1001 1668 1301 3120
rect 1001 1612 1041 1668
rect 1097 1612 1121 1668
rect 1177 1612 1201 1668
rect 1257 1612 1301 1668
rect 1001 578 1301 1612
rect 1001 522 1041 578
rect 1097 522 1121 578
rect 1177 522 1201 578
rect 1257 522 1301 578
rect 1001 -514 1301 522
rect 1001 -570 1041 -514
rect 1097 -570 1121 -514
rect 1177 -570 1201 -514
rect 1257 -570 1301 -514
rect 1001 -1881 1301 -570
rect 1001 -1937 1041 -1881
rect 1097 -1937 1121 -1881
rect 1177 -1937 1201 -1881
rect 1257 -1937 1301 -1881
rect 1001 -3385 1301 -1937
rect 1001 -3441 1041 -3385
rect 1097 -3441 1121 -3385
rect 1177 -3441 1201 -3385
rect 1257 -3441 1301 -3385
rect 1001 -4889 1301 -3441
rect 1001 -4945 1041 -4889
rect 1097 -4945 1121 -4889
rect 1177 -4945 1201 -4889
rect 1257 -4945 1301 -4889
rect 1001 -4985 1301 -4945
rect 2241 4000 2541 5278
rect 2241 3944 2281 4000
rect 2337 3944 2361 4000
rect 2417 3944 2441 4000
rect 2497 3944 2541 4000
rect 2241 3830 2541 3944
rect 2241 3774 2281 3830
rect 2337 3774 2361 3830
rect 2417 3774 2441 3830
rect 2497 3774 2541 3830
rect 2241 2496 2541 3774
rect 2241 2440 2281 2496
rect 2337 2440 2361 2496
rect 2417 2440 2441 2496
rect 2497 2440 2541 2496
rect 2241 2316 2541 2440
rect 2241 2260 2281 2316
rect 2337 2260 2361 2316
rect 2417 2260 2441 2316
rect 2497 2260 2541 2316
rect 2241 1498 2541 2260
rect 2241 1442 2281 1498
rect 2337 1442 2361 1498
rect 2417 1442 2441 1498
rect 2497 1442 2541 1498
rect 2241 1129 2541 1442
rect 2241 1073 2281 1129
rect 2337 1073 2361 1129
rect 2417 1073 2441 1129
rect 2497 1073 2541 1129
rect 2241 949 2541 1073
rect 2241 893 2281 949
rect 2337 893 2361 949
rect 2417 893 2441 949
rect 2497 893 2541 949
rect 2241 411 2541 893
rect 2241 355 2281 411
rect 2337 355 2361 411
rect 2417 355 2441 411
rect 2497 355 2541 411
rect 2241 35 2541 355
rect 2241 -21 2281 35
rect 2337 -21 2361 35
rect 2417 -21 2441 35
rect 2497 -21 2541 35
rect 2241 -146 2541 -21
rect 2241 -202 2281 -146
rect 2337 -202 2361 -146
rect 2417 -202 2441 -146
rect 2497 -202 2541 -146
rect 2241 -684 2541 -202
rect 2241 -740 2281 -684
rect 2337 -740 2361 -684
rect 2417 -740 2441 -684
rect 2497 -740 2541 -684
rect 2241 -1057 2541 -740
rect 2241 -1113 2281 -1057
rect 2337 -1113 2361 -1057
rect 2417 -1113 2441 -1057
rect 2497 -1113 2541 -1057
rect 2241 -1227 2541 -1113
rect 2241 -1283 2281 -1227
rect 2337 -1283 2361 -1227
rect 2417 -1283 2441 -1227
rect 2497 -1283 2541 -1227
rect 2241 -2561 2541 -1283
rect 2241 -2617 2281 -2561
rect 2337 -2617 2361 -2561
rect 2417 -2617 2441 -2561
rect 2497 -2617 2541 -2561
rect 2241 -2731 2541 -2617
rect 2241 -2787 2281 -2731
rect 2337 -2787 2361 -2731
rect 2417 -2787 2441 -2731
rect 2497 -2787 2541 -2731
rect 2241 -4065 2541 -2787
rect 2241 -4121 2281 -4065
rect 2337 -4121 2361 -4065
rect 2417 -4121 2441 -4065
rect 2497 -4121 2541 -4065
rect 2241 -4235 2541 -4121
rect 2241 -4291 2281 -4235
rect 2337 -4291 2361 -4235
rect 2417 -4291 2441 -4235
rect 2497 -4291 2541 -4235
rect 2241 -5031 2541 -4291
rect 3986 4802 4286 5379
rect 3986 4746 4026 4802
rect 4082 4746 4106 4802
rect 4162 4746 4186 4802
rect 4242 4746 4286 4802
rect 3986 4371 4286 4746
rect 3986 4315 4026 4371
rect 4082 4315 4106 4371
rect 4162 4315 4186 4371
rect 4242 4315 4286 4371
rect 3986 3298 4286 4315
rect 3986 3242 4026 3298
rect 4082 3242 4106 3298
rect 4162 3242 4186 3298
rect 4242 3242 4286 3298
rect 3986 2867 4286 3242
rect 3986 2811 4026 2867
rect 4082 2811 4106 2867
rect 4162 2811 4186 2867
rect 4242 2811 4286 2867
rect 3986 1807 4286 2811
rect 3986 1751 4026 1807
rect 4082 1751 4106 1807
rect 4162 1751 4186 1807
rect 4242 1751 4286 1807
rect 3986 -1602 4286 1751
rect 3986 -1658 4026 -1602
rect 4082 -1658 4106 -1602
rect 4162 -1658 4186 -1602
rect 4242 -1658 4286 -1602
rect 3986 -2038 4286 -1658
rect 3986 -2094 4026 -2038
rect 4082 -2094 4106 -2038
rect 4162 -2094 4186 -2038
rect 4242 -2094 4286 -2038
rect 3986 -3106 4286 -2094
rect 3986 -3162 4026 -3106
rect 4082 -3162 4106 -3106
rect 4162 -3162 4186 -3106
rect 4242 -3162 4286 -3106
rect 3986 -3542 4286 -3162
rect 3986 -3598 4026 -3542
rect 4082 -3598 4106 -3542
rect 4162 -3598 4186 -3542
rect 4242 -3598 4286 -3542
rect 3986 -4610 4286 -3598
rect 3986 -4666 4026 -4610
rect 4082 -4666 4106 -4610
rect 4162 -4666 4186 -4610
rect 4242 -4666 4286 -4610
rect 3986 -5043 4286 -4666
rect 5204 4959 5504 5380
rect 5204 4903 5244 4959
rect 5300 4903 5324 4959
rect 5380 4903 5404 4959
rect 5460 4903 5504 4959
rect 5204 4523 5504 4903
rect 5204 4467 5244 4523
rect 5300 4467 5324 4523
rect 5380 4467 5404 4523
rect 5460 4467 5504 4523
rect 5204 3455 5504 4467
rect 5204 3399 5244 3455
rect 5300 3399 5324 3455
rect 5380 3399 5404 3455
rect 5460 3399 5504 3455
rect 5204 3019 5504 3399
rect 5204 2963 5244 3019
rect 5300 2963 5324 3019
rect 5380 2963 5404 3019
rect 5460 2963 5504 3019
rect 5204 1947 5504 2963
rect 5204 1891 5244 1947
rect 5300 1891 5324 1947
rect 5380 1891 5404 1947
rect 5460 1891 5504 1947
rect 5204 -1750 5504 1891
rect 5204 -1806 5244 -1750
rect 5300 -1806 5324 -1750
rect 5380 -1806 5404 -1750
rect 5460 -1806 5504 -1750
rect 5204 -2190 5504 -1806
rect 5204 -2246 5244 -2190
rect 5300 -2246 5324 -2190
rect 5380 -2246 5404 -2190
rect 5460 -2246 5504 -2190
rect 5204 -3246 5504 -2246
rect 5204 -3302 5244 -3246
rect 5300 -3302 5324 -3246
rect 5380 -3302 5404 -3246
rect 5460 -3302 5504 -3246
rect 5204 -3694 5504 -3302
rect 5204 -3750 5244 -3694
rect 5300 -3750 5324 -3694
rect 5380 -3750 5404 -3694
rect 5460 -3750 5504 -3694
rect 5204 -4767 5504 -3750
rect 5204 -4823 5244 -4767
rect 5300 -4823 5324 -4767
rect 5380 -4823 5404 -4767
rect 5460 -4823 5504 -4767
rect 5204 -5038 5504 -4823
use pfet_2series  pfet_2series_0
timestamp 1698888477
transform 1 0 1107 0 1 -86
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_1
timestamp 1698888477
transform 1 0 1107 0 -1 -1171
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_2
timestamp 1698888477
transform 1 0 -119 0 -1 -1171
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_3
timestamp 1698888477
transform 1 0 591 0 1 -86
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_4
timestamp 1698888477
transform 1 0 591 0 1 -3096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_5
timestamp 1698888477
transform 1 0 -119 0 -1 -5265
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_6
timestamp 1698888477
transform 1 0 1107 0 -1 -5265
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_7
timestamp 1698888477
transform 1 0 591 0 -1 -5265
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_8
timestamp 1698888477
transform 1 0 -119 0 -1 -2257
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_9
timestamp 1698888477
transform 1 0 591 0 -1 -2257
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_10
timestamp 1698888477
transform 1 0 591 0 1 -1592
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_11
timestamp 1698888477
transform 1 0 1107 0 1 -1592
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_12
timestamp 1698888477
transform 1 0 1107 0 1 -3096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_13
timestamp 1698888477
transform 1 0 -119 0 1 -3096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_14
timestamp 1698888477
transform 1 0 1107 0 -1 -3761
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_15
timestamp 1698888477
transform 1 0 -119 0 -1 -3761
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_16
timestamp 1698888477
transform 1 0 591 0 -1 -3761
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_17
timestamp 1698888477
transform 1 0 -119 0 1 -1592
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_18
timestamp 1698888477
transform 1 0 -119 0 1 -86
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_19
timestamp 1698888477
transform 1 0 1107 0 -1 -2257
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_20
timestamp 1698888477
transform 1 0 591 0 -1 -1171
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_21
timestamp 1698888477
transform 1 0 -2377 0 -1 -1171
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_22
timestamp 1698888477
transform 1 0 -1151 0 1 -1592
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_23
timestamp 1698888477
transform 1 0 -1151 0 -1 -3761
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_24
timestamp 1698888477
transform 1 0 -2377 0 1 -3096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_25
timestamp 1698888477
transform 1 0 -1151 0 1 -3096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_26
timestamp 1698888477
transform 1 0 -1861 0 1 -86
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_27
timestamp 1698888477
transform 1 0 -2377 0 1 -86
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_28
timestamp 1698888477
transform 1 0 -1861 0 -1 -5265
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_29
timestamp 1698888477
transform 1 0 -1151 0 -1 -1171
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_30
timestamp 1698888477
transform 1 0 -1861 0 1 -1592
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_31
timestamp 1698888477
transform 1 0 -1151 0 -1 -5265
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_32
timestamp 1698888477
transform 1 0 -1861 0 1 -3096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_33
timestamp 1698888477
transform 1 0 -2377 0 -1 -5265
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_34
timestamp 1698888477
transform 1 0 -1151 0 1 -86
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_35
timestamp 1698888477
transform 1 0 -2377 0 -1 -3761
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_36
timestamp 1698888477
transform 1 0 -1151 0 -1 -2257
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_37
timestamp 1698888477
transform 1 0 -1861 0 -1 -3761
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_38
timestamp 1698888477
transform 1 0 -1861 0 -1 -1171
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_39
timestamp 1698888477
transform 1 0 -2377 0 -1 -2257
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_40
timestamp 1698888477
transform 1 0 -1861 0 -1 -2257
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_41
timestamp 1698888477
transform 1 0 -2377 0 1 -1592
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_42
timestamp 1698888477
transform 1 0 -2377 0 -1 2800
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_43
timestamp 1698888477
transform 1 0 -1861 0 -1 2800
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_44
timestamp 1698888477
transform 1 0 -1151 0 -1 1292
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_45
timestamp 1698888477
transform 1 0 -1151 0 1 3465
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_46
timestamp 1698888477
transform 1 0 -1861 0 1 2096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_47
timestamp 1698888477
transform 1 0 -1861 0 -1 -77
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_48
timestamp 1698888477
transform 1 0 -2377 0 -1 1292
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_49
timestamp 1698888477
transform 1 0 -1861 0 -1 1292
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_50
timestamp 1698888477
transform 1 0 -1861 0 1 3465
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_51
timestamp 1698888477
transform 1 0 -2377 0 1 3465
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_52
timestamp 1698888477
transform 1 0 -1151 0 1 2096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_53
timestamp 1698888477
transform 1 0 -2377 0 -1 -77
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_54
timestamp 1698888477
transform 1 0 -1151 0 -1 -77
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_55
timestamp 1698888477
transform 1 0 -2377 0 1 4969
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_56
timestamp 1698888477
transform 1 0 -1151 0 -1 2800
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_57
timestamp 1698888477
transform 1 0 -1861 0 1 4969
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_58
timestamp 1698888477
transform 1 0 -2377 0 1 2096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_59
timestamp 1698888477
transform 1 0 -1151 0 1 4969
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_60
timestamp 1698888477
transform 1 0 -1861 0 -1 4304
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_61
timestamp 1698888477
transform 1 0 -1151 0 -1 4304
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_62
timestamp 1698888477
transform 1 0 -2377 0 -1 4304
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_63
timestamp 1698888477
transform 1 0 1107 0 -1 2800
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_64
timestamp 1698888477
transform 1 0 -119 0 -1 4304
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_65
timestamp 1698888477
transform 1 0 591 0 -1 2800
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_66
timestamp 1698888477
transform 1 0 -119 0 -1 1292
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_67
timestamp 1698888477
transform 1 0 591 0 -1 1292
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_68
timestamp 1698888477
transform 1 0 591 0 1 3465
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_69
timestamp 1698888477
transform 1 0 -119 0 1 4969
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_70
timestamp 1698888477
transform 1 0 1107 0 -1 1292
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_71
timestamp 1698888477
transform 1 0 591 0 -1 4304
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_72
timestamp 1698888477
transform 1 0 -119 0 1 2096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_73
timestamp 1698888477
transform 1 0 591 0 -1 -77
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_74
timestamp 1698888477
transform 1 0 1107 0 1 2096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_75
timestamp 1698888477
transform 1 0 591 0 1 4969
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_76
timestamp 1698888477
transform 1 0 1107 0 1 4969
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_77
timestamp 1698888477
transform 1 0 1107 0 -1 -77
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_78
timestamp 1698888477
transform 1 0 591 0 1 2096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_79
timestamp 1698888477
transform 1 0 1107 0 1 3465
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_80
timestamp 1698888477
transform 1 0 -119 0 1 3465
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_81
timestamp 1698888477
transform 1 0 1107 0 -1 4304
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_82
timestamp 1698888477
transform 1 0 -119 0 -1 -77
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_83
timestamp 1698888477
transform 1 0 -119 0 -1 2800
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_84
timestamp 1698888477
transform 1 0 -635 0 1 4969
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_85
timestamp 1698888477
transform 1 0 -635 0 -1 -5265
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_86
timestamp 1698888477
transform 1 0 -635 0 -1 -2257
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_87
timestamp 1698888477
transform 1 0 -635 0 1 -1592
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_88
timestamp 1698888477
transform 1 0 -635 0 -1 -3761
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_89
timestamp 1698888477
transform 1 0 -635 0 1 -3096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_90
timestamp 1698888477
transform 1 0 -635 0 1 -86
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_91
timestamp 1698888477
transform 1 0 -635 0 1 1010
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_92
timestamp 1698888477
transform 1 0 -635 0 -1 4304
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_93
timestamp 1698888477
transform 1 0 -2377 0 1 1010
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_94
timestamp 1698888477
transform 1 0 -635 0 -1 2800
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_95
timestamp 1698888477
transform 1 0 -635 0 -1 1292
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_96
timestamp 1698888477
transform 1 0 -635 0 1 3465
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_97
timestamp 1698888477
transform 1 0 -635 0 -1 -1171
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_98
timestamp 1698888477
transform 1 0 1107 0 1 1010
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_99
timestamp 1698888477
transform 1 0 -1151 0 1 1010
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_100
timestamp 1698888477
transform 1 0 -119 0 1 1010
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_101
timestamp 1698888477
transform 1 0 591 0 1 1010
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_102
timestamp 1698888477
transform 1 0 -1861 0 1 1010
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_103
timestamp 1698888477
transform 1 0 -635 0 1 2096
box 3549 -998 4227 -608
use pfet_2series  pfet_2series_104
timestamp 1698888477
transform 1 0 -635 0 -1 -77
box 3549 -998 4227 -608
<< labels >>
flabel metal3 s 4002 -2148 4248 -1692 2 FreeSans 3126 0 0 0 VB3
port 1 nsew
flabel metal3 s 5220 -2142 5466 -1716 2 FreeSans 3126 0 0 0 VB2
port 2 nsew
flabel metal3 s 1028 -2329 1267 -1449 2 FreeSans 3126 0 0 0 AVDD
port 3 nsew
flabel metal3 s 2273 -2106 2511 -1710 2 FreeSans 3126 0 0 0 VB1
port 4 nsew
<< end >>
