magic
tech sky130A
magscale 1 2
timestamp 1698710451
<< pwell >>
rect -270 592 6894 1015
rect -270 398 -184 592
rect 3269 398 3355 592
rect 6808 398 6894 592
rect -270 312 6894 398
rect -270 118 -184 312
rect 3269 118 3355 312
rect 6808 118 6894 312
rect -270 -134 6894 118
rect -270 -555 -184 -134
rect 3269 -555 3355 -134
rect 6808 -555 6894 -134
rect -270 -807 6894 -555
rect -270 -1000 -184 -807
rect 3269 -1000 3355 -807
rect 6808 -1000 6894 -807
rect -270 -1086 6894 -1000
rect -270 -1279 -184 -1086
rect 3269 -1279 3355 -1086
rect 6808 -1279 6894 -1086
rect -270 -1531 6894 -1279
rect -270 -1952 -184 -1531
rect 3269 -1952 3355 -1531
rect 6808 -1952 6894 -1531
rect -270 -2204 6894 -1952
rect -270 -2398 -184 -2204
rect 3269 -2398 3355 -2204
rect 6808 -2398 6894 -2204
rect -270 -2484 6894 -2398
rect -270 -2678 -184 -2484
rect 3269 -2678 3355 -2484
rect 6808 -2678 6894 -2484
rect -270 -3101 6894 -2678
<< nmos >>
rect -84 618 116 818
rect 421 618 621 818
rect 679 618 879 818
rect 1184 618 1384 818
rect 1442 618 1642 818
rect 1700 618 1900 818
rect 2205 618 2405 818
rect 2463 618 2663 818
rect 2969 618 3169 818
rect 3455 618 3655 818
rect 3961 618 4161 818
rect 4219 618 4419 818
rect 4724 618 4924 818
rect 4982 618 5182 818
rect 5240 618 5440 818
rect 5745 618 5945 818
rect 6003 618 6203 818
rect 6508 618 6708 818
rect -84 -108 116 92
rect 421 -108 621 92
rect 679 -108 879 92
rect 1184 -108 1384 92
rect 1442 -108 1642 92
rect 1700 -108 1900 92
rect 2205 -108 2405 92
rect 2463 -108 2663 92
rect 2969 -108 3169 92
rect 3455 -108 3655 92
rect 3961 -108 4161 92
rect 4219 -108 4419 92
rect 4724 -108 4924 92
rect 4982 -108 5182 92
rect 5240 -108 5440 92
rect 5745 -108 5945 92
rect 6003 -108 6203 92
rect 6508 -108 6708 92
rect -84 -781 116 -581
rect 421 -781 621 -581
rect 679 -781 879 -581
rect 1184 -781 1384 -581
rect 1442 -781 1642 -581
rect 1700 -781 1900 -581
rect 2205 -781 2405 -581
rect 2463 -781 2663 -581
rect 2969 -781 3169 -581
rect 3455 -781 3655 -581
rect 3961 -781 4161 -581
rect 4219 -781 4419 -581
rect 4724 -781 4924 -581
rect 4982 -781 5182 -581
rect 5240 -781 5440 -581
rect 5745 -781 5945 -581
rect 6003 -781 6203 -581
rect 6508 -781 6708 -581
rect -84 -1505 116 -1305
rect 421 -1505 621 -1305
rect 679 -1505 879 -1305
rect 1184 -1505 1384 -1305
rect 1442 -1505 1642 -1305
rect 1700 -1505 1900 -1305
rect 2205 -1505 2405 -1305
rect 2463 -1505 2663 -1305
rect 2969 -1505 3169 -1305
rect 3455 -1505 3655 -1305
rect 3961 -1505 4161 -1305
rect 4219 -1505 4419 -1305
rect 4724 -1505 4924 -1305
rect 4982 -1505 5182 -1305
rect 5240 -1505 5440 -1305
rect 5745 -1505 5945 -1305
rect 6003 -1505 6203 -1305
rect 6508 -1505 6708 -1305
rect -84 -2178 116 -1978
rect 421 -2178 621 -1978
rect 679 -2178 879 -1978
rect 1184 -2178 1384 -1978
rect 1442 -2178 1642 -1978
rect 1700 -2178 1900 -1978
rect 2205 -2178 2405 -1978
rect 2463 -2178 2663 -1978
rect 2969 -2178 3169 -1978
rect 3455 -2178 3655 -1978
rect 3961 -2178 4161 -1978
rect 4219 -2178 4419 -1978
rect 4724 -2178 4924 -1978
rect 4982 -2178 5182 -1978
rect 5240 -2178 5440 -1978
rect 5745 -2178 5945 -1978
rect 6003 -2178 6203 -1978
rect 6508 -2178 6708 -1978
rect -84 -2904 116 -2704
rect 421 -2904 621 -2704
rect 679 -2904 879 -2704
rect 1184 -2904 1384 -2704
rect 1442 -2904 1642 -2704
rect 1700 -2904 1900 -2704
rect 2205 -2904 2405 -2704
rect 2463 -2904 2663 -2704
rect 2969 -2904 3169 -2704
rect 3455 -2904 3655 -2704
rect 3961 -2904 4161 -2704
rect 4219 -2904 4419 -2704
rect 4724 -2904 4924 -2704
rect 4982 -2904 5182 -2704
rect 5240 -2904 5440 -2704
rect 5745 -2904 5945 -2704
rect 6003 -2904 6203 -2704
rect 6508 -2904 6708 -2704
<< ndiff >>
rect -142 803 -84 818
rect -142 769 -130 803
rect -96 769 -84 803
rect -142 735 -84 769
rect -142 701 -130 735
rect -96 701 -84 735
rect -142 667 -84 701
rect -142 633 -130 667
rect -96 633 -84 667
rect -142 618 -84 633
rect 116 803 174 818
rect 116 769 128 803
rect 162 769 174 803
rect 116 735 174 769
rect 116 701 128 735
rect 162 701 174 735
rect 116 667 174 701
rect 116 633 128 667
rect 162 633 174 667
rect 116 618 174 633
rect 363 803 421 818
rect 363 769 375 803
rect 409 769 421 803
rect 363 735 421 769
rect 363 701 375 735
rect 409 701 421 735
rect 363 667 421 701
rect 363 633 375 667
rect 409 633 421 667
rect 363 618 421 633
rect 621 803 679 818
rect 621 769 633 803
rect 667 769 679 803
rect 621 735 679 769
rect 621 701 633 735
rect 667 701 679 735
rect 621 667 679 701
rect 621 633 633 667
rect 667 633 679 667
rect 621 618 679 633
rect 879 803 937 818
rect 879 769 891 803
rect 925 769 937 803
rect 879 735 937 769
rect 879 701 891 735
rect 925 701 937 735
rect 879 667 937 701
rect 879 633 891 667
rect 925 633 937 667
rect 879 618 937 633
rect 1126 803 1184 818
rect 1126 769 1138 803
rect 1172 769 1184 803
rect 1126 735 1184 769
rect 1126 701 1138 735
rect 1172 701 1184 735
rect 1126 667 1184 701
rect 1126 633 1138 667
rect 1172 633 1184 667
rect 1126 618 1184 633
rect 1384 803 1442 818
rect 1384 769 1396 803
rect 1430 769 1442 803
rect 1384 735 1442 769
rect 1384 701 1396 735
rect 1430 701 1442 735
rect 1384 667 1442 701
rect 1384 633 1396 667
rect 1430 633 1442 667
rect 1384 618 1442 633
rect 1642 803 1700 818
rect 1642 769 1654 803
rect 1688 769 1700 803
rect 1642 735 1700 769
rect 1642 701 1654 735
rect 1688 701 1700 735
rect 1642 667 1700 701
rect 1642 633 1654 667
rect 1688 633 1700 667
rect 1642 618 1700 633
rect 1900 803 1958 818
rect 1900 769 1912 803
rect 1946 769 1958 803
rect 1900 735 1958 769
rect 1900 701 1912 735
rect 1946 701 1958 735
rect 1900 667 1958 701
rect 1900 633 1912 667
rect 1946 633 1958 667
rect 1900 618 1958 633
rect 2147 803 2205 818
rect 2147 769 2159 803
rect 2193 769 2205 803
rect 2147 735 2205 769
rect 2147 701 2159 735
rect 2193 701 2205 735
rect 2147 667 2205 701
rect 2147 633 2159 667
rect 2193 633 2205 667
rect 2147 618 2205 633
rect 2405 803 2463 818
rect 2405 769 2417 803
rect 2451 769 2463 803
rect 2405 735 2463 769
rect 2405 701 2417 735
rect 2451 701 2463 735
rect 2405 667 2463 701
rect 2405 633 2417 667
rect 2451 633 2463 667
rect 2405 618 2463 633
rect 2663 803 2721 818
rect 2663 769 2675 803
rect 2709 769 2721 803
rect 2663 735 2721 769
rect 2663 701 2675 735
rect 2709 701 2721 735
rect 2663 667 2721 701
rect 2663 633 2675 667
rect 2709 633 2721 667
rect 2663 618 2721 633
rect 2911 803 2969 818
rect 2911 769 2923 803
rect 2957 769 2969 803
rect 2911 735 2969 769
rect 2911 701 2923 735
rect 2957 701 2969 735
rect 2911 667 2969 701
rect 2911 633 2923 667
rect 2957 633 2969 667
rect 2911 618 2969 633
rect 3169 803 3227 818
rect 3169 769 3181 803
rect 3215 769 3227 803
rect 3169 735 3227 769
rect 3169 701 3181 735
rect 3215 701 3227 735
rect 3169 667 3227 701
rect 3169 633 3181 667
rect 3215 633 3227 667
rect 3169 618 3227 633
rect 3397 803 3455 818
rect 3397 769 3409 803
rect 3443 769 3455 803
rect 3397 735 3455 769
rect 3397 701 3409 735
rect 3443 701 3455 735
rect 3397 667 3455 701
rect 3397 633 3409 667
rect 3443 633 3455 667
rect 3397 618 3455 633
rect 3655 803 3713 818
rect 3655 769 3667 803
rect 3701 769 3713 803
rect 3655 735 3713 769
rect 3655 701 3667 735
rect 3701 701 3713 735
rect 3655 667 3713 701
rect 3655 633 3667 667
rect 3701 633 3713 667
rect 3655 618 3713 633
rect 3903 803 3961 818
rect 3903 769 3915 803
rect 3949 769 3961 803
rect 3903 735 3961 769
rect 3903 701 3915 735
rect 3949 701 3961 735
rect 3903 667 3961 701
rect 3903 633 3915 667
rect 3949 633 3961 667
rect 3903 618 3961 633
rect 4161 803 4219 818
rect 4161 769 4173 803
rect 4207 769 4219 803
rect 4161 735 4219 769
rect 4161 701 4173 735
rect 4207 701 4219 735
rect 4161 667 4219 701
rect 4161 633 4173 667
rect 4207 633 4219 667
rect 4161 618 4219 633
rect 4419 803 4477 818
rect 4419 769 4431 803
rect 4465 769 4477 803
rect 4419 735 4477 769
rect 4419 701 4431 735
rect 4465 701 4477 735
rect 4419 667 4477 701
rect 4419 633 4431 667
rect 4465 633 4477 667
rect 4419 618 4477 633
rect 4666 803 4724 818
rect 4666 769 4678 803
rect 4712 769 4724 803
rect 4666 735 4724 769
rect 4666 701 4678 735
rect 4712 701 4724 735
rect 4666 667 4724 701
rect 4666 633 4678 667
rect 4712 633 4724 667
rect 4666 618 4724 633
rect 4924 803 4982 818
rect 4924 769 4936 803
rect 4970 769 4982 803
rect 4924 735 4982 769
rect 4924 701 4936 735
rect 4970 701 4982 735
rect 4924 667 4982 701
rect 4924 633 4936 667
rect 4970 633 4982 667
rect 4924 618 4982 633
rect 5182 803 5240 818
rect 5182 769 5194 803
rect 5228 769 5240 803
rect 5182 735 5240 769
rect 5182 701 5194 735
rect 5228 701 5240 735
rect 5182 667 5240 701
rect 5182 633 5194 667
rect 5228 633 5240 667
rect 5182 618 5240 633
rect 5440 803 5498 818
rect 5440 769 5452 803
rect 5486 769 5498 803
rect 5440 735 5498 769
rect 5440 701 5452 735
rect 5486 701 5498 735
rect 5440 667 5498 701
rect 5440 633 5452 667
rect 5486 633 5498 667
rect 5440 618 5498 633
rect 5687 803 5745 818
rect 5687 769 5699 803
rect 5733 769 5745 803
rect 5687 735 5745 769
rect 5687 701 5699 735
rect 5733 701 5745 735
rect 5687 667 5745 701
rect 5687 633 5699 667
rect 5733 633 5745 667
rect 5687 618 5745 633
rect 5945 803 6003 818
rect 5945 769 5957 803
rect 5991 769 6003 803
rect 5945 735 6003 769
rect 5945 701 5957 735
rect 5991 701 6003 735
rect 5945 667 6003 701
rect 5945 633 5957 667
rect 5991 633 6003 667
rect 5945 618 6003 633
rect 6203 803 6261 818
rect 6203 769 6215 803
rect 6249 769 6261 803
rect 6203 735 6261 769
rect 6203 701 6215 735
rect 6249 701 6261 735
rect 6203 667 6261 701
rect 6203 633 6215 667
rect 6249 633 6261 667
rect 6203 618 6261 633
rect 6450 803 6508 818
rect 6450 769 6462 803
rect 6496 769 6508 803
rect 6450 735 6508 769
rect 6450 701 6462 735
rect 6496 701 6508 735
rect 6450 667 6508 701
rect 6450 633 6462 667
rect 6496 633 6508 667
rect 6450 618 6508 633
rect 6708 803 6766 818
rect 6708 769 6720 803
rect 6754 769 6766 803
rect 6708 735 6766 769
rect 6708 701 6720 735
rect 6754 701 6766 735
rect 6708 667 6766 701
rect 6708 633 6720 667
rect 6754 633 6766 667
rect 6708 618 6766 633
rect -142 77 -84 92
rect -142 43 -130 77
rect -96 43 -84 77
rect -142 9 -84 43
rect -142 -25 -130 9
rect -96 -25 -84 9
rect -142 -59 -84 -25
rect -142 -93 -130 -59
rect -96 -93 -84 -59
rect -142 -108 -84 -93
rect 116 77 174 92
rect 116 43 128 77
rect 162 43 174 77
rect 116 9 174 43
rect 116 -25 128 9
rect 162 -25 174 9
rect 116 -59 174 -25
rect 116 -93 128 -59
rect 162 -93 174 -59
rect 116 -108 174 -93
rect 363 77 421 92
rect 363 43 375 77
rect 409 43 421 77
rect 363 9 421 43
rect 363 -25 375 9
rect 409 -25 421 9
rect 363 -59 421 -25
rect 363 -93 375 -59
rect 409 -93 421 -59
rect 363 -108 421 -93
rect 621 77 679 92
rect 621 43 633 77
rect 667 43 679 77
rect 621 9 679 43
rect 621 -25 633 9
rect 667 -25 679 9
rect 621 -59 679 -25
rect 621 -93 633 -59
rect 667 -93 679 -59
rect 621 -108 679 -93
rect 879 77 937 92
rect 879 43 891 77
rect 925 43 937 77
rect 879 9 937 43
rect 879 -25 891 9
rect 925 -25 937 9
rect 879 -59 937 -25
rect 879 -93 891 -59
rect 925 -93 937 -59
rect 879 -108 937 -93
rect 1126 77 1184 92
rect 1126 43 1138 77
rect 1172 43 1184 77
rect 1126 9 1184 43
rect 1126 -25 1138 9
rect 1172 -25 1184 9
rect 1126 -59 1184 -25
rect 1126 -93 1138 -59
rect 1172 -93 1184 -59
rect 1126 -108 1184 -93
rect 1384 77 1442 92
rect 1384 43 1396 77
rect 1430 43 1442 77
rect 1384 9 1442 43
rect 1384 -25 1396 9
rect 1430 -25 1442 9
rect 1384 -59 1442 -25
rect 1384 -93 1396 -59
rect 1430 -93 1442 -59
rect 1384 -108 1442 -93
rect 1642 77 1700 92
rect 1642 43 1654 77
rect 1688 43 1700 77
rect 1642 9 1700 43
rect 1642 -25 1654 9
rect 1688 -25 1700 9
rect 1642 -59 1700 -25
rect 1642 -93 1654 -59
rect 1688 -93 1700 -59
rect 1642 -108 1700 -93
rect 1900 77 1958 92
rect 1900 43 1912 77
rect 1946 43 1958 77
rect 1900 9 1958 43
rect 1900 -25 1912 9
rect 1946 -25 1958 9
rect 1900 -59 1958 -25
rect 1900 -93 1912 -59
rect 1946 -93 1958 -59
rect 1900 -108 1958 -93
rect 2147 77 2205 92
rect 2147 43 2159 77
rect 2193 43 2205 77
rect 2147 9 2205 43
rect 2147 -25 2159 9
rect 2193 -25 2205 9
rect 2147 -59 2205 -25
rect 2147 -93 2159 -59
rect 2193 -93 2205 -59
rect 2147 -108 2205 -93
rect 2405 77 2463 92
rect 2405 43 2417 77
rect 2451 43 2463 77
rect 2405 9 2463 43
rect 2405 -25 2417 9
rect 2451 -25 2463 9
rect 2405 -59 2463 -25
rect 2405 -93 2417 -59
rect 2451 -93 2463 -59
rect 2405 -108 2463 -93
rect 2663 77 2721 92
rect 2663 43 2675 77
rect 2709 43 2721 77
rect 2663 9 2721 43
rect 2663 -25 2675 9
rect 2709 -25 2721 9
rect 2663 -59 2721 -25
rect 2663 -93 2675 -59
rect 2709 -93 2721 -59
rect 2663 -108 2721 -93
rect 2911 77 2969 92
rect 2911 43 2923 77
rect 2957 43 2969 77
rect 2911 9 2969 43
rect 2911 -25 2923 9
rect 2957 -25 2969 9
rect 2911 -59 2969 -25
rect 2911 -93 2923 -59
rect 2957 -93 2969 -59
rect 2911 -108 2969 -93
rect 3169 77 3227 92
rect 3169 43 3181 77
rect 3215 43 3227 77
rect 3169 9 3227 43
rect 3169 -25 3181 9
rect 3215 -25 3227 9
rect 3169 -59 3227 -25
rect 3169 -93 3181 -59
rect 3215 -93 3227 -59
rect 3169 -108 3227 -93
rect 3397 77 3455 92
rect 3397 43 3409 77
rect 3443 43 3455 77
rect 3397 9 3455 43
rect 3397 -25 3409 9
rect 3443 -25 3455 9
rect 3397 -59 3455 -25
rect 3397 -93 3409 -59
rect 3443 -93 3455 -59
rect 3397 -108 3455 -93
rect 3655 77 3713 92
rect 3655 43 3667 77
rect 3701 43 3713 77
rect 3655 9 3713 43
rect 3655 -25 3667 9
rect 3701 -25 3713 9
rect 3655 -59 3713 -25
rect 3655 -93 3667 -59
rect 3701 -93 3713 -59
rect 3655 -108 3713 -93
rect 3903 77 3961 92
rect 3903 43 3915 77
rect 3949 43 3961 77
rect 3903 9 3961 43
rect 3903 -25 3915 9
rect 3949 -25 3961 9
rect 3903 -59 3961 -25
rect 3903 -93 3915 -59
rect 3949 -93 3961 -59
rect 3903 -108 3961 -93
rect 4161 77 4219 92
rect 4161 43 4173 77
rect 4207 43 4219 77
rect 4161 9 4219 43
rect 4161 -25 4173 9
rect 4207 -25 4219 9
rect 4161 -59 4219 -25
rect 4161 -93 4173 -59
rect 4207 -93 4219 -59
rect 4161 -108 4219 -93
rect 4419 77 4477 92
rect 4419 43 4431 77
rect 4465 43 4477 77
rect 4419 9 4477 43
rect 4419 -25 4431 9
rect 4465 -25 4477 9
rect 4419 -59 4477 -25
rect 4419 -93 4431 -59
rect 4465 -93 4477 -59
rect 4419 -108 4477 -93
rect 4666 77 4724 92
rect 4666 43 4678 77
rect 4712 43 4724 77
rect 4666 9 4724 43
rect 4666 -25 4678 9
rect 4712 -25 4724 9
rect 4666 -59 4724 -25
rect 4666 -93 4678 -59
rect 4712 -93 4724 -59
rect 4666 -108 4724 -93
rect 4924 77 4982 92
rect 4924 43 4936 77
rect 4970 43 4982 77
rect 4924 9 4982 43
rect 4924 -25 4936 9
rect 4970 -25 4982 9
rect 4924 -59 4982 -25
rect 4924 -93 4936 -59
rect 4970 -93 4982 -59
rect 4924 -108 4982 -93
rect 5182 77 5240 92
rect 5182 43 5194 77
rect 5228 43 5240 77
rect 5182 9 5240 43
rect 5182 -25 5194 9
rect 5228 -25 5240 9
rect 5182 -59 5240 -25
rect 5182 -93 5194 -59
rect 5228 -93 5240 -59
rect 5182 -108 5240 -93
rect 5440 77 5498 92
rect 5440 43 5452 77
rect 5486 43 5498 77
rect 5440 9 5498 43
rect 5440 -25 5452 9
rect 5486 -25 5498 9
rect 5440 -59 5498 -25
rect 5440 -93 5452 -59
rect 5486 -93 5498 -59
rect 5440 -108 5498 -93
rect 5687 77 5745 92
rect 5687 43 5699 77
rect 5733 43 5745 77
rect 5687 9 5745 43
rect 5687 -25 5699 9
rect 5733 -25 5745 9
rect 5687 -59 5745 -25
rect 5687 -93 5699 -59
rect 5733 -93 5745 -59
rect 5687 -108 5745 -93
rect 5945 77 6003 92
rect 5945 43 5957 77
rect 5991 43 6003 77
rect 5945 9 6003 43
rect 5945 -25 5957 9
rect 5991 -25 6003 9
rect 5945 -59 6003 -25
rect 5945 -93 5957 -59
rect 5991 -93 6003 -59
rect 5945 -108 6003 -93
rect 6203 77 6261 92
rect 6203 43 6215 77
rect 6249 43 6261 77
rect 6203 9 6261 43
rect 6203 -25 6215 9
rect 6249 -25 6261 9
rect 6203 -59 6261 -25
rect 6203 -93 6215 -59
rect 6249 -93 6261 -59
rect 6203 -108 6261 -93
rect 6450 77 6508 92
rect 6450 43 6462 77
rect 6496 43 6508 77
rect 6450 9 6508 43
rect 6450 -25 6462 9
rect 6496 -25 6508 9
rect 6450 -59 6508 -25
rect 6450 -93 6462 -59
rect 6496 -93 6508 -59
rect 6450 -108 6508 -93
rect 6708 77 6766 92
rect 6708 43 6720 77
rect 6754 43 6766 77
rect 6708 9 6766 43
rect 6708 -25 6720 9
rect 6754 -25 6766 9
rect 6708 -59 6766 -25
rect 6708 -93 6720 -59
rect 6754 -93 6766 -59
rect 6708 -108 6766 -93
rect -142 -596 -84 -581
rect -142 -630 -130 -596
rect -96 -630 -84 -596
rect -142 -664 -84 -630
rect -142 -698 -130 -664
rect -96 -698 -84 -664
rect -142 -732 -84 -698
rect -142 -766 -130 -732
rect -96 -766 -84 -732
rect -142 -781 -84 -766
rect 116 -596 174 -581
rect 116 -630 128 -596
rect 162 -630 174 -596
rect 116 -664 174 -630
rect 116 -698 128 -664
rect 162 -698 174 -664
rect 116 -732 174 -698
rect 116 -766 128 -732
rect 162 -766 174 -732
rect 116 -781 174 -766
rect 363 -596 421 -581
rect 363 -630 375 -596
rect 409 -630 421 -596
rect 363 -664 421 -630
rect 363 -698 375 -664
rect 409 -698 421 -664
rect 363 -732 421 -698
rect 363 -766 375 -732
rect 409 -766 421 -732
rect 363 -781 421 -766
rect 621 -596 679 -581
rect 621 -630 633 -596
rect 667 -630 679 -596
rect 621 -664 679 -630
rect 621 -698 633 -664
rect 667 -698 679 -664
rect 621 -732 679 -698
rect 621 -766 633 -732
rect 667 -766 679 -732
rect 621 -781 679 -766
rect 879 -596 937 -581
rect 879 -630 891 -596
rect 925 -630 937 -596
rect 879 -664 937 -630
rect 879 -698 891 -664
rect 925 -698 937 -664
rect 879 -732 937 -698
rect 879 -766 891 -732
rect 925 -766 937 -732
rect 879 -781 937 -766
rect 1126 -596 1184 -581
rect 1126 -630 1138 -596
rect 1172 -630 1184 -596
rect 1126 -664 1184 -630
rect 1126 -698 1138 -664
rect 1172 -698 1184 -664
rect 1126 -732 1184 -698
rect 1126 -766 1138 -732
rect 1172 -766 1184 -732
rect 1126 -781 1184 -766
rect 1384 -596 1442 -581
rect 1384 -630 1396 -596
rect 1430 -630 1442 -596
rect 1384 -664 1442 -630
rect 1384 -698 1396 -664
rect 1430 -698 1442 -664
rect 1384 -732 1442 -698
rect 1384 -766 1396 -732
rect 1430 -766 1442 -732
rect 1384 -781 1442 -766
rect 1642 -596 1700 -581
rect 1642 -630 1654 -596
rect 1688 -630 1700 -596
rect 1642 -664 1700 -630
rect 1642 -698 1654 -664
rect 1688 -698 1700 -664
rect 1642 -732 1700 -698
rect 1642 -766 1654 -732
rect 1688 -766 1700 -732
rect 1642 -781 1700 -766
rect 1900 -596 1958 -581
rect 1900 -630 1912 -596
rect 1946 -630 1958 -596
rect 1900 -664 1958 -630
rect 1900 -698 1912 -664
rect 1946 -698 1958 -664
rect 1900 -732 1958 -698
rect 1900 -766 1912 -732
rect 1946 -766 1958 -732
rect 1900 -781 1958 -766
rect 2147 -596 2205 -581
rect 2147 -630 2159 -596
rect 2193 -630 2205 -596
rect 2147 -664 2205 -630
rect 2147 -698 2159 -664
rect 2193 -698 2205 -664
rect 2147 -732 2205 -698
rect 2147 -766 2159 -732
rect 2193 -766 2205 -732
rect 2147 -781 2205 -766
rect 2405 -596 2463 -581
rect 2405 -630 2417 -596
rect 2451 -630 2463 -596
rect 2405 -664 2463 -630
rect 2405 -698 2417 -664
rect 2451 -698 2463 -664
rect 2405 -732 2463 -698
rect 2405 -766 2417 -732
rect 2451 -766 2463 -732
rect 2405 -781 2463 -766
rect 2663 -596 2721 -581
rect 2663 -630 2675 -596
rect 2709 -630 2721 -596
rect 2663 -664 2721 -630
rect 2663 -698 2675 -664
rect 2709 -698 2721 -664
rect 2663 -732 2721 -698
rect 2663 -766 2675 -732
rect 2709 -766 2721 -732
rect 2663 -781 2721 -766
rect 2911 -596 2969 -581
rect 2911 -630 2923 -596
rect 2957 -630 2969 -596
rect 2911 -664 2969 -630
rect 2911 -698 2923 -664
rect 2957 -698 2969 -664
rect 2911 -732 2969 -698
rect 2911 -766 2923 -732
rect 2957 -766 2969 -732
rect 2911 -781 2969 -766
rect 3169 -596 3227 -581
rect 3169 -630 3181 -596
rect 3215 -630 3227 -596
rect 3169 -664 3227 -630
rect 3169 -698 3181 -664
rect 3215 -698 3227 -664
rect 3169 -732 3227 -698
rect 3169 -766 3181 -732
rect 3215 -766 3227 -732
rect 3169 -781 3227 -766
rect 3397 -596 3455 -581
rect 3397 -630 3409 -596
rect 3443 -630 3455 -596
rect 3397 -664 3455 -630
rect 3397 -698 3409 -664
rect 3443 -698 3455 -664
rect 3397 -732 3455 -698
rect 3397 -766 3409 -732
rect 3443 -766 3455 -732
rect 3397 -781 3455 -766
rect 3655 -596 3713 -581
rect 3655 -630 3667 -596
rect 3701 -630 3713 -596
rect 3655 -664 3713 -630
rect 3655 -698 3667 -664
rect 3701 -698 3713 -664
rect 3655 -732 3713 -698
rect 3655 -766 3667 -732
rect 3701 -766 3713 -732
rect 3655 -781 3713 -766
rect 3903 -596 3961 -581
rect 3903 -630 3915 -596
rect 3949 -630 3961 -596
rect 3903 -664 3961 -630
rect 3903 -698 3915 -664
rect 3949 -698 3961 -664
rect 3903 -732 3961 -698
rect 3903 -766 3915 -732
rect 3949 -766 3961 -732
rect 3903 -781 3961 -766
rect 4161 -596 4219 -581
rect 4161 -630 4173 -596
rect 4207 -630 4219 -596
rect 4161 -664 4219 -630
rect 4161 -698 4173 -664
rect 4207 -698 4219 -664
rect 4161 -732 4219 -698
rect 4161 -766 4173 -732
rect 4207 -766 4219 -732
rect 4161 -781 4219 -766
rect 4419 -596 4477 -581
rect 4419 -630 4431 -596
rect 4465 -630 4477 -596
rect 4419 -664 4477 -630
rect 4419 -698 4431 -664
rect 4465 -698 4477 -664
rect 4419 -732 4477 -698
rect 4419 -766 4431 -732
rect 4465 -766 4477 -732
rect 4419 -781 4477 -766
rect 4666 -596 4724 -581
rect 4666 -630 4678 -596
rect 4712 -630 4724 -596
rect 4666 -664 4724 -630
rect 4666 -698 4678 -664
rect 4712 -698 4724 -664
rect 4666 -732 4724 -698
rect 4666 -766 4678 -732
rect 4712 -766 4724 -732
rect 4666 -781 4724 -766
rect 4924 -596 4982 -581
rect 4924 -630 4936 -596
rect 4970 -630 4982 -596
rect 4924 -664 4982 -630
rect 4924 -698 4936 -664
rect 4970 -698 4982 -664
rect 4924 -732 4982 -698
rect 4924 -766 4936 -732
rect 4970 -766 4982 -732
rect 4924 -781 4982 -766
rect 5182 -596 5240 -581
rect 5182 -630 5194 -596
rect 5228 -630 5240 -596
rect 5182 -664 5240 -630
rect 5182 -698 5194 -664
rect 5228 -698 5240 -664
rect 5182 -732 5240 -698
rect 5182 -766 5194 -732
rect 5228 -766 5240 -732
rect 5182 -781 5240 -766
rect 5440 -596 5498 -581
rect 5440 -630 5452 -596
rect 5486 -630 5498 -596
rect 5440 -664 5498 -630
rect 5440 -698 5452 -664
rect 5486 -698 5498 -664
rect 5440 -732 5498 -698
rect 5440 -766 5452 -732
rect 5486 -766 5498 -732
rect 5440 -781 5498 -766
rect 5687 -596 5745 -581
rect 5687 -630 5699 -596
rect 5733 -630 5745 -596
rect 5687 -664 5745 -630
rect 5687 -698 5699 -664
rect 5733 -698 5745 -664
rect 5687 -732 5745 -698
rect 5687 -766 5699 -732
rect 5733 -766 5745 -732
rect 5687 -781 5745 -766
rect 5945 -596 6003 -581
rect 5945 -630 5957 -596
rect 5991 -630 6003 -596
rect 5945 -664 6003 -630
rect 5945 -698 5957 -664
rect 5991 -698 6003 -664
rect 5945 -732 6003 -698
rect 5945 -766 5957 -732
rect 5991 -766 6003 -732
rect 5945 -781 6003 -766
rect 6203 -596 6261 -581
rect 6203 -630 6215 -596
rect 6249 -630 6261 -596
rect 6203 -664 6261 -630
rect 6203 -698 6215 -664
rect 6249 -698 6261 -664
rect 6203 -732 6261 -698
rect 6203 -766 6215 -732
rect 6249 -766 6261 -732
rect 6203 -781 6261 -766
rect 6450 -596 6508 -581
rect 6450 -630 6462 -596
rect 6496 -630 6508 -596
rect 6450 -664 6508 -630
rect 6450 -698 6462 -664
rect 6496 -698 6508 -664
rect 6450 -732 6508 -698
rect 6450 -766 6462 -732
rect 6496 -766 6508 -732
rect 6450 -781 6508 -766
rect 6708 -596 6766 -581
rect 6708 -630 6720 -596
rect 6754 -630 6766 -596
rect 6708 -664 6766 -630
rect 6708 -698 6720 -664
rect 6754 -698 6766 -664
rect 6708 -732 6766 -698
rect 6708 -766 6720 -732
rect 6754 -766 6766 -732
rect 6708 -781 6766 -766
rect -142 -1320 -84 -1305
rect -142 -1354 -130 -1320
rect -96 -1354 -84 -1320
rect -142 -1388 -84 -1354
rect -142 -1422 -130 -1388
rect -96 -1422 -84 -1388
rect -142 -1456 -84 -1422
rect -142 -1490 -130 -1456
rect -96 -1490 -84 -1456
rect -142 -1505 -84 -1490
rect 116 -1320 174 -1305
rect 116 -1354 128 -1320
rect 162 -1354 174 -1320
rect 116 -1388 174 -1354
rect 116 -1422 128 -1388
rect 162 -1422 174 -1388
rect 116 -1456 174 -1422
rect 116 -1490 128 -1456
rect 162 -1490 174 -1456
rect 116 -1505 174 -1490
rect 363 -1320 421 -1305
rect 363 -1354 375 -1320
rect 409 -1354 421 -1320
rect 363 -1388 421 -1354
rect 363 -1422 375 -1388
rect 409 -1422 421 -1388
rect 363 -1456 421 -1422
rect 363 -1490 375 -1456
rect 409 -1490 421 -1456
rect 363 -1505 421 -1490
rect 621 -1320 679 -1305
rect 621 -1354 633 -1320
rect 667 -1354 679 -1320
rect 621 -1388 679 -1354
rect 621 -1422 633 -1388
rect 667 -1422 679 -1388
rect 621 -1456 679 -1422
rect 621 -1490 633 -1456
rect 667 -1490 679 -1456
rect 621 -1505 679 -1490
rect 879 -1320 937 -1305
rect 879 -1354 891 -1320
rect 925 -1354 937 -1320
rect 879 -1388 937 -1354
rect 879 -1422 891 -1388
rect 925 -1422 937 -1388
rect 879 -1456 937 -1422
rect 879 -1490 891 -1456
rect 925 -1490 937 -1456
rect 879 -1505 937 -1490
rect 1126 -1320 1184 -1305
rect 1126 -1354 1138 -1320
rect 1172 -1354 1184 -1320
rect 1126 -1388 1184 -1354
rect 1126 -1422 1138 -1388
rect 1172 -1422 1184 -1388
rect 1126 -1456 1184 -1422
rect 1126 -1490 1138 -1456
rect 1172 -1490 1184 -1456
rect 1126 -1505 1184 -1490
rect 1384 -1320 1442 -1305
rect 1384 -1354 1396 -1320
rect 1430 -1354 1442 -1320
rect 1384 -1388 1442 -1354
rect 1384 -1422 1396 -1388
rect 1430 -1422 1442 -1388
rect 1384 -1456 1442 -1422
rect 1384 -1490 1396 -1456
rect 1430 -1490 1442 -1456
rect 1384 -1505 1442 -1490
rect 1642 -1320 1700 -1305
rect 1642 -1354 1654 -1320
rect 1688 -1354 1700 -1320
rect 1642 -1388 1700 -1354
rect 1642 -1422 1654 -1388
rect 1688 -1422 1700 -1388
rect 1642 -1456 1700 -1422
rect 1642 -1490 1654 -1456
rect 1688 -1490 1700 -1456
rect 1642 -1505 1700 -1490
rect 1900 -1320 1958 -1305
rect 1900 -1354 1912 -1320
rect 1946 -1354 1958 -1320
rect 1900 -1388 1958 -1354
rect 1900 -1422 1912 -1388
rect 1946 -1422 1958 -1388
rect 1900 -1456 1958 -1422
rect 1900 -1490 1912 -1456
rect 1946 -1490 1958 -1456
rect 1900 -1505 1958 -1490
rect 2147 -1320 2205 -1305
rect 2147 -1354 2159 -1320
rect 2193 -1354 2205 -1320
rect 2147 -1388 2205 -1354
rect 2147 -1422 2159 -1388
rect 2193 -1422 2205 -1388
rect 2147 -1456 2205 -1422
rect 2147 -1490 2159 -1456
rect 2193 -1490 2205 -1456
rect 2147 -1505 2205 -1490
rect 2405 -1320 2463 -1305
rect 2405 -1354 2417 -1320
rect 2451 -1354 2463 -1320
rect 2405 -1388 2463 -1354
rect 2405 -1422 2417 -1388
rect 2451 -1422 2463 -1388
rect 2405 -1456 2463 -1422
rect 2405 -1490 2417 -1456
rect 2451 -1490 2463 -1456
rect 2405 -1505 2463 -1490
rect 2663 -1320 2721 -1305
rect 2663 -1354 2675 -1320
rect 2709 -1354 2721 -1320
rect 2663 -1388 2721 -1354
rect 2663 -1422 2675 -1388
rect 2709 -1422 2721 -1388
rect 2663 -1456 2721 -1422
rect 2663 -1490 2675 -1456
rect 2709 -1490 2721 -1456
rect 2663 -1505 2721 -1490
rect 2911 -1320 2969 -1305
rect 2911 -1354 2923 -1320
rect 2957 -1354 2969 -1320
rect 2911 -1388 2969 -1354
rect 2911 -1422 2923 -1388
rect 2957 -1422 2969 -1388
rect 2911 -1456 2969 -1422
rect 2911 -1490 2923 -1456
rect 2957 -1490 2969 -1456
rect 2911 -1505 2969 -1490
rect 3169 -1320 3227 -1305
rect 3169 -1354 3181 -1320
rect 3215 -1354 3227 -1320
rect 3169 -1388 3227 -1354
rect 3169 -1422 3181 -1388
rect 3215 -1422 3227 -1388
rect 3169 -1456 3227 -1422
rect 3169 -1490 3181 -1456
rect 3215 -1490 3227 -1456
rect 3169 -1505 3227 -1490
rect 3397 -1320 3455 -1305
rect 3397 -1354 3409 -1320
rect 3443 -1354 3455 -1320
rect 3397 -1388 3455 -1354
rect 3397 -1422 3409 -1388
rect 3443 -1422 3455 -1388
rect 3397 -1456 3455 -1422
rect 3397 -1490 3409 -1456
rect 3443 -1490 3455 -1456
rect 3397 -1505 3455 -1490
rect 3655 -1320 3713 -1305
rect 3655 -1354 3667 -1320
rect 3701 -1354 3713 -1320
rect 3655 -1388 3713 -1354
rect 3655 -1422 3667 -1388
rect 3701 -1422 3713 -1388
rect 3655 -1456 3713 -1422
rect 3655 -1490 3667 -1456
rect 3701 -1490 3713 -1456
rect 3655 -1505 3713 -1490
rect 3903 -1320 3961 -1305
rect 3903 -1354 3915 -1320
rect 3949 -1354 3961 -1320
rect 3903 -1388 3961 -1354
rect 3903 -1422 3915 -1388
rect 3949 -1422 3961 -1388
rect 3903 -1456 3961 -1422
rect 3903 -1490 3915 -1456
rect 3949 -1490 3961 -1456
rect 3903 -1505 3961 -1490
rect 4161 -1320 4219 -1305
rect 4161 -1354 4173 -1320
rect 4207 -1354 4219 -1320
rect 4161 -1388 4219 -1354
rect 4161 -1422 4173 -1388
rect 4207 -1422 4219 -1388
rect 4161 -1456 4219 -1422
rect 4161 -1490 4173 -1456
rect 4207 -1490 4219 -1456
rect 4161 -1505 4219 -1490
rect 4419 -1320 4477 -1305
rect 4419 -1354 4431 -1320
rect 4465 -1354 4477 -1320
rect 4419 -1388 4477 -1354
rect 4419 -1422 4431 -1388
rect 4465 -1422 4477 -1388
rect 4419 -1456 4477 -1422
rect 4419 -1490 4431 -1456
rect 4465 -1490 4477 -1456
rect 4419 -1505 4477 -1490
rect 4666 -1320 4724 -1305
rect 4666 -1354 4678 -1320
rect 4712 -1354 4724 -1320
rect 4666 -1388 4724 -1354
rect 4666 -1422 4678 -1388
rect 4712 -1422 4724 -1388
rect 4666 -1456 4724 -1422
rect 4666 -1490 4678 -1456
rect 4712 -1490 4724 -1456
rect 4666 -1505 4724 -1490
rect 4924 -1320 4982 -1305
rect 4924 -1354 4936 -1320
rect 4970 -1354 4982 -1320
rect 4924 -1388 4982 -1354
rect 4924 -1422 4936 -1388
rect 4970 -1422 4982 -1388
rect 4924 -1456 4982 -1422
rect 4924 -1490 4936 -1456
rect 4970 -1490 4982 -1456
rect 4924 -1505 4982 -1490
rect 5182 -1320 5240 -1305
rect 5182 -1354 5194 -1320
rect 5228 -1354 5240 -1320
rect 5182 -1388 5240 -1354
rect 5182 -1422 5194 -1388
rect 5228 -1422 5240 -1388
rect 5182 -1456 5240 -1422
rect 5182 -1490 5194 -1456
rect 5228 -1490 5240 -1456
rect 5182 -1505 5240 -1490
rect 5440 -1320 5498 -1305
rect 5440 -1354 5452 -1320
rect 5486 -1354 5498 -1320
rect 5440 -1388 5498 -1354
rect 5440 -1422 5452 -1388
rect 5486 -1422 5498 -1388
rect 5440 -1456 5498 -1422
rect 5440 -1490 5452 -1456
rect 5486 -1490 5498 -1456
rect 5440 -1505 5498 -1490
rect 5687 -1320 5745 -1305
rect 5687 -1354 5699 -1320
rect 5733 -1354 5745 -1320
rect 5687 -1388 5745 -1354
rect 5687 -1422 5699 -1388
rect 5733 -1422 5745 -1388
rect 5687 -1456 5745 -1422
rect 5687 -1490 5699 -1456
rect 5733 -1490 5745 -1456
rect 5687 -1505 5745 -1490
rect 5945 -1320 6003 -1305
rect 5945 -1354 5957 -1320
rect 5991 -1354 6003 -1320
rect 5945 -1388 6003 -1354
rect 5945 -1422 5957 -1388
rect 5991 -1422 6003 -1388
rect 5945 -1456 6003 -1422
rect 5945 -1490 5957 -1456
rect 5991 -1490 6003 -1456
rect 5945 -1505 6003 -1490
rect 6203 -1320 6261 -1305
rect 6203 -1354 6215 -1320
rect 6249 -1354 6261 -1320
rect 6203 -1388 6261 -1354
rect 6203 -1422 6215 -1388
rect 6249 -1422 6261 -1388
rect 6203 -1456 6261 -1422
rect 6203 -1490 6215 -1456
rect 6249 -1490 6261 -1456
rect 6203 -1505 6261 -1490
rect 6450 -1320 6508 -1305
rect 6450 -1354 6462 -1320
rect 6496 -1354 6508 -1320
rect 6450 -1388 6508 -1354
rect 6450 -1422 6462 -1388
rect 6496 -1422 6508 -1388
rect 6450 -1456 6508 -1422
rect 6450 -1490 6462 -1456
rect 6496 -1490 6508 -1456
rect 6450 -1505 6508 -1490
rect 6708 -1320 6766 -1305
rect 6708 -1354 6720 -1320
rect 6754 -1354 6766 -1320
rect 6708 -1388 6766 -1354
rect 6708 -1422 6720 -1388
rect 6754 -1422 6766 -1388
rect 6708 -1456 6766 -1422
rect 6708 -1490 6720 -1456
rect 6754 -1490 6766 -1456
rect 6708 -1505 6766 -1490
rect -142 -1993 -84 -1978
rect -142 -2027 -130 -1993
rect -96 -2027 -84 -1993
rect -142 -2061 -84 -2027
rect -142 -2095 -130 -2061
rect -96 -2095 -84 -2061
rect -142 -2129 -84 -2095
rect -142 -2163 -130 -2129
rect -96 -2163 -84 -2129
rect -142 -2178 -84 -2163
rect 116 -1993 174 -1978
rect 116 -2027 128 -1993
rect 162 -2027 174 -1993
rect 116 -2061 174 -2027
rect 116 -2095 128 -2061
rect 162 -2095 174 -2061
rect 116 -2129 174 -2095
rect 116 -2163 128 -2129
rect 162 -2163 174 -2129
rect 116 -2178 174 -2163
rect 363 -1993 421 -1978
rect 363 -2027 375 -1993
rect 409 -2027 421 -1993
rect 363 -2061 421 -2027
rect 363 -2095 375 -2061
rect 409 -2095 421 -2061
rect 363 -2129 421 -2095
rect 363 -2163 375 -2129
rect 409 -2163 421 -2129
rect 363 -2178 421 -2163
rect 621 -1993 679 -1978
rect 621 -2027 633 -1993
rect 667 -2027 679 -1993
rect 621 -2061 679 -2027
rect 621 -2095 633 -2061
rect 667 -2095 679 -2061
rect 621 -2129 679 -2095
rect 621 -2163 633 -2129
rect 667 -2163 679 -2129
rect 621 -2178 679 -2163
rect 879 -1993 937 -1978
rect 879 -2027 891 -1993
rect 925 -2027 937 -1993
rect 879 -2061 937 -2027
rect 879 -2095 891 -2061
rect 925 -2095 937 -2061
rect 879 -2129 937 -2095
rect 879 -2163 891 -2129
rect 925 -2163 937 -2129
rect 879 -2178 937 -2163
rect 1126 -1993 1184 -1978
rect 1126 -2027 1138 -1993
rect 1172 -2027 1184 -1993
rect 1126 -2061 1184 -2027
rect 1126 -2095 1138 -2061
rect 1172 -2095 1184 -2061
rect 1126 -2129 1184 -2095
rect 1126 -2163 1138 -2129
rect 1172 -2163 1184 -2129
rect 1126 -2178 1184 -2163
rect 1384 -1993 1442 -1978
rect 1384 -2027 1396 -1993
rect 1430 -2027 1442 -1993
rect 1384 -2061 1442 -2027
rect 1384 -2095 1396 -2061
rect 1430 -2095 1442 -2061
rect 1384 -2129 1442 -2095
rect 1384 -2163 1396 -2129
rect 1430 -2163 1442 -2129
rect 1384 -2178 1442 -2163
rect 1642 -1993 1700 -1978
rect 1642 -2027 1654 -1993
rect 1688 -2027 1700 -1993
rect 1642 -2061 1700 -2027
rect 1642 -2095 1654 -2061
rect 1688 -2095 1700 -2061
rect 1642 -2129 1700 -2095
rect 1642 -2163 1654 -2129
rect 1688 -2163 1700 -2129
rect 1642 -2178 1700 -2163
rect 1900 -1993 1958 -1978
rect 1900 -2027 1912 -1993
rect 1946 -2027 1958 -1993
rect 1900 -2061 1958 -2027
rect 1900 -2095 1912 -2061
rect 1946 -2095 1958 -2061
rect 1900 -2129 1958 -2095
rect 1900 -2163 1912 -2129
rect 1946 -2163 1958 -2129
rect 1900 -2178 1958 -2163
rect 2147 -1993 2205 -1978
rect 2147 -2027 2159 -1993
rect 2193 -2027 2205 -1993
rect 2147 -2061 2205 -2027
rect 2147 -2095 2159 -2061
rect 2193 -2095 2205 -2061
rect 2147 -2129 2205 -2095
rect 2147 -2163 2159 -2129
rect 2193 -2163 2205 -2129
rect 2147 -2178 2205 -2163
rect 2405 -1993 2463 -1978
rect 2405 -2027 2417 -1993
rect 2451 -2027 2463 -1993
rect 2405 -2061 2463 -2027
rect 2405 -2095 2417 -2061
rect 2451 -2095 2463 -2061
rect 2405 -2129 2463 -2095
rect 2405 -2163 2417 -2129
rect 2451 -2163 2463 -2129
rect 2405 -2178 2463 -2163
rect 2663 -1993 2721 -1978
rect 2663 -2027 2675 -1993
rect 2709 -2027 2721 -1993
rect 2663 -2061 2721 -2027
rect 2663 -2095 2675 -2061
rect 2709 -2095 2721 -2061
rect 2663 -2129 2721 -2095
rect 2663 -2163 2675 -2129
rect 2709 -2163 2721 -2129
rect 2663 -2178 2721 -2163
rect 2911 -1993 2969 -1978
rect 2911 -2027 2923 -1993
rect 2957 -2027 2969 -1993
rect 2911 -2061 2969 -2027
rect 2911 -2095 2923 -2061
rect 2957 -2095 2969 -2061
rect 2911 -2129 2969 -2095
rect 2911 -2163 2923 -2129
rect 2957 -2163 2969 -2129
rect 2911 -2178 2969 -2163
rect 3169 -1993 3227 -1978
rect 3169 -2027 3181 -1993
rect 3215 -2027 3227 -1993
rect 3169 -2061 3227 -2027
rect 3169 -2095 3181 -2061
rect 3215 -2095 3227 -2061
rect 3169 -2129 3227 -2095
rect 3169 -2163 3181 -2129
rect 3215 -2163 3227 -2129
rect 3169 -2178 3227 -2163
rect 3397 -1993 3455 -1978
rect 3397 -2027 3409 -1993
rect 3443 -2027 3455 -1993
rect 3397 -2061 3455 -2027
rect 3397 -2095 3409 -2061
rect 3443 -2095 3455 -2061
rect 3397 -2129 3455 -2095
rect 3397 -2163 3409 -2129
rect 3443 -2163 3455 -2129
rect 3397 -2178 3455 -2163
rect 3655 -1993 3713 -1978
rect 3655 -2027 3667 -1993
rect 3701 -2027 3713 -1993
rect 3655 -2061 3713 -2027
rect 3655 -2095 3667 -2061
rect 3701 -2095 3713 -2061
rect 3655 -2129 3713 -2095
rect 3655 -2163 3667 -2129
rect 3701 -2163 3713 -2129
rect 3655 -2178 3713 -2163
rect 3903 -1993 3961 -1978
rect 3903 -2027 3915 -1993
rect 3949 -2027 3961 -1993
rect 3903 -2061 3961 -2027
rect 3903 -2095 3915 -2061
rect 3949 -2095 3961 -2061
rect 3903 -2129 3961 -2095
rect 3903 -2163 3915 -2129
rect 3949 -2163 3961 -2129
rect 3903 -2178 3961 -2163
rect 4161 -1993 4219 -1978
rect 4161 -2027 4173 -1993
rect 4207 -2027 4219 -1993
rect 4161 -2061 4219 -2027
rect 4161 -2095 4173 -2061
rect 4207 -2095 4219 -2061
rect 4161 -2129 4219 -2095
rect 4161 -2163 4173 -2129
rect 4207 -2163 4219 -2129
rect 4161 -2178 4219 -2163
rect 4419 -1993 4477 -1978
rect 4419 -2027 4431 -1993
rect 4465 -2027 4477 -1993
rect 4419 -2061 4477 -2027
rect 4419 -2095 4431 -2061
rect 4465 -2095 4477 -2061
rect 4419 -2129 4477 -2095
rect 4419 -2163 4431 -2129
rect 4465 -2163 4477 -2129
rect 4419 -2178 4477 -2163
rect 4666 -1993 4724 -1978
rect 4666 -2027 4678 -1993
rect 4712 -2027 4724 -1993
rect 4666 -2061 4724 -2027
rect 4666 -2095 4678 -2061
rect 4712 -2095 4724 -2061
rect 4666 -2129 4724 -2095
rect 4666 -2163 4678 -2129
rect 4712 -2163 4724 -2129
rect 4666 -2178 4724 -2163
rect 4924 -1993 4982 -1978
rect 4924 -2027 4936 -1993
rect 4970 -2027 4982 -1993
rect 4924 -2061 4982 -2027
rect 4924 -2095 4936 -2061
rect 4970 -2095 4982 -2061
rect 4924 -2129 4982 -2095
rect 4924 -2163 4936 -2129
rect 4970 -2163 4982 -2129
rect 4924 -2178 4982 -2163
rect 5182 -1993 5240 -1978
rect 5182 -2027 5194 -1993
rect 5228 -2027 5240 -1993
rect 5182 -2061 5240 -2027
rect 5182 -2095 5194 -2061
rect 5228 -2095 5240 -2061
rect 5182 -2129 5240 -2095
rect 5182 -2163 5194 -2129
rect 5228 -2163 5240 -2129
rect 5182 -2178 5240 -2163
rect 5440 -1993 5498 -1978
rect 5440 -2027 5452 -1993
rect 5486 -2027 5498 -1993
rect 5440 -2061 5498 -2027
rect 5440 -2095 5452 -2061
rect 5486 -2095 5498 -2061
rect 5440 -2129 5498 -2095
rect 5440 -2163 5452 -2129
rect 5486 -2163 5498 -2129
rect 5440 -2178 5498 -2163
rect 5687 -1993 5745 -1978
rect 5687 -2027 5699 -1993
rect 5733 -2027 5745 -1993
rect 5687 -2061 5745 -2027
rect 5687 -2095 5699 -2061
rect 5733 -2095 5745 -2061
rect 5687 -2129 5745 -2095
rect 5687 -2163 5699 -2129
rect 5733 -2163 5745 -2129
rect 5687 -2178 5745 -2163
rect 5945 -1993 6003 -1978
rect 5945 -2027 5957 -1993
rect 5991 -2027 6003 -1993
rect 5945 -2061 6003 -2027
rect 5945 -2095 5957 -2061
rect 5991 -2095 6003 -2061
rect 5945 -2129 6003 -2095
rect 5945 -2163 5957 -2129
rect 5991 -2163 6003 -2129
rect 5945 -2178 6003 -2163
rect 6203 -1993 6261 -1978
rect 6203 -2027 6215 -1993
rect 6249 -2027 6261 -1993
rect 6203 -2061 6261 -2027
rect 6203 -2095 6215 -2061
rect 6249 -2095 6261 -2061
rect 6203 -2129 6261 -2095
rect 6203 -2163 6215 -2129
rect 6249 -2163 6261 -2129
rect 6203 -2178 6261 -2163
rect 6450 -1993 6508 -1978
rect 6450 -2027 6462 -1993
rect 6496 -2027 6508 -1993
rect 6450 -2061 6508 -2027
rect 6450 -2095 6462 -2061
rect 6496 -2095 6508 -2061
rect 6450 -2129 6508 -2095
rect 6450 -2163 6462 -2129
rect 6496 -2163 6508 -2129
rect 6450 -2178 6508 -2163
rect 6708 -1993 6766 -1978
rect 6708 -2027 6720 -1993
rect 6754 -2027 6766 -1993
rect 6708 -2061 6766 -2027
rect 6708 -2095 6720 -2061
rect 6754 -2095 6766 -2061
rect 6708 -2129 6766 -2095
rect 6708 -2163 6720 -2129
rect 6754 -2163 6766 -2129
rect 6708 -2178 6766 -2163
rect -142 -2719 -84 -2704
rect -142 -2753 -130 -2719
rect -96 -2753 -84 -2719
rect -142 -2787 -84 -2753
rect -142 -2821 -130 -2787
rect -96 -2821 -84 -2787
rect -142 -2855 -84 -2821
rect -142 -2889 -130 -2855
rect -96 -2889 -84 -2855
rect -142 -2904 -84 -2889
rect 116 -2719 174 -2704
rect 116 -2753 128 -2719
rect 162 -2753 174 -2719
rect 116 -2787 174 -2753
rect 116 -2821 128 -2787
rect 162 -2821 174 -2787
rect 116 -2855 174 -2821
rect 116 -2889 128 -2855
rect 162 -2889 174 -2855
rect 116 -2904 174 -2889
rect 363 -2719 421 -2704
rect 363 -2753 375 -2719
rect 409 -2753 421 -2719
rect 363 -2787 421 -2753
rect 363 -2821 375 -2787
rect 409 -2821 421 -2787
rect 363 -2855 421 -2821
rect 363 -2889 375 -2855
rect 409 -2889 421 -2855
rect 363 -2904 421 -2889
rect 621 -2719 679 -2704
rect 621 -2753 633 -2719
rect 667 -2753 679 -2719
rect 621 -2787 679 -2753
rect 621 -2821 633 -2787
rect 667 -2821 679 -2787
rect 621 -2855 679 -2821
rect 621 -2889 633 -2855
rect 667 -2889 679 -2855
rect 621 -2904 679 -2889
rect 879 -2719 937 -2704
rect 879 -2753 891 -2719
rect 925 -2753 937 -2719
rect 879 -2787 937 -2753
rect 879 -2821 891 -2787
rect 925 -2821 937 -2787
rect 879 -2855 937 -2821
rect 879 -2889 891 -2855
rect 925 -2889 937 -2855
rect 879 -2904 937 -2889
rect 1126 -2719 1184 -2704
rect 1126 -2753 1138 -2719
rect 1172 -2753 1184 -2719
rect 1126 -2787 1184 -2753
rect 1126 -2821 1138 -2787
rect 1172 -2821 1184 -2787
rect 1126 -2855 1184 -2821
rect 1126 -2889 1138 -2855
rect 1172 -2889 1184 -2855
rect 1126 -2904 1184 -2889
rect 1384 -2719 1442 -2704
rect 1384 -2753 1396 -2719
rect 1430 -2753 1442 -2719
rect 1384 -2787 1442 -2753
rect 1384 -2821 1396 -2787
rect 1430 -2821 1442 -2787
rect 1384 -2855 1442 -2821
rect 1384 -2889 1396 -2855
rect 1430 -2889 1442 -2855
rect 1384 -2904 1442 -2889
rect 1642 -2719 1700 -2704
rect 1642 -2753 1654 -2719
rect 1688 -2753 1700 -2719
rect 1642 -2787 1700 -2753
rect 1642 -2821 1654 -2787
rect 1688 -2821 1700 -2787
rect 1642 -2855 1700 -2821
rect 1642 -2889 1654 -2855
rect 1688 -2889 1700 -2855
rect 1642 -2904 1700 -2889
rect 1900 -2719 1958 -2704
rect 1900 -2753 1912 -2719
rect 1946 -2753 1958 -2719
rect 1900 -2787 1958 -2753
rect 1900 -2821 1912 -2787
rect 1946 -2821 1958 -2787
rect 1900 -2855 1958 -2821
rect 1900 -2889 1912 -2855
rect 1946 -2889 1958 -2855
rect 1900 -2904 1958 -2889
rect 2147 -2719 2205 -2704
rect 2147 -2753 2159 -2719
rect 2193 -2753 2205 -2719
rect 2147 -2787 2205 -2753
rect 2147 -2821 2159 -2787
rect 2193 -2821 2205 -2787
rect 2147 -2855 2205 -2821
rect 2147 -2889 2159 -2855
rect 2193 -2889 2205 -2855
rect 2147 -2904 2205 -2889
rect 2405 -2719 2463 -2704
rect 2405 -2753 2417 -2719
rect 2451 -2753 2463 -2719
rect 2405 -2787 2463 -2753
rect 2405 -2821 2417 -2787
rect 2451 -2821 2463 -2787
rect 2405 -2855 2463 -2821
rect 2405 -2889 2417 -2855
rect 2451 -2889 2463 -2855
rect 2405 -2904 2463 -2889
rect 2663 -2719 2721 -2704
rect 2663 -2753 2675 -2719
rect 2709 -2753 2721 -2719
rect 2663 -2787 2721 -2753
rect 2663 -2821 2675 -2787
rect 2709 -2821 2721 -2787
rect 2663 -2855 2721 -2821
rect 2663 -2889 2675 -2855
rect 2709 -2889 2721 -2855
rect 2663 -2904 2721 -2889
rect 2911 -2719 2969 -2704
rect 2911 -2753 2923 -2719
rect 2957 -2753 2969 -2719
rect 2911 -2787 2969 -2753
rect 2911 -2821 2923 -2787
rect 2957 -2821 2969 -2787
rect 2911 -2855 2969 -2821
rect 2911 -2889 2923 -2855
rect 2957 -2889 2969 -2855
rect 2911 -2904 2969 -2889
rect 3169 -2719 3227 -2704
rect 3169 -2753 3181 -2719
rect 3215 -2753 3227 -2719
rect 3169 -2787 3227 -2753
rect 3169 -2821 3181 -2787
rect 3215 -2821 3227 -2787
rect 3169 -2855 3227 -2821
rect 3169 -2889 3181 -2855
rect 3215 -2889 3227 -2855
rect 3169 -2904 3227 -2889
rect 3397 -2719 3455 -2704
rect 3397 -2753 3409 -2719
rect 3443 -2753 3455 -2719
rect 3397 -2787 3455 -2753
rect 3397 -2821 3409 -2787
rect 3443 -2821 3455 -2787
rect 3397 -2855 3455 -2821
rect 3397 -2889 3409 -2855
rect 3443 -2889 3455 -2855
rect 3397 -2904 3455 -2889
rect 3655 -2719 3713 -2704
rect 3655 -2753 3667 -2719
rect 3701 -2753 3713 -2719
rect 3655 -2787 3713 -2753
rect 3655 -2821 3667 -2787
rect 3701 -2821 3713 -2787
rect 3655 -2855 3713 -2821
rect 3655 -2889 3667 -2855
rect 3701 -2889 3713 -2855
rect 3655 -2904 3713 -2889
rect 3903 -2719 3961 -2704
rect 3903 -2753 3915 -2719
rect 3949 -2753 3961 -2719
rect 3903 -2787 3961 -2753
rect 3903 -2821 3915 -2787
rect 3949 -2821 3961 -2787
rect 3903 -2855 3961 -2821
rect 3903 -2889 3915 -2855
rect 3949 -2889 3961 -2855
rect 3903 -2904 3961 -2889
rect 4161 -2719 4219 -2704
rect 4161 -2753 4173 -2719
rect 4207 -2753 4219 -2719
rect 4161 -2787 4219 -2753
rect 4161 -2821 4173 -2787
rect 4207 -2821 4219 -2787
rect 4161 -2855 4219 -2821
rect 4161 -2889 4173 -2855
rect 4207 -2889 4219 -2855
rect 4161 -2904 4219 -2889
rect 4419 -2719 4477 -2704
rect 4419 -2753 4431 -2719
rect 4465 -2753 4477 -2719
rect 4419 -2787 4477 -2753
rect 4419 -2821 4431 -2787
rect 4465 -2821 4477 -2787
rect 4419 -2855 4477 -2821
rect 4419 -2889 4431 -2855
rect 4465 -2889 4477 -2855
rect 4419 -2904 4477 -2889
rect 4666 -2719 4724 -2704
rect 4666 -2753 4678 -2719
rect 4712 -2753 4724 -2719
rect 4666 -2787 4724 -2753
rect 4666 -2821 4678 -2787
rect 4712 -2821 4724 -2787
rect 4666 -2855 4724 -2821
rect 4666 -2889 4678 -2855
rect 4712 -2889 4724 -2855
rect 4666 -2904 4724 -2889
rect 4924 -2719 4982 -2704
rect 4924 -2753 4936 -2719
rect 4970 -2753 4982 -2719
rect 4924 -2787 4982 -2753
rect 4924 -2821 4936 -2787
rect 4970 -2821 4982 -2787
rect 4924 -2855 4982 -2821
rect 4924 -2889 4936 -2855
rect 4970 -2889 4982 -2855
rect 4924 -2904 4982 -2889
rect 5182 -2719 5240 -2704
rect 5182 -2753 5194 -2719
rect 5228 -2753 5240 -2719
rect 5182 -2787 5240 -2753
rect 5182 -2821 5194 -2787
rect 5228 -2821 5240 -2787
rect 5182 -2855 5240 -2821
rect 5182 -2889 5194 -2855
rect 5228 -2889 5240 -2855
rect 5182 -2904 5240 -2889
rect 5440 -2719 5498 -2704
rect 5440 -2753 5452 -2719
rect 5486 -2753 5498 -2719
rect 5440 -2787 5498 -2753
rect 5440 -2821 5452 -2787
rect 5486 -2821 5498 -2787
rect 5440 -2855 5498 -2821
rect 5440 -2889 5452 -2855
rect 5486 -2889 5498 -2855
rect 5440 -2904 5498 -2889
rect 5687 -2719 5745 -2704
rect 5687 -2753 5699 -2719
rect 5733 -2753 5745 -2719
rect 5687 -2787 5745 -2753
rect 5687 -2821 5699 -2787
rect 5733 -2821 5745 -2787
rect 5687 -2855 5745 -2821
rect 5687 -2889 5699 -2855
rect 5733 -2889 5745 -2855
rect 5687 -2904 5745 -2889
rect 5945 -2719 6003 -2704
rect 5945 -2753 5957 -2719
rect 5991 -2753 6003 -2719
rect 5945 -2787 6003 -2753
rect 5945 -2821 5957 -2787
rect 5991 -2821 6003 -2787
rect 5945 -2855 6003 -2821
rect 5945 -2889 5957 -2855
rect 5991 -2889 6003 -2855
rect 5945 -2904 6003 -2889
rect 6203 -2719 6261 -2704
rect 6203 -2753 6215 -2719
rect 6249 -2753 6261 -2719
rect 6203 -2787 6261 -2753
rect 6203 -2821 6215 -2787
rect 6249 -2821 6261 -2787
rect 6203 -2855 6261 -2821
rect 6203 -2889 6215 -2855
rect 6249 -2889 6261 -2855
rect 6203 -2904 6261 -2889
rect 6450 -2719 6508 -2704
rect 6450 -2753 6462 -2719
rect 6496 -2753 6508 -2719
rect 6450 -2787 6508 -2753
rect 6450 -2821 6462 -2787
rect 6496 -2821 6508 -2787
rect 6450 -2855 6508 -2821
rect 6450 -2889 6462 -2855
rect 6496 -2889 6508 -2855
rect 6450 -2904 6508 -2889
rect 6708 -2719 6766 -2704
rect 6708 -2753 6720 -2719
rect 6754 -2753 6766 -2719
rect 6708 -2787 6766 -2753
rect 6708 -2821 6720 -2787
rect 6754 -2821 6766 -2787
rect 6708 -2855 6766 -2821
rect 6708 -2889 6720 -2855
rect 6754 -2889 6766 -2855
rect 6708 -2904 6766 -2889
<< ndiffc >>
rect -130 769 -96 803
rect -130 701 -96 735
rect -130 633 -96 667
rect 128 769 162 803
rect 128 701 162 735
rect 128 633 162 667
rect 375 769 409 803
rect 375 701 409 735
rect 375 633 409 667
rect 633 769 667 803
rect 633 701 667 735
rect 633 633 667 667
rect 891 769 925 803
rect 891 701 925 735
rect 891 633 925 667
rect 1138 769 1172 803
rect 1138 701 1172 735
rect 1138 633 1172 667
rect 1396 769 1430 803
rect 1396 701 1430 735
rect 1396 633 1430 667
rect 1654 769 1688 803
rect 1654 701 1688 735
rect 1654 633 1688 667
rect 1912 769 1946 803
rect 1912 701 1946 735
rect 1912 633 1946 667
rect 2159 769 2193 803
rect 2159 701 2193 735
rect 2159 633 2193 667
rect 2417 769 2451 803
rect 2417 701 2451 735
rect 2417 633 2451 667
rect 2675 769 2709 803
rect 2675 701 2709 735
rect 2675 633 2709 667
rect 2923 769 2957 803
rect 2923 701 2957 735
rect 2923 633 2957 667
rect 3181 769 3215 803
rect 3181 701 3215 735
rect 3181 633 3215 667
rect 3409 769 3443 803
rect 3409 701 3443 735
rect 3409 633 3443 667
rect 3667 769 3701 803
rect 3667 701 3701 735
rect 3667 633 3701 667
rect 3915 769 3949 803
rect 3915 701 3949 735
rect 3915 633 3949 667
rect 4173 769 4207 803
rect 4173 701 4207 735
rect 4173 633 4207 667
rect 4431 769 4465 803
rect 4431 701 4465 735
rect 4431 633 4465 667
rect 4678 769 4712 803
rect 4678 701 4712 735
rect 4678 633 4712 667
rect 4936 769 4970 803
rect 4936 701 4970 735
rect 4936 633 4970 667
rect 5194 769 5228 803
rect 5194 701 5228 735
rect 5194 633 5228 667
rect 5452 769 5486 803
rect 5452 701 5486 735
rect 5452 633 5486 667
rect 5699 769 5733 803
rect 5699 701 5733 735
rect 5699 633 5733 667
rect 5957 769 5991 803
rect 5957 701 5991 735
rect 5957 633 5991 667
rect 6215 769 6249 803
rect 6215 701 6249 735
rect 6215 633 6249 667
rect 6462 769 6496 803
rect 6462 701 6496 735
rect 6462 633 6496 667
rect 6720 769 6754 803
rect 6720 701 6754 735
rect 6720 633 6754 667
rect -130 43 -96 77
rect -130 -25 -96 9
rect -130 -93 -96 -59
rect 128 43 162 77
rect 128 -25 162 9
rect 128 -93 162 -59
rect 375 43 409 77
rect 375 -25 409 9
rect 375 -93 409 -59
rect 633 43 667 77
rect 633 -25 667 9
rect 633 -93 667 -59
rect 891 43 925 77
rect 891 -25 925 9
rect 891 -93 925 -59
rect 1138 43 1172 77
rect 1138 -25 1172 9
rect 1138 -93 1172 -59
rect 1396 43 1430 77
rect 1396 -25 1430 9
rect 1396 -93 1430 -59
rect 1654 43 1688 77
rect 1654 -25 1688 9
rect 1654 -93 1688 -59
rect 1912 43 1946 77
rect 1912 -25 1946 9
rect 1912 -93 1946 -59
rect 2159 43 2193 77
rect 2159 -25 2193 9
rect 2159 -93 2193 -59
rect 2417 43 2451 77
rect 2417 -25 2451 9
rect 2417 -93 2451 -59
rect 2675 43 2709 77
rect 2675 -25 2709 9
rect 2675 -93 2709 -59
rect 2923 43 2957 77
rect 2923 -25 2957 9
rect 2923 -93 2957 -59
rect 3181 43 3215 77
rect 3181 -25 3215 9
rect 3181 -93 3215 -59
rect 3409 43 3443 77
rect 3409 -25 3443 9
rect 3409 -93 3443 -59
rect 3667 43 3701 77
rect 3667 -25 3701 9
rect 3667 -93 3701 -59
rect 3915 43 3949 77
rect 3915 -25 3949 9
rect 3915 -93 3949 -59
rect 4173 43 4207 77
rect 4173 -25 4207 9
rect 4173 -93 4207 -59
rect 4431 43 4465 77
rect 4431 -25 4465 9
rect 4431 -93 4465 -59
rect 4678 43 4712 77
rect 4678 -25 4712 9
rect 4678 -93 4712 -59
rect 4936 43 4970 77
rect 4936 -25 4970 9
rect 4936 -93 4970 -59
rect 5194 43 5228 77
rect 5194 -25 5228 9
rect 5194 -93 5228 -59
rect 5452 43 5486 77
rect 5452 -25 5486 9
rect 5452 -93 5486 -59
rect 5699 43 5733 77
rect 5699 -25 5733 9
rect 5699 -93 5733 -59
rect 5957 43 5991 77
rect 5957 -25 5991 9
rect 5957 -93 5991 -59
rect 6215 43 6249 77
rect 6215 -25 6249 9
rect 6215 -93 6249 -59
rect 6462 43 6496 77
rect 6462 -25 6496 9
rect 6462 -93 6496 -59
rect 6720 43 6754 77
rect 6720 -25 6754 9
rect 6720 -93 6754 -59
rect -130 -630 -96 -596
rect -130 -698 -96 -664
rect -130 -766 -96 -732
rect 128 -630 162 -596
rect 128 -698 162 -664
rect 128 -766 162 -732
rect 375 -630 409 -596
rect 375 -698 409 -664
rect 375 -766 409 -732
rect 633 -630 667 -596
rect 633 -698 667 -664
rect 633 -766 667 -732
rect 891 -630 925 -596
rect 891 -698 925 -664
rect 891 -766 925 -732
rect 1138 -630 1172 -596
rect 1138 -698 1172 -664
rect 1138 -766 1172 -732
rect 1396 -630 1430 -596
rect 1396 -698 1430 -664
rect 1396 -766 1430 -732
rect 1654 -630 1688 -596
rect 1654 -698 1688 -664
rect 1654 -766 1688 -732
rect 1912 -630 1946 -596
rect 1912 -698 1946 -664
rect 1912 -766 1946 -732
rect 2159 -630 2193 -596
rect 2159 -698 2193 -664
rect 2159 -766 2193 -732
rect 2417 -630 2451 -596
rect 2417 -698 2451 -664
rect 2417 -766 2451 -732
rect 2675 -630 2709 -596
rect 2675 -698 2709 -664
rect 2675 -766 2709 -732
rect 2923 -630 2957 -596
rect 2923 -698 2957 -664
rect 2923 -766 2957 -732
rect 3181 -630 3215 -596
rect 3181 -698 3215 -664
rect 3181 -766 3215 -732
rect 3409 -630 3443 -596
rect 3409 -698 3443 -664
rect 3409 -766 3443 -732
rect 3667 -630 3701 -596
rect 3667 -698 3701 -664
rect 3667 -766 3701 -732
rect 3915 -630 3949 -596
rect 3915 -698 3949 -664
rect 3915 -766 3949 -732
rect 4173 -630 4207 -596
rect 4173 -698 4207 -664
rect 4173 -766 4207 -732
rect 4431 -630 4465 -596
rect 4431 -698 4465 -664
rect 4431 -766 4465 -732
rect 4678 -630 4712 -596
rect 4678 -698 4712 -664
rect 4678 -766 4712 -732
rect 4936 -630 4970 -596
rect 4936 -698 4970 -664
rect 4936 -766 4970 -732
rect 5194 -630 5228 -596
rect 5194 -698 5228 -664
rect 5194 -766 5228 -732
rect 5452 -630 5486 -596
rect 5452 -698 5486 -664
rect 5452 -766 5486 -732
rect 5699 -630 5733 -596
rect 5699 -698 5733 -664
rect 5699 -766 5733 -732
rect 5957 -630 5991 -596
rect 5957 -698 5991 -664
rect 5957 -766 5991 -732
rect 6215 -630 6249 -596
rect 6215 -698 6249 -664
rect 6215 -766 6249 -732
rect 6462 -630 6496 -596
rect 6462 -698 6496 -664
rect 6462 -766 6496 -732
rect 6720 -630 6754 -596
rect 6720 -698 6754 -664
rect 6720 -766 6754 -732
rect -130 -1354 -96 -1320
rect -130 -1422 -96 -1388
rect -130 -1490 -96 -1456
rect 128 -1354 162 -1320
rect 128 -1422 162 -1388
rect 128 -1490 162 -1456
rect 375 -1354 409 -1320
rect 375 -1422 409 -1388
rect 375 -1490 409 -1456
rect 633 -1354 667 -1320
rect 633 -1422 667 -1388
rect 633 -1490 667 -1456
rect 891 -1354 925 -1320
rect 891 -1422 925 -1388
rect 891 -1490 925 -1456
rect 1138 -1354 1172 -1320
rect 1138 -1422 1172 -1388
rect 1138 -1490 1172 -1456
rect 1396 -1354 1430 -1320
rect 1396 -1422 1430 -1388
rect 1396 -1490 1430 -1456
rect 1654 -1354 1688 -1320
rect 1654 -1422 1688 -1388
rect 1654 -1490 1688 -1456
rect 1912 -1354 1946 -1320
rect 1912 -1422 1946 -1388
rect 1912 -1490 1946 -1456
rect 2159 -1354 2193 -1320
rect 2159 -1422 2193 -1388
rect 2159 -1490 2193 -1456
rect 2417 -1354 2451 -1320
rect 2417 -1422 2451 -1388
rect 2417 -1490 2451 -1456
rect 2675 -1354 2709 -1320
rect 2675 -1422 2709 -1388
rect 2675 -1490 2709 -1456
rect 2923 -1354 2957 -1320
rect 2923 -1422 2957 -1388
rect 2923 -1490 2957 -1456
rect 3181 -1354 3215 -1320
rect 3181 -1422 3215 -1388
rect 3181 -1490 3215 -1456
rect 3409 -1354 3443 -1320
rect 3409 -1422 3443 -1388
rect 3409 -1490 3443 -1456
rect 3667 -1354 3701 -1320
rect 3667 -1422 3701 -1388
rect 3667 -1490 3701 -1456
rect 3915 -1354 3949 -1320
rect 3915 -1422 3949 -1388
rect 3915 -1490 3949 -1456
rect 4173 -1354 4207 -1320
rect 4173 -1422 4207 -1388
rect 4173 -1490 4207 -1456
rect 4431 -1354 4465 -1320
rect 4431 -1422 4465 -1388
rect 4431 -1490 4465 -1456
rect 4678 -1354 4712 -1320
rect 4678 -1422 4712 -1388
rect 4678 -1490 4712 -1456
rect 4936 -1354 4970 -1320
rect 4936 -1422 4970 -1388
rect 4936 -1490 4970 -1456
rect 5194 -1354 5228 -1320
rect 5194 -1422 5228 -1388
rect 5194 -1490 5228 -1456
rect 5452 -1354 5486 -1320
rect 5452 -1422 5486 -1388
rect 5452 -1490 5486 -1456
rect 5699 -1354 5733 -1320
rect 5699 -1422 5733 -1388
rect 5699 -1490 5733 -1456
rect 5957 -1354 5991 -1320
rect 5957 -1422 5991 -1388
rect 5957 -1490 5991 -1456
rect 6215 -1354 6249 -1320
rect 6215 -1422 6249 -1388
rect 6215 -1490 6249 -1456
rect 6462 -1354 6496 -1320
rect 6462 -1422 6496 -1388
rect 6462 -1490 6496 -1456
rect 6720 -1354 6754 -1320
rect 6720 -1422 6754 -1388
rect 6720 -1490 6754 -1456
rect -130 -2027 -96 -1993
rect -130 -2095 -96 -2061
rect -130 -2163 -96 -2129
rect 128 -2027 162 -1993
rect 128 -2095 162 -2061
rect 128 -2163 162 -2129
rect 375 -2027 409 -1993
rect 375 -2095 409 -2061
rect 375 -2163 409 -2129
rect 633 -2027 667 -1993
rect 633 -2095 667 -2061
rect 633 -2163 667 -2129
rect 891 -2027 925 -1993
rect 891 -2095 925 -2061
rect 891 -2163 925 -2129
rect 1138 -2027 1172 -1993
rect 1138 -2095 1172 -2061
rect 1138 -2163 1172 -2129
rect 1396 -2027 1430 -1993
rect 1396 -2095 1430 -2061
rect 1396 -2163 1430 -2129
rect 1654 -2027 1688 -1993
rect 1654 -2095 1688 -2061
rect 1654 -2163 1688 -2129
rect 1912 -2027 1946 -1993
rect 1912 -2095 1946 -2061
rect 1912 -2163 1946 -2129
rect 2159 -2027 2193 -1993
rect 2159 -2095 2193 -2061
rect 2159 -2163 2193 -2129
rect 2417 -2027 2451 -1993
rect 2417 -2095 2451 -2061
rect 2417 -2163 2451 -2129
rect 2675 -2027 2709 -1993
rect 2675 -2095 2709 -2061
rect 2675 -2163 2709 -2129
rect 2923 -2027 2957 -1993
rect 2923 -2095 2957 -2061
rect 2923 -2163 2957 -2129
rect 3181 -2027 3215 -1993
rect 3181 -2095 3215 -2061
rect 3181 -2163 3215 -2129
rect 3409 -2027 3443 -1993
rect 3409 -2095 3443 -2061
rect 3409 -2163 3443 -2129
rect 3667 -2027 3701 -1993
rect 3667 -2095 3701 -2061
rect 3667 -2163 3701 -2129
rect 3915 -2027 3949 -1993
rect 3915 -2095 3949 -2061
rect 3915 -2163 3949 -2129
rect 4173 -2027 4207 -1993
rect 4173 -2095 4207 -2061
rect 4173 -2163 4207 -2129
rect 4431 -2027 4465 -1993
rect 4431 -2095 4465 -2061
rect 4431 -2163 4465 -2129
rect 4678 -2027 4712 -1993
rect 4678 -2095 4712 -2061
rect 4678 -2163 4712 -2129
rect 4936 -2027 4970 -1993
rect 4936 -2095 4970 -2061
rect 4936 -2163 4970 -2129
rect 5194 -2027 5228 -1993
rect 5194 -2095 5228 -2061
rect 5194 -2163 5228 -2129
rect 5452 -2027 5486 -1993
rect 5452 -2095 5486 -2061
rect 5452 -2163 5486 -2129
rect 5699 -2027 5733 -1993
rect 5699 -2095 5733 -2061
rect 5699 -2163 5733 -2129
rect 5957 -2027 5991 -1993
rect 5957 -2095 5991 -2061
rect 5957 -2163 5991 -2129
rect 6215 -2027 6249 -1993
rect 6215 -2095 6249 -2061
rect 6215 -2163 6249 -2129
rect 6462 -2027 6496 -1993
rect 6462 -2095 6496 -2061
rect 6462 -2163 6496 -2129
rect 6720 -2027 6754 -1993
rect 6720 -2095 6754 -2061
rect 6720 -2163 6754 -2129
rect -130 -2753 -96 -2719
rect -130 -2821 -96 -2787
rect -130 -2889 -96 -2855
rect 128 -2753 162 -2719
rect 128 -2821 162 -2787
rect 128 -2889 162 -2855
rect 375 -2753 409 -2719
rect 375 -2821 409 -2787
rect 375 -2889 409 -2855
rect 633 -2753 667 -2719
rect 633 -2821 667 -2787
rect 633 -2889 667 -2855
rect 891 -2753 925 -2719
rect 891 -2821 925 -2787
rect 891 -2889 925 -2855
rect 1138 -2753 1172 -2719
rect 1138 -2821 1172 -2787
rect 1138 -2889 1172 -2855
rect 1396 -2753 1430 -2719
rect 1396 -2821 1430 -2787
rect 1396 -2889 1430 -2855
rect 1654 -2753 1688 -2719
rect 1654 -2821 1688 -2787
rect 1654 -2889 1688 -2855
rect 1912 -2753 1946 -2719
rect 1912 -2821 1946 -2787
rect 1912 -2889 1946 -2855
rect 2159 -2753 2193 -2719
rect 2159 -2821 2193 -2787
rect 2159 -2889 2193 -2855
rect 2417 -2753 2451 -2719
rect 2417 -2821 2451 -2787
rect 2417 -2889 2451 -2855
rect 2675 -2753 2709 -2719
rect 2675 -2821 2709 -2787
rect 2675 -2889 2709 -2855
rect 2923 -2753 2957 -2719
rect 2923 -2821 2957 -2787
rect 2923 -2889 2957 -2855
rect 3181 -2753 3215 -2719
rect 3181 -2821 3215 -2787
rect 3181 -2889 3215 -2855
rect 3409 -2753 3443 -2719
rect 3409 -2821 3443 -2787
rect 3409 -2889 3443 -2855
rect 3667 -2753 3701 -2719
rect 3667 -2821 3701 -2787
rect 3667 -2889 3701 -2855
rect 3915 -2753 3949 -2719
rect 3915 -2821 3949 -2787
rect 3915 -2889 3949 -2855
rect 4173 -2753 4207 -2719
rect 4173 -2821 4207 -2787
rect 4173 -2889 4207 -2855
rect 4431 -2753 4465 -2719
rect 4431 -2821 4465 -2787
rect 4431 -2889 4465 -2855
rect 4678 -2753 4712 -2719
rect 4678 -2821 4712 -2787
rect 4678 -2889 4712 -2855
rect 4936 -2753 4970 -2719
rect 4936 -2821 4970 -2787
rect 4936 -2889 4970 -2855
rect 5194 -2753 5228 -2719
rect 5194 -2821 5228 -2787
rect 5194 -2889 5228 -2855
rect 5452 -2753 5486 -2719
rect 5452 -2821 5486 -2787
rect 5452 -2889 5486 -2855
rect 5699 -2753 5733 -2719
rect 5699 -2821 5733 -2787
rect 5699 -2889 5733 -2855
rect 5957 -2753 5991 -2719
rect 5957 -2821 5991 -2787
rect 5957 -2889 5991 -2855
rect 6215 -2753 6249 -2719
rect 6215 -2821 6249 -2787
rect 6215 -2889 6249 -2855
rect 6462 -2753 6496 -2719
rect 6462 -2821 6496 -2787
rect 6462 -2889 6496 -2855
rect 6720 -2753 6754 -2719
rect 6720 -2821 6754 -2787
rect 6720 -2889 6754 -2855
<< psubdiff >>
rect -244 955 -59 989
rect -25 955 9 989
rect 43 955 77 989
rect 111 955 145 989
rect 179 955 213 989
rect 247 955 281 989
rect 315 955 349 989
rect 383 955 417 989
rect 451 955 485 989
rect 519 955 553 989
rect 587 955 621 989
rect 655 955 689 989
rect 723 955 757 989
rect 791 955 825 989
rect 859 955 893 989
rect 927 955 961 989
rect 995 955 1029 989
rect 1063 955 1097 989
rect 1131 955 1165 989
rect 1199 955 1233 989
rect 1267 955 1301 989
rect 1335 955 1369 989
rect 1403 955 1437 989
rect 1471 955 1505 989
rect 1539 955 1573 989
rect 1607 955 1641 989
rect 1675 955 1709 989
rect 1743 955 1777 989
rect 1811 955 1845 989
rect 1879 955 1913 989
rect 1947 955 1981 989
rect 2015 955 2049 989
rect 2083 955 2117 989
rect 2151 955 2185 989
rect 2219 955 2253 989
rect 2287 955 2321 989
rect 2355 955 2389 989
rect 2423 955 2457 989
rect 2491 955 2525 989
rect 2559 955 2593 989
rect 2627 955 2661 989
rect 2695 955 2729 989
rect 2763 955 2797 989
rect 2831 955 2865 989
rect 2899 955 2933 989
rect 2967 955 3001 989
rect 3035 955 3069 989
rect 3103 955 3137 989
rect 3171 955 3453 989
rect 3487 955 3521 989
rect 3555 955 3589 989
rect 3623 955 3657 989
rect 3691 955 3725 989
rect 3759 955 3793 989
rect 3827 955 3861 989
rect 3895 955 3929 989
rect 3963 955 3997 989
rect 4031 955 4065 989
rect 4099 955 4133 989
rect 4167 955 4201 989
rect 4235 955 4269 989
rect 4303 955 4337 989
rect 4371 955 4405 989
rect 4439 955 4473 989
rect 4507 955 4541 989
rect 4575 955 4609 989
rect 4643 955 4677 989
rect 4711 955 4745 989
rect 4779 955 4813 989
rect 4847 955 4881 989
rect 4915 955 4949 989
rect 4983 955 5017 989
rect 5051 955 5085 989
rect 5119 955 5153 989
rect 5187 955 5221 989
rect 5255 955 5289 989
rect 5323 955 5357 989
rect 5391 955 5425 989
rect 5459 955 5493 989
rect 5527 955 5561 989
rect 5595 955 5629 989
rect 5663 955 5697 989
rect 5731 955 5765 989
rect 5799 955 5833 989
rect 5867 955 5901 989
rect 5935 955 5969 989
rect 6003 955 6037 989
rect 6071 955 6105 989
rect 6139 955 6173 989
rect 6207 955 6241 989
rect 6275 955 6309 989
rect 6343 955 6377 989
rect 6411 955 6445 989
rect 6479 955 6513 989
rect 6547 955 6581 989
rect 6615 955 6649 989
rect 6683 955 6868 989
rect -244 848 -210 955
rect 3295 848 3329 955
rect -244 780 -210 814
rect -244 712 -210 746
rect -244 644 -210 678
rect 6834 848 6868 955
rect 3295 780 3329 814
rect 3295 712 3329 746
rect 3295 644 3329 678
rect -244 576 -210 610
rect 6834 780 6868 814
rect 6834 712 6868 746
rect 6834 644 6868 678
rect -244 508 -210 542
rect -244 440 -210 474
rect -244 372 -210 406
rect 3295 576 3329 610
rect 3295 508 3329 542
rect 3295 440 3329 474
rect 3295 372 3329 406
rect 6834 576 6868 610
rect 6834 508 6868 542
rect 6834 440 6868 474
rect 6834 372 6868 406
rect -210 338 -59 372
rect -25 338 9 372
rect 43 338 77 372
rect 111 338 145 372
rect 179 338 213 372
rect 247 338 281 372
rect 315 338 349 372
rect 383 338 417 372
rect 451 338 485 372
rect 519 338 553 372
rect 587 338 621 372
rect 655 338 689 372
rect 723 338 757 372
rect 791 338 825 372
rect 859 338 893 372
rect 927 338 961 372
rect 995 338 1029 372
rect 1063 338 1097 372
rect 1131 338 1165 372
rect 1199 338 1233 372
rect 1267 338 1301 372
rect 1335 338 1369 372
rect 1403 338 1437 372
rect 1471 338 1505 372
rect 1539 338 1573 372
rect 1607 338 1641 372
rect 1675 338 1709 372
rect 1743 338 1777 372
rect 1811 338 1845 372
rect 1879 338 1913 372
rect 1947 338 1981 372
rect 2015 338 2049 372
rect 2083 338 2117 372
rect 2151 338 2185 372
rect 2219 338 2253 372
rect 2287 338 2321 372
rect 2355 338 2389 372
rect 2423 338 2457 372
rect 2491 338 2525 372
rect 2559 338 2593 372
rect 2627 338 2661 372
rect 2695 338 2729 372
rect 2763 338 2797 372
rect 2831 338 2865 372
rect 2899 338 2933 372
rect 2967 338 3001 372
rect 3035 338 3069 372
rect 3103 338 3137 372
rect 3171 338 3295 372
rect 3329 338 3453 372
rect 3487 338 3521 372
rect 3555 338 3589 372
rect 3623 338 3657 372
rect 3691 338 3725 372
rect 3759 338 3793 372
rect 3827 338 3861 372
rect 3895 338 3929 372
rect 3963 338 3997 372
rect 4031 338 4065 372
rect 4099 338 4133 372
rect 4167 338 4201 372
rect 4235 338 4269 372
rect 4303 338 4337 372
rect 4371 338 4405 372
rect 4439 338 4473 372
rect 4507 338 4541 372
rect 4575 338 4609 372
rect 4643 338 4677 372
rect 4711 338 4745 372
rect 4779 338 4813 372
rect 4847 338 4881 372
rect 4915 338 4949 372
rect 4983 338 5017 372
rect 5051 338 5085 372
rect 5119 338 5153 372
rect 5187 338 5221 372
rect 5255 338 5289 372
rect 5323 338 5357 372
rect 5391 338 5425 372
rect 5459 338 5493 372
rect 5527 338 5561 372
rect 5595 338 5629 372
rect 5663 338 5697 372
rect 5731 338 5765 372
rect 5799 338 5833 372
rect 5867 338 5901 372
rect 5935 338 5969 372
rect 6003 338 6037 372
rect 6071 338 6105 372
rect 6139 338 6173 372
rect 6207 338 6241 372
rect 6275 338 6309 372
rect 6343 338 6377 372
rect 6411 338 6445 372
rect 6479 338 6513 372
rect 6547 338 6581 372
rect 6615 338 6649 372
rect 6683 338 6834 372
rect -244 304 -210 338
rect -244 236 -210 270
rect -244 168 -210 202
rect -244 100 -210 134
rect 3295 304 3329 338
rect 3295 236 3329 270
rect 3295 168 3329 202
rect 3295 100 3329 134
rect 6834 304 6868 338
rect 6834 236 6868 270
rect 6834 168 6868 202
rect -244 32 -210 66
rect -244 -36 -210 -2
rect -244 -104 -210 -70
rect 6834 100 6868 134
rect 3295 32 3329 66
rect 3295 -36 3329 -2
rect 3295 -104 3329 -70
rect -244 -172 -210 -138
rect 6834 32 6868 66
rect 6834 -36 6868 -2
rect 6834 -104 6868 -70
rect 3295 -172 3329 -138
rect -244 -240 -210 -206
rect -244 -308 -210 -274
rect -244 -376 -210 -342
rect -244 -444 -210 -410
rect -244 -512 -210 -478
rect 6834 -172 6868 -138
rect 3295 -240 3329 -206
rect 3295 -308 3329 -274
rect 3295 -376 3329 -342
rect 3295 -444 3329 -410
rect -244 -580 -210 -546
rect 3295 -512 3329 -478
rect 6834 -240 6868 -206
rect 6834 -308 6868 -274
rect 6834 -376 6868 -342
rect 6834 -444 6868 -410
rect 3295 -580 3329 -546
rect -244 -648 -210 -614
rect -244 -716 -210 -682
rect -244 -784 -210 -750
rect 6834 -512 6868 -478
rect 6834 -580 6868 -546
rect 3295 -648 3329 -614
rect 3295 -716 3329 -682
rect 3295 -784 3329 -750
rect 6834 -648 6868 -614
rect 6834 -716 6868 -682
rect -244 -852 -210 -818
rect -244 -1026 -210 -886
rect 6834 -784 6868 -750
rect 3295 -852 3329 -818
rect 3295 -1026 3329 -886
rect 6834 -852 6868 -818
rect 6834 -1026 6868 -886
rect -244 -1060 -59 -1026
rect -25 -1060 9 -1026
rect 43 -1060 77 -1026
rect 111 -1060 145 -1026
rect 179 -1060 213 -1026
rect 247 -1060 281 -1026
rect 315 -1060 349 -1026
rect 383 -1060 417 -1026
rect 451 -1060 485 -1026
rect 519 -1060 553 -1026
rect 587 -1060 621 -1026
rect 655 -1060 689 -1026
rect 723 -1060 757 -1026
rect 791 -1060 825 -1026
rect 859 -1060 893 -1026
rect 927 -1060 961 -1026
rect 995 -1060 1029 -1026
rect 1063 -1060 1097 -1026
rect 1131 -1060 1165 -1026
rect 1199 -1060 1233 -1026
rect 1267 -1060 1301 -1026
rect 1335 -1060 1369 -1026
rect 1403 -1060 1437 -1026
rect 1471 -1060 1505 -1026
rect 1539 -1060 1573 -1026
rect 1607 -1060 1641 -1026
rect 1675 -1060 1709 -1026
rect 1743 -1060 1777 -1026
rect 1811 -1060 1845 -1026
rect 1879 -1060 1913 -1026
rect 1947 -1060 1981 -1026
rect 2015 -1060 2049 -1026
rect 2083 -1060 2117 -1026
rect 2151 -1060 2185 -1026
rect 2219 -1060 2253 -1026
rect 2287 -1060 2321 -1026
rect 2355 -1060 2389 -1026
rect 2423 -1060 2457 -1026
rect 2491 -1060 2525 -1026
rect 2559 -1060 2593 -1026
rect 2627 -1060 2661 -1026
rect 2695 -1060 2729 -1026
rect 2763 -1060 2797 -1026
rect 2831 -1060 2865 -1026
rect 2899 -1060 2933 -1026
rect 2967 -1060 3001 -1026
rect 3035 -1060 3069 -1026
rect 3103 -1060 3137 -1026
rect 3171 -1060 3453 -1026
rect 3487 -1060 3521 -1026
rect 3555 -1060 3589 -1026
rect 3623 -1060 3657 -1026
rect 3691 -1060 3725 -1026
rect 3759 -1060 3793 -1026
rect 3827 -1060 3861 -1026
rect 3895 -1060 3929 -1026
rect 3963 -1060 3997 -1026
rect 4031 -1060 4065 -1026
rect 4099 -1060 4133 -1026
rect 4167 -1060 4201 -1026
rect 4235 -1060 4269 -1026
rect 4303 -1060 4337 -1026
rect 4371 -1060 4405 -1026
rect 4439 -1060 4473 -1026
rect 4507 -1060 4541 -1026
rect 4575 -1060 4609 -1026
rect 4643 -1060 4677 -1026
rect 4711 -1060 4745 -1026
rect 4779 -1060 4813 -1026
rect 4847 -1060 4881 -1026
rect 4915 -1060 4949 -1026
rect 4983 -1060 5017 -1026
rect 5051 -1060 5085 -1026
rect 5119 -1060 5153 -1026
rect 5187 -1060 5221 -1026
rect 5255 -1060 5289 -1026
rect 5323 -1060 5357 -1026
rect 5391 -1060 5425 -1026
rect 5459 -1060 5493 -1026
rect 5527 -1060 5561 -1026
rect 5595 -1060 5629 -1026
rect 5663 -1060 5697 -1026
rect 5731 -1060 5765 -1026
rect 5799 -1060 5833 -1026
rect 5867 -1060 5901 -1026
rect 5935 -1060 5969 -1026
rect 6003 -1060 6037 -1026
rect 6071 -1060 6105 -1026
rect 6139 -1060 6173 -1026
rect 6207 -1060 6241 -1026
rect 6275 -1060 6309 -1026
rect 6343 -1060 6377 -1026
rect 6411 -1060 6445 -1026
rect 6479 -1060 6513 -1026
rect 6547 -1060 6581 -1026
rect 6615 -1060 6649 -1026
rect 6683 -1060 6868 -1026
rect -244 -1200 -210 -1060
rect -244 -1268 -210 -1234
rect 3295 -1200 3329 -1060
rect 3295 -1268 3329 -1234
rect -244 -1336 -210 -1302
rect 6834 -1200 6868 -1060
rect 6834 -1268 6868 -1234
rect -244 -1404 -210 -1370
rect -244 -1472 -210 -1438
rect 3295 -1336 3329 -1302
rect 3295 -1404 3329 -1370
rect 3295 -1472 3329 -1438
rect -244 -1540 -210 -1506
rect -244 -1608 -210 -1574
rect 6834 -1336 6868 -1302
rect 6834 -1404 6868 -1370
rect 6834 -1472 6868 -1438
rect 3295 -1540 3329 -1506
rect -244 -1676 -210 -1642
rect -244 -1744 -210 -1710
rect -244 -1812 -210 -1778
rect -244 -1880 -210 -1846
rect 3295 -1608 3329 -1574
rect 6834 -1540 6868 -1506
rect 3295 -1676 3329 -1642
rect 3295 -1744 3329 -1710
rect 3295 -1812 3329 -1778
rect 3295 -1880 3329 -1846
rect -244 -1948 -210 -1914
rect 6834 -1608 6868 -1574
rect 6834 -1676 6868 -1642
rect 6834 -1744 6868 -1710
rect 6834 -1812 6868 -1778
rect 6834 -1880 6868 -1846
rect 3295 -1948 3329 -1914
rect -244 -2016 -210 -1982
rect -244 -2084 -210 -2050
rect -244 -2152 -210 -2118
rect 6834 -1948 6868 -1914
rect 3295 -2016 3329 -1982
rect 3295 -2084 3329 -2050
rect 3295 -2152 3329 -2118
rect -244 -2220 -210 -2186
rect 6834 -2016 6868 -1982
rect 6834 -2084 6868 -2050
rect 6834 -2152 6868 -2118
rect -244 -2288 -210 -2254
rect -244 -2356 -210 -2322
rect -244 -2424 -210 -2390
rect 3295 -2220 3329 -2186
rect 3295 -2288 3329 -2254
rect 3295 -2356 3329 -2322
rect 3295 -2424 3329 -2390
rect 6834 -2220 6868 -2186
rect 6834 -2288 6868 -2254
rect 6834 -2356 6868 -2322
rect 6834 -2424 6868 -2390
rect -210 -2458 -59 -2424
rect -25 -2458 9 -2424
rect 43 -2458 77 -2424
rect 111 -2458 145 -2424
rect 179 -2458 213 -2424
rect 247 -2458 281 -2424
rect 315 -2458 349 -2424
rect 383 -2458 417 -2424
rect 451 -2458 485 -2424
rect 519 -2458 553 -2424
rect 587 -2458 621 -2424
rect 655 -2458 689 -2424
rect 723 -2458 757 -2424
rect 791 -2458 825 -2424
rect 859 -2458 893 -2424
rect 927 -2458 961 -2424
rect 995 -2458 1029 -2424
rect 1063 -2458 1097 -2424
rect 1131 -2458 1165 -2424
rect 1199 -2458 1233 -2424
rect 1267 -2458 1301 -2424
rect 1335 -2458 1369 -2424
rect 1403 -2458 1437 -2424
rect 1471 -2458 1505 -2424
rect 1539 -2458 1573 -2424
rect 1607 -2458 1641 -2424
rect 1675 -2458 1709 -2424
rect 1743 -2458 1777 -2424
rect 1811 -2458 1845 -2424
rect 1879 -2458 1913 -2424
rect 1947 -2458 1981 -2424
rect 2015 -2458 2049 -2424
rect 2083 -2458 2117 -2424
rect 2151 -2458 2185 -2424
rect 2219 -2458 2253 -2424
rect 2287 -2458 2321 -2424
rect 2355 -2458 2389 -2424
rect 2423 -2458 2457 -2424
rect 2491 -2458 2525 -2424
rect 2559 -2458 2593 -2424
rect 2627 -2458 2661 -2424
rect 2695 -2458 2729 -2424
rect 2763 -2458 2797 -2424
rect 2831 -2458 2865 -2424
rect 2899 -2458 2933 -2424
rect 2967 -2458 3001 -2424
rect 3035 -2458 3069 -2424
rect 3103 -2458 3137 -2424
rect 3171 -2458 3295 -2424
rect 3329 -2458 3453 -2424
rect 3487 -2458 3521 -2424
rect 3555 -2458 3589 -2424
rect 3623 -2458 3657 -2424
rect 3691 -2458 3725 -2424
rect 3759 -2458 3793 -2424
rect 3827 -2458 3861 -2424
rect 3895 -2458 3929 -2424
rect 3963 -2458 3997 -2424
rect 4031 -2458 4065 -2424
rect 4099 -2458 4133 -2424
rect 4167 -2458 4201 -2424
rect 4235 -2458 4269 -2424
rect 4303 -2458 4337 -2424
rect 4371 -2458 4405 -2424
rect 4439 -2458 4473 -2424
rect 4507 -2458 4541 -2424
rect 4575 -2458 4609 -2424
rect 4643 -2458 4677 -2424
rect 4711 -2458 4745 -2424
rect 4779 -2458 4813 -2424
rect 4847 -2458 4881 -2424
rect 4915 -2458 4949 -2424
rect 4983 -2458 5017 -2424
rect 5051 -2458 5085 -2424
rect 5119 -2458 5153 -2424
rect 5187 -2458 5221 -2424
rect 5255 -2458 5289 -2424
rect 5323 -2458 5357 -2424
rect 5391 -2458 5425 -2424
rect 5459 -2458 5493 -2424
rect 5527 -2458 5561 -2424
rect 5595 -2458 5629 -2424
rect 5663 -2458 5697 -2424
rect 5731 -2458 5765 -2424
rect 5799 -2458 5833 -2424
rect 5867 -2458 5901 -2424
rect 5935 -2458 5969 -2424
rect 6003 -2458 6037 -2424
rect 6071 -2458 6105 -2424
rect 6139 -2458 6173 -2424
rect 6207 -2458 6241 -2424
rect 6275 -2458 6309 -2424
rect 6343 -2458 6377 -2424
rect 6411 -2458 6445 -2424
rect 6479 -2458 6513 -2424
rect 6547 -2458 6581 -2424
rect 6615 -2458 6649 -2424
rect 6683 -2458 6834 -2424
rect -244 -2492 -210 -2458
rect -244 -2560 -210 -2526
rect -244 -2628 -210 -2594
rect -244 -2696 -210 -2662
rect 3295 -2492 3329 -2458
rect 3295 -2560 3329 -2526
rect 3295 -2628 3329 -2594
rect 3295 -2696 3329 -2662
rect 6834 -2492 6868 -2458
rect 6834 -2560 6868 -2526
rect 6834 -2628 6868 -2594
rect -244 -2764 -210 -2730
rect -244 -2832 -210 -2798
rect -244 -2900 -210 -2866
rect 6834 -2696 6868 -2662
rect 3295 -2764 3329 -2730
rect 3295 -2832 3329 -2798
rect 3295 -2900 3329 -2866
rect -244 -3041 -210 -2934
rect 6834 -2764 6868 -2730
rect 6834 -2832 6868 -2798
rect 6834 -2900 6868 -2866
rect 3295 -3041 3329 -2934
rect 6834 -3041 6868 -2934
rect -244 -3075 -59 -3041
rect -25 -3075 9 -3041
rect 43 -3075 77 -3041
rect 111 -3075 145 -3041
rect 179 -3075 213 -3041
rect 247 -3075 281 -3041
rect 315 -3075 349 -3041
rect 383 -3075 417 -3041
rect 451 -3075 485 -3041
rect 519 -3075 553 -3041
rect 587 -3075 621 -3041
rect 655 -3075 689 -3041
rect 723 -3075 757 -3041
rect 791 -3075 825 -3041
rect 859 -3075 893 -3041
rect 927 -3075 961 -3041
rect 995 -3075 1029 -3041
rect 1063 -3075 1097 -3041
rect 1131 -3075 1165 -3041
rect 1199 -3075 1233 -3041
rect 1267 -3075 1301 -3041
rect 1335 -3075 1369 -3041
rect 1403 -3075 1437 -3041
rect 1471 -3075 1505 -3041
rect 1539 -3075 1573 -3041
rect 1607 -3075 1641 -3041
rect 1675 -3075 1709 -3041
rect 1743 -3075 1777 -3041
rect 1811 -3075 1845 -3041
rect 1879 -3075 1913 -3041
rect 1947 -3075 1981 -3041
rect 2015 -3075 2049 -3041
rect 2083 -3075 2117 -3041
rect 2151 -3075 2185 -3041
rect 2219 -3075 2253 -3041
rect 2287 -3075 2321 -3041
rect 2355 -3075 2389 -3041
rect 2423 -3075 2457 -3041
rect 2491 -3075 2525 -3041
rect 2559 -3075 2593 -3041
rect 2627 -3075 2661 -3041
rect 2695 -3075 2729 -3041
rect 2763 -3075 2797 -3041
rect 2831 -3075 2865 -3041
rect 2899 -3075 2933 -3041
rect 2967 -3075 3001 -3041
rect 3035 -3075 3069 -3041
rect 3103 -3075 3137 -3041
rect 3171 -3075 3453 -3041
rect 3487 -3075 3521 -3041
rect 3555 -3075 3589 -3041
rect 3623 -3075 3657 -3041
rect 3691 -3075 3725 -3041
rect 3759 -3075 3793 -3041
rect 3827 -3075 3861 -3041
rect 3895 -3075 3929 -3041
rect 3963 -3075 3997 -3041
rect 4031 -3075 4065 -3041
rect 4099 -3075 4133 -3041
rect 4167 -3075 4201 -3041
rect 4235 -3075 4269 -3041
rect 4303 -3075 4337 -3041
rect 4371 -3075 4405 -3041
rect 4439 -3075 4473 -3041
rect 4507 -3075 4541 -3041
rect 4575 -3075 4609 -3041
rect 4643 -3075 4677 -3041
rect 4711 -3075 4745 -3041
rect 4779 -3075 4813 -3041
rect 4847 -3075 4881 -3041
rect 4915 -3075 4949 -3041
rect 4983 -3075 5017 -3041
rect 5051 -3075 5085 -3041
rect 5119 -3075 5153 -3041
rect 5187 -3075 5221 -3041
rect 5255 -3075 5289 -3041
rect 5323 -3075 5357 -3041
rect 5391 -3075 5425 -3041
rect 5459 -3075 5493 -3041
rect 5527 -3075 5561 -3041
rect 5595 -3075 5629 -3041
rect 5663 -3075 5697 -3041
rect 5731 -3075 5765 -3041
rect 5799 -3075 5833 -3041
rect 5867 -3075 5901 -3041
rect 5935 -3075 5969 -3041
rect 6003 -3075 6037 -3041
rect 6071 -3075 6105 -3041
rect 6139 -3075 6173 -3041
rect 6207 -3075 6241 -3041
rect 6275 -3075 6309 -3041
rect 6343 -3075 6377 -3041
rect 6411 -3075 6445 -3041
rect 6479 -3075 6513 -3041
rect 6547 -3075 6581 -3041
rect 6615 -3075 6649 -3041
rect 6683 -3075 6868 -3041
<< psubdiffcont >>
rect -59 955 -25 989
rect 9 955 43 989
rect 77 955 111 989
rect 145 955 179 989
rect 213 955 247 989
rect 281 955 315 989
rect 349 955 383 989
rect 417 955 451 989
rect 485 955 519 989
rect 553 955 587 989
rect 621 955 655 989
rect 689 955 723 989
rect 757 955 791 989
rect 825 955 859 989
rect 893 955 927 989
rect 961 955 995 989
rect 1029 955 1063 989
rect 1097 955 1131 989
rect 1165 955 1199 989
rect 1233 955 1267 989
rect 1301 955 1335 989
rect 1369 955 1403 989
rect 1437 955 1471 989
rect 1505 955 1539 989
rect 1573 955 1607 989
rect 1641 955 1675 989
rect 1709 955 1743 989
rect 1777 955 1811 989
rect 1845 955 1879 989
rect 1913 955 1947 989
rect 1981 955 2015 989
rect 2049 955 2083 989
rect 2117 955 2151 989
rect 2185 955 2219 989
rect 2253 955 2287 989
rect 2321 955 2355 989
rect 2389 955 2423 989
rect 2457 955 2491 989
rect 2525 955 2559 989
rect 2593 955 2627 989
rect 2661 955 2695 989
rect 2729 955 2763 989
rect 2797 955 2831 989
rect 2865 955 2899 989
rect 2933 955 2967 989
rect 3001 955 3035 989
rect 3069 955 3103 989
rect 3137 955 3171 989
rect 3453 955 3487 989
rect 3521 955 3555 989
rect 3589 955 3623 989
rect 3657 955 3691 989
rect 3725 955 3759 989
rect 3793 955 3827 989
rect 3861 955 3895 989
rect 3929 955 3963 989
rect 3997 955 4031 989
rect 4065 955 4099 989
rect 4133 955 4167 989
rect 4201 955 4235 989
rect 4269 955 4303 989
rect 4337 955 4371 989
rect 4405 955 4439 989
rect 4473 955 4507 989
rect 4541 955 4575 989
rect 4609 955 4643 989
rect 4677 955 4711 989
rect 4745 955 4779 989
rect 4813 955 4847 989
rect 4881 955 4915 989
rect 4949 955 4983 989
rect 5017 955 5051 989
rect 5085 955 5119 989
rect 5153 955 5187 989
rect 5221 955 5255 989
rect 5289 955 5323 989
rect 5357 955 5391 989
rect 5425 955 5459 989
rect 5493 955 5527 989
rect 5561 955 5595 989
rect 5629 955 5663 989
rect 5697 955 5731 989
rect 5765 955 5799 989
rect 5833 955 5867 989
rect 5901 955 5935 989
rect 5969 955 6003 989
rect 6037 955 6071 989
rect 6105 955 6139 989
rect 6173 955 6207 989
rect 6241 955 6275 989
rect 6309 955 6343 989
rect 6377 955 6411 989
rect 6445 955 6479 989
rect 6513 955 6547 989
rect 6581 955 6615 989
rect 6649 955 6683 989
rect -244 814 -210 848
rect -244 746 -210 780
rect -244 678 -210 712
rect -244 610 -210 644
rect 3295 814 3329 848
rect 3295 746 3329 780
rect 3295 678 3329 712
rect 3295 610 3329 644
rect 6834 814 6868 848
rect 6834 746 6868 780
rect 6834 678 6868 712
rect -244 542 -210 576
rect -244 474 -210 508
rect -244 406 -210 440
rect 6834 610 6868 644
rect 3295 542 3329 576
rect 3295 474 3329 508
rect 3295 406 3329 440
rect 6834 542 6868 576
rect 6834 474 6868 508
rect 6834 406 6868 440
rect -244 338 -210 372
rect -59 338 -25 372
rect 9 338 43 372
rect 77 338 111 372
rect 145 338 179 372
rect 213 338 247 372
rect 281 338 315 372
rect 349 338 383 372
rect 417 338 451 372
rect 485 338 519 372
rect 553 338 587 372
rect 621 338 655 372
rect 689 338 723 372
rect 757 338 791 372
rect 825 338 859 372
rect 893 338 927 372
rect 961 338 995 372
rect 1029 338 1063 372
rect 1097 338 1131 372
rect 1165 338 1199 372
rect 1233 338 1267 372
rect 1301 338 1335 372
rect 1369 338 1403 372
rect 1437 338 1471 372
rect 1505 338 1539 372
rect 1573 338 1607 372
rect 1641 338 1675 372
rect 1709 338 1743 372
rect 1777 338 1811 372
rect 1845 338 1879 372
rect 1913 338 1947 372
rect 1981 338 2015 372
rect 2049 338 2083 372
rect 2117 338 2151 372
rect 2185 338 2219 372
rect 2253 338 2287 372
rect 2321 338 2355 372
rect 2389 338 2423 372
rect 2457 338 2491 372
rect 2525 338 2559 372
rect 2593 338 2627 372
rect 2661 338 2695 372
rect 2729 338 2763 372
rect 2797 338 2831 372
rect 2865 338 2899 372
rect 2933 338 2967 372
rect 3001 338 3035 372
rect 3069 338 3103 372
rect 3137 338 3171 372
rect 3295 338 3329 372
rect 3453 338 3487 372
rect 3521 338 3555 372
rect 3589 338 3623 372
rect 3657 338 3691 372
rect 3725 338 3759 372
rect 3793 338 3827 372
rect 3861 338 3895 372
rect 3929 338 3963 372
rect 3997 338 4031 372
rect 4065 338 4099 372
rect 4133 338 4167 372
rect 4201 338 4235 372
rect 4269 338 4303 372
rect 4337 338 4371 372
rect 4405 338 4439 372
rect 4473 338 4507 372
rect 4541 338 4575 372
rect 4609 338 4643 372
rect 4677 338 4711 372
rect 4745 338 4779 372
rect 4813 338 4847 372
rect 4881 338 4915 372
rect 4949 338 4983 372
rect 5017 338 5051 372
rect 5085 338 5119 372
rect 5153 338 5187 372
rect 5221 338 5255 372
rect 5289 338 5323 372
rect 5357 338 5391 372
rect 5425 338 5459 372
rect 5493 338 5527 372
rect 5561 338 5595 372
rect 5629 338 5663 372
rect 5697 338 5731 372
rect 5765 338 5799 372
rect 5833 338 5867 372
rect 5901 338 5935 372
rect 5969 338 6003 372
rect 6037 338 6071 372
rect 6105 338 6139 372
rect 6173 338 6207 372
rect 6241 338 6275 372
rect 6309 338 6343 372
rect 6377 338 6411 372
rect 6445 338 6479 372
rect 6513 338 6547 372
rect 6581 338 6615 372
rect 6649 338 6683 372
rect 6834 338 6868 372
rect -244 270 -210 304
rect -244 202 -210 236
rect -244 134 -210 168
rect 3295 270 3329 304
rect 3295 202 3329 236
rect 3295 134 3329 168
rect -244 66 -210 100
rect 6834 270 6868 304
rect 6834 202 6868 236
rect 6834 134 6868 168
rect -244 -2 -210 32
rect -244 -70 -210 -36
rect -244 -138 -210 -104
rect 3295 66 3329 100
rect 3295 -2 3329 32
rect 3295 -70 3329 -36
rect -244 -206 -210 -172
rect 3295 -138 3329 -104
rect 6834 66 6868 100
rect 6834 -2 6868 32
rect 6834 -70 6868 -36
rect -244 -274 -210 -240
rect -244 -342 -210 -308
rect -244 -410 -210 -376
rect -244 -478 -210 -444
rect 3295 -206 3329 -172
rect 6834 -138 6868 -104
rect 3295 -274 3329 -240
rect 3295 -342 3329 -308
rect 3295 -410 3329 -376
rect 3295 -478 3329 -444
rect -244 -546 -210 -512
rect -244 -614 -210 -580
rect 6834 -206 6868 -172
rect 6834 -274 6868 -240
rect 6834 -342 6868 -308
rect 6834 -410 6868 -376
rect 6834 -478 6868 -444
rect 3295 -546 3329 -512
rect -244 -682 -210 -648
rect -244 -750 -210 -716
rect 3295 -614 3329 -580
rect 6834 -546 6868 -512
rect 3295 -682 3329 -648
rect 3295 -750 3329 -716
rect -244 -818 -210 -784
rect 6834 -614 6868 -580
rect 6834 -682 6868 -648
rect 6834 -750 6868 -716
rect -244 -886 -210 -852
rect 3295 -818 3329 -784
rect 3295 -886 3329 -852
rect 6834 -818 6868 -784
rect 6834 -886 6868 -852
rect -59 -1060 -25 -1026
rect 9 -1060 43 -1026
rect 77 -1060 111 -1026
rect 145 -1060 179 -1026
rect 213 -1060 247 -1026
rect 281 -1060 315 -1026
rect 349 -1060 383 -1026
rect 417 -1060 451 -1026
rect 485 -1060 519 -1026
rect 553 -1060 587 -1026
rect 621 -1060 655 -1026
rect 689 -1060 723 -1026
rect 757 -1060 791 -1026
rect 825 -1060 859 -1026
rect 893 -1060 927 -1026
rect 961 -1060 995 -1026
rect 1029 -1060 1063 -1026
rect 1097 -1060 1131 -1026
rect 1165 -1060 1199 -1026
rect 1233 -1060 1267 -1026
rect 1301 -1060 1335 -1026
rect 1369 -1060 1403 -1026
rect 1437 -1060 1471 -1026
rect 1505 -1060 1539 -1026
rect 1573 -1060 1607 -1026
rect 1641 -1060 1675 -1026
rect 1709 -1060 1743 -1026
rect 1777 -1060 1811 -1026
rect 1845 -1060 1879 -1026
rect 1913 -1060 1947 -1026
rect 1981 -1060 2015 -1026
rect 2049 -1060 2083 -1026
rect 2117 -1060 2151 -1026
rect 2185 -1060 2219 -1026
rect 2253 -1060 2287 -1026
rect 2321 -1060 2355 -1026
rect 2389 -1060 2423 -1026
rect 2457 -1060 2491 -1026
rect 2525 -1060 2559 -1026
rect 2593 -1060 2627 -1026
rect 2661 -1060 2695 -1026
rect 2729 -1060 2763 -1026
rect 2797 -1060 2831 -1026
rect 2865 -1060 2899 -1026
rect 2933 -1060 2967 -1026
rect 3001 -1060 3035 -1026
rect 3069 -1060 3103 -1026
rect 3137 -1060 3171 -1026
rect 3453 -1060 3487 -1026
rect 3521 -1060 3555 -1026
rect 3589 -1060 3623 -1026
rect 3657 -1060 3691 -1026
rect 3725 -1060 3759 -1026
rect 3793 -1060 3827 -1026
rect 3861 -1060 3895 -1026
rect 3929 -1060 3963 -1026
rect 3997 -1060 4031 -1026
rect 4065 -1060 4099 -1026
rect 4133 -1060 4167 -1026
rect 4201 -1060 4235 -1026
rect 4269 -1060 4303 -1026
rect 4337 -1060 4371 -1026
rect 4405 -1060 4439 -1026
rect 4473 -1060 4507 -1026
rect 4541 -1060 4575 -1026
rect 4609 -1060 4643 -1026
rect 4677 -1060 4711 -1026
rect 4745 -1060 4779 -1026
rect 4813 -1060 4847 -1026
rect 4881 -1060 4915 -1026
rect 4949 -1060 4983 -1026
rect 5017 -1060 5051 -1026
rect 5085 -1060 5119 -1026
rect 5153 -1060 5187 -1026
rect 5221 -1060 5255 -1026
rect 5289 -1060 5323 -1026
rect 5357 -1060 5391 -1026
rect 5425 -1060 5459 -1026
rect 5493 -1060 5527 -1026
rect 5561 -1060 5595 -1026
rect 5629 -1060 5663 -1026
rect 5697 -1060 5731 -1026
rect 5765 -1060 5799 -1026
rect 5833 -1060 5867 -1026
rect 5901 -1060 5935 -1026
rect 5969 -1060 6003 -1026
rect 6037 -1060 6071 -1026
rect 6105 -1060 6139 -1026
rect 6173 -1060 6207 -1026
rect 6241 -1060 6275 -1026
rect 6309 -1060 6343 -1026
rect 6377 -1060 6411 -1026
rect 6445 -1060 6479 -1026
rect 6513 -1060 6547 -1026
rect 6581 -1060 6615 -1026
rect 6649 -1060 6683 -1026
rect -244 -1234 -210 -1200
rect -244 -1302 -210 -1268
rect 3295 -1234 3329 -1200
rect 3295 -1302 3329 -1268
rect 6834 -1234 6868 -1200
rect -244 -1370 -210 -1336
rect -244 -1438 -210 -1404
rect -244 -1506 -210 -1472
rect 6834 -1302 6868 -1268
rect 3295 -1370 3329 -1336
rect 3295 -1438 3329 -1404
rect -244 -1574 -210 -1540
rect 3295 -1506 3329 -1472
rect 6834 -1370 6868 -1336
rect 6834 -1438 6868 -1404
rect 3295 -1574 3329 -1540
rect -244 -1642 -210 -1608
rect -244 -1710 -210 -1676
rect -244 -1778 -210 -1744
rect -244 -1846 -210 -1812
rect -244 -1914 -210 -1880
rect 6834 -1506 6868 -1472
rect 6834 -1574 6868 -1540
rect 3295 -1642 3329 -1608
rect 3295 -1710 3329 -1676
rect 3295 -1778 3329 -1744
rect 3295 -1846 3329 -1812
rect -244 -1982 -210 -1948
rect 3295 -1914 3329 -1880
rect 6834 -1642 6868 -1608
rect 6834 -1710 6868 -1676
rect 6834 -1778 6868 -1744
rect 6834 -1846 6868 -1812
rect -244 -2050 -210 -2016
rect -244 -2118 -210 -2084
rect -244 -2186 -210 -2152
rect 3295 -1982 3329 -1948
rect 6834 -1914 6868 -1880
rect 3295 -2050 3329 -2016
rect 3295 -2118 3329 -2084
rect 3295 -2186 3329 -2152
rect 6834 -1982 6868 -1948
rect 6834 -2050 6868 -2016
rect 6834 -2118 6868 -2084
rect -244 -2254 -210 -2220
rect -244 -2322 -210 -2288
rect -244 -2390 -210 -2356
rect 6834 -2186 6868 -2152
rect 3295 -2254 3329 -2220
rect 3295 -2322 3329 -2288
rect 3295 -2390 3329 -2356
rect 6834 -2254 6868 -2220
rect 6834 -2322 6868 -2288
rect 6834 -2390 6868 -2356
rect -244 -2458 -210 -2424
rect -59 -2458 -25 -2424
rect 9 -2458 43 -2424
rect 77 -2458 111 -2424
rect 145 -2458 179 -2424
rect 213 -2458 247 -2424
rect 281 -2458 315 -2424
rect 349 -2458 383 -2424
rect 417 -2458 451 -2424
rect 485 -2458 519 -2424
rect 553 -2458 587 -2424
rect 621 -2458 655 -2424
rect 689 -2458 723 -2424
rect 757 -2458 791 -2424
rect 825 -2458 859 -2424
rect 893 -2458 927 -2424
rect 961 -2458 995 -2424
rect 1029 -2458 1063 -2424
rect 1097 -2458 1131 -2424
rect 1165 -2458 1199 -2424
rect 1233 -2458 1267 -2424
rect 1301 -2458 1335 -2424
rect 1369 -2458 1403 -2424
rect 1437 -2458 1471 -2424
rect 1505 -2458 1539 -2424
rect 1573 -2458 1607 -2424
rect 1641 -2458 1675 -2424
rect 1709 -2458 1743 -2424
rect 1777 -2458 1811 -2424
rect 1845 -2458 1879 -2424
rect 1913 -2458 1947 -2424
rect 1981 -2458 2015 -2424
rect 2049 -2458 2083 -2424
rect 2117 -2458 2151 -2424
rect 2185 -2458 2219 -2424
rect 2253 -2458 2287 -2424
rect 2321 -2458 2355 -2424
rect 2389 -2458 2423 -2424
rect 2457 -2458 2491 -2424
rect 2525 -2458 2559 -2424
rect 2593 -2458 2627 -2424
rect 2661 -2458 2695 -2424
rect 2729 -2458 2763 -2424
rect 2797 -2458 2831 -2424
rect 2865 -2458 2899 -2424
rect 2933 -2458 2967 -2424
rect 3001 -2458 3035 -2424
rect 3069 -2458 3103 -2424
rect 3137 -2458 3171 -2424
rect 3295 -2458 3329 -2424
rect 3453 -2458 3487 -2424
rect 3521 -2458 3555 -2424
rect 3589 -2458 3623 -2424
rect 3657 -2458 3691 -2424
rect 3725 -2458 3759 -2424
rect 3793 -2458 3827 -2424
rect 3861 -2458 3895 -2424
rect 3929 -2458 3963 -2424
rect 3997 -2458 4031 -2424
rect 4065 -2458 4099 -2424
rect 4133 -2458 4167 -2424
rect 4201 -2458 4235 -2424
rect 4269 -2458 4303 -2424
rect 4337 -2458 4371 -2424
rect 4405 -2458 4439 -2424
rect 4473 -2458 4507 -2424
rect 4541 -2458 4575 -2424
rect 4609 -2458 4643 -2424
rect 4677 -2458 4711 -2424
rect 4745 -2458 4779 -2424
rect 4813 -2458 4847 -2424
rect 4881 -2458 4915 -2424
rect 4949 -2458 4983 -2424
rect 5017 -2458 5051 -2424
rect 5085 -2458 5119 -2424
rect 5153 -2458 5187 -2424
rect 5221 -2458 5255 -2424
rect 5289 -2458 5323 -2424
rect 5357 -2458 5391 -2424
rect 5425 -2458 5459 -2424
rect 5493 -2458 5527 -2424
rect 5561 -2458 5595 -2424
rect 5629 -2458 5663 -2424
rect 5697 -2458 5731 -2424
rect 5765 -2458 5799 -2424
rect 5833 -2458 5867 -2424
rect 5901 -2458 5935 -2424
rect 5969 -2458 6003 -2424
rect 6037 -2458 6071 -2424
rect 6105 -2458 6139 -2424
rect 6173 -2458 6207 -2424
rect 6241 -2458 6275 -2424
rect 6309 -2458 6343 -2424
rect 6377 -2458 6411 -2424
rect 6445 -2458 6479 -2424
rect 6513 -2458 6547 -2424
rect 6581 -2458 6615 -2424
rect 6649 -2458 6683 -2424
rect 6834 -2458 6868 -2424
rect -244 -2526 -210 -2492
rect -244 -2594 -210 -2560
rect -244 -2662 -210 -2628
rect 3295 -2526 3329 -2492
rect 3295 -2594 3329 -2560
rect 3295 -2662 3329 -2628
rect -244 -2730 -210 -2696
rect 6834 -2526 6868 -2492
rect 6834 -2594 6868 -2560
rect 6834 -2662 6868 -2628
rect -244 -2798 -210 -2764
rect -244 -2866 -210 -2832
rect -244 -2934 -210 -2900
rect 3295 -2730 3329 -2696
rect 3295 -2798 3329 -2764
rect 3295 -2866 3329 -2832
rect 3295 -2934 3329 -2900
rect 6834 -2730 6868 -2696
rect 6834 -2798 6868 -2764
rect 6834 -2866 6868 -2832
rect 6834 -2934 6868 -2900
rect -59 -3075 -25 -3041
rect 9 -3075 43 -3041
rect 77 -3075 111 -3041
rect 145 -3075 179 -3041
rect 213 -3075 247 -3041
rect 281 -3075 315 -3041
rect 349 -3075 383 -3041
rect 417 -3075 451 -3041
rect 485 -3075 519 -3041
rect 553 -3075 587 -3041
rect 621 -3075 655 -3041
rect 689 -3075 723 -3041
rect 757 -3075 791 -3041
rect 825 -3075 859 -3041
rect 893 -3075 927 -3041
rect 961 -3075 995 -3041
rect 1029 -3075 1063 -3041
rect 1097 -3075 1131 -3041
rect 1165 -3075 1199 -3041
rect 1233 -3075 1267 -3041
rect 1301 -3075 1335 -3041
rect 1369 -3075 1403 -3041
rect 1437 -3075 1471 -3041
rect 1505 -3075 1539 -3041
rect 1573 -3075 1607 -3041
rect 1641 -3075 1675 -3041
rect 1709 -3075 1743 -3041
rect 1777 -3075 1811 -3041
rect 1845 -3075 1879 -3041
rect 1913 -3075 1947 -3041
rect 1981 -3075 2015 -3041
rect 2049 -3075 2083 -3041
rect 2117 -3075 2151 -3041
rect 2185 -3075 2219 -3041
rect 2253 -3075 2287 -3041
rect 2321 -3075 2355 -3041
rect 2389 -3075 2423 -3041
rect 2457 -3075 2491 -3041
rect 2525 -3075 2559 -3041
rect 2593 -3075 2627 -3041
rect 2661 -3075 2695 -3041
rect 2729 -3075 2763 -3041
rect 2797 -3075 2831 -3041
rect 2865 -3075 2899 -3041
rect 2933 -3075 2967 -3041
rect 3001 -3075 3035 -3041
rect 3069 -3075 3103 -3041
rect 3137 -3075 3171 -3041
rect 3453 -3075 3487 -3041
rect 3521 -3075 3555 -3041
rect 3589 -3075 3623 -3041
rect 3657 -3075 3691 -3041
rect 3725 -3075 3759 -3041
rect 3793 -3075 3827 -3041
rect 3861 -3075 3895 -3041
rect 3929 -3075 3963 -3041
rect 3997 -3075 4031 -3041
rect 4065 -3075 4099 -3041
rect 4133 -3075 4167 -3041
rect 4201 -3075 4235 -3041
rect 4269 -3075 4303 -3041
rect 4337 -3075 4371 -3041
rect 4405 -3075 4439 -3041
rect 4473 -3075 4507 -3041
rect 4541 -3075 4575 -3041
rect 4609 -3075 4643 -3041
rect 4677 -3075 4711 -3041
rect 4745 -3075 4779 -3041
rect 4813 -3075 4847 -3041
rect 4881 -3075 4915 -3041
rect 4949 -3075 4983 -3041
rect 5017 -3075 5051 -3041
rect 5085 -3075 5119 -3041
rect 5153 -3075 5187 -3041
rect 5221 -3075 5255 -3041
rect 5289 -3075 5323 -3041
rect 5357 -3075 5391 -3041
rect 5425 -3075 5459 -3041
rect 5493 -3075 5527 -3041
rect 5561 -3075 5595 -3041
rect 5629 -3075 5663 -3041
rect 5697 -3075 5731 -3041
rect 5765 -3075 5799 -3041
rect 5833 -3075 5867 -3041
rect 5901 -3075 5935 -3041
rect 5969 -3075 6003 -3041
rect 6037 -3075 6071 -3041
rect 6105 -3075 6139 -3041
rect 6173 -3075 6207 -3041
rect 6241 -3075 6275 -3041
rect 6309 -3075 6343 -3041
rect 6377 -3075 6411 -3041
rect 6445 -3075 6479 -3041
rect 6513 -3075 6547 -3041
rect 6581 -3075 6615 -3041
rect 6649 -3075 6683 -3041
<< poly >>
rect -84 890 116 906
rect -84 856 -35 890
rect -1 856 33 890
rect 67 856 116 890
rect -84 818 116 856
rect 421 890 621 906
rect 421 856 470 890
rect 504 856 538 890
rect 572 856 621 890
rect 421 818 621 856
rect 679 890 879 906
rect 679 856 728 890
rect 762 856 796 890
rect 830 856 879 890
rect 679 818 879 856
rect 1184 890 1384 906
rect 1184 856 1233 890
rect 1267 856 1301 890
rect 1335 856 1384 890
rect 1184 818 1384 856
rect 1442 890 1642 906
rect 1442 856 1491 890
rect 1525 856 1559 890
rect 1593 856 1642 890
rect 1442 818 1642 856
rect 1700 890 1900 906
rect 1700 856 1749 890
rect 1783 856 1817 890
rect 1851 856 1900 890
rect 1700 818 1900 856
rect 2205 890 2405 906
rect 2205 856 2254 890
rect 2288 856 2322 890
rect 2356 856 2405 890
rect 2205 818 2405 856
rect 2463 890 2663 906
rect 2463 856 2512 890
rect 2546 856 2580 890
rect 2614 856 2663 890
rect 2463 818 2663 856
rect 2969 890 3169 906
rect 2969 856 3018 890
rect 3052 856 3086 890
rect 3120 856 3169 890
rect 2969 818 3169 856
rect 3455 890 3655 906
rect 3455 856 3504 890
rect 3538 856 3572 890
rect 3606 856 3655 890
rect 3455 818 3655 856
rect 3961 890 4161 906
rect 3961 856 4010 890
rect 4044 856 4078 890
rect 4112 856 4161 890
rect 3961 818 4161 856
rect 4219 890 4419 906
rect 4219 856 4268 890
rect 4302 856 4336 890
rect 4370 856 4419 890
rect 4219 818 4419 856
rect 4724 890 4924 906
rect 4724 856 4773 890
rect 4807 856 4841 890
rect 4875 856 4924 890
rect 4724 818 4924 856
rect 4982 890 5182 906
rect 4982 856 5031 890
rect 5065 856 5099 890
rect 5133 856 5182 890
rect 4982 818 5182 856
rect 5240 890 5440 906
rect 5240 856 5289 890
rect 5323 856 5357 890
rect 5391 856 5440 890
rect 5240 818 5440 856
rect 5745 890 5945 906
rect 5745 856 5794 890
rect 5828 856 5862 890
rect 5896 856 5945 890
rect 5745 818 5945 856
rect 6003 890 6203 906
rect 6003 856 6052 890
rect 6086 856 6120 890
rect 6154 856 6203 890
rect 6003 818 6203 856
rect 6508 890 6708 906
rect 6508 856 6557 890
rect 6591 856 6625 890
rect 6659 856 6708 890
rect 6508 818 6708 856
rect -84 592 116 618
rect 421 592 621 618
rect 679 592 879 618
rect 1184 592 1384 618
rect 1442 592 1642 618
rect 1700 592 1900 618
rect 2205 592 2405 618
rect 2463 592 2663 618
rect 2969 592 3169 618
rect 3455 592 3655 618
rect 3961 592 4161 618
rect 4219 592 4419 618
rect 4724 592 4924 618
rect 4982 592 5182 618
rect 5240 592 5440 618
rect 5745 592 5945 618
rect 6003 592 6203 618
rect 6508 592 6708 618
rect -84 92 116 118
rect 421 92 621 118
rect 679 92 879 118
rect 1184 92 1384 118
rect 1442 92 1642 118
rect 1700 92 1900 118
rect 2205 92 2405 118
rect 2463 92 2663 118
rect 2969 92 3169 118
rect 3455 92 3655 118
rect 3961 92 4161 118
rect 4219 92 4419 118
rect 4724 92 4924 118
rect 4982 92 5182 118
rect 5240 92 5440 118
rect 5745 92 5945 118
rect 6003 92 6203 118
rect 6508 92 6708 118
rect -84 -146 116 -108
rect -84 -180 -35 -146
rect -1 -180 33 -146
rect 67 -180 116 -146
rect -84 -196 116 -180
rect 421 -146 621 -108
rect 421 -180 470 -146
rect 504 -180 538 -146
rect 572 -180 621 -146
rect 421 -196 621 -180
rect 679 -146 879 -108
rect 679 -180 728 -146
rect 762 -180 796 -146
rect 830 -180 879 -146
rect 679 -196 879 -180
rect 1184 -146 1384 -108
rect 1184 -180 1233 -146
rect 1267 -180 1301 -146
rect 1335 -180 1384 -146
rect 1184 -196 1384 -180
rect 1442 -146 1642 -108
rect 1442 -180 1491 -146
rect 1525 -180 1559 -146
rect 1593 -180 1642 -146
rect 1442 -196 1642 -180
rect 1700 -146 1900 -108
rect 1700 -180 1749 -146
rect 1783 -180 1817 -146
rect 1851 -180 1900 -146
rect 1700 -196 1900 -180
rect 2205 -146 2405 -108
rect 2205 -180 2254 -146
rect 2288 -180 2322 -146
rect 2356 -180 2405 -146
rect 2205 -196 2405 -180
rect 2463 -146 2663 -108
rect 2463 -180 2512 -146
rect 2546 -180 2580 -146
rect 2614 -180 2663 -146
rect 2463 -196 2663 -180
rect 2969 -146 3169 -108
rect 2969 -180 3018 -146
rect 3052 -180 3086 -146
rect 3120 -180 3169 -146
rect 2969 -196 3169 -180
rect 3455 -146 3655 -108
rect 3455 -180 3504 -146
rect 3538 -180 3572 -146
rect 3606 -180 3655 -146
rect 3455 -196 3655 -180
rect 3961 -146 4161 -108
rect 3961 -180 4010 -146
rect 4044 -180 4078 -146
rect 4112 -180 4161 -146
rect 3961 -196 4161 -180
rect 4219 -146 4419 -108
rect 4219 -180 4268 -146
rect 4302 -180 4336 -146
rect 4370 -180 4419 -146
rect 4219 -196 4419 -180
rect 4724 -146 4924 -108
rect 4724 -180 4773 -146
rect 4807 -180 4841 -146
rect 4875 -180 4924 -146
rect 4724 -196 4924 -180
rect 4982 -146 5182 -108
rect 4982 -180 5031 -146
rect 5065 -180 5099 -146
rect 5133 -180 5182 -146
rect 4982 -196 5182 -180
rect 5240 -146 5440 -108
rect 5240 -180 5289 -146
rect 5323 -180 5357 -146
rect 5391 -180 5440 -146
rect 5240 -196 5440 -180
rect 5745 -146 5945 -108
rect 5745 -180 5794 -146
rect 5828 -180 5862 -146
rect 5896 -180 5945 -146
rect 5745 -196 5945 -180
rect 6003 -146 6203 -108
rect 6003 -180 6052 -146
rect 6086 -180 6120 -146
rect 6154 -180 6203 -146
rect 6003 -196 6203 -180
rect 6508 -146 6708 -108
rect 6508 -180 6557 -146
rect 6591 -180 6625 -146
rect 6659 -180 6708 -146
rect 6508 -196 6708 -180
rect -84 -509 116 -493
rect -84 -543 -35 -509
rect -1 -543 33 -509
rect 67 -543 116 -509
rect -84 -581 116 -543
rect 421 -509 621 -493
rect 421 -543 470 -509
rect 504 -543 538 -509
rect 572 -543 621 -509
rect 421 -581 621 -543
rect 679 -509 879 -493
rect 679 -543 728 -509
rect 762 -543 796 -509
rect 830 -543 879 -509
rect 679 -581 879 -543
rect 1184 -509 1384 -493
rect 1184 -543 1233 -509
rect 1267 -543 1301 -509
rect 1335 -543 1384 -509
rect 1184 -581 1384 -543
rect 1442 -509 1642 -493
rect 1442 -543 1491 -509
rect 1525 -543 1559 -509
rect 1593 -543 1642 -509
rect 1442 -581 1642 -543
rect 1700 -509 1900 -493
rect 1700 -543 1749 -509
rect 1783 -543 1817 -509
rect 1851 -543 1900 -509
rect 1700 -581 1900 -543
rect 2205 -509 2405 -493
rect 2205 -543 2254 -509
rect 2288 -543 2322 -509
rect 2356 -543 2405 -509
rect 2205 -581 2405 -543
rect 2463 -509 2663 -493
rect 2463 -543 2512 -509
rect 2546 -543 2580 -509
rect 2614 -543 2663 -509
rect 2463 -581 2663 -543
rect 2969 -509 3169 -493
rect 2969 -543 3018 -509
rect 3052 -543 3086 -509
rect 3120 -543 3169 -509
rect 2969 -581 3169 -543
rect 3455 -509 3655 -493
rect 3455 -543 3504 -509
rect 3538 -543 3572 -509
rect 3606 -543 3655 -509
rect 3455 -581 3655 -543
rect 3961 -509 4161 -493
rect 3961 -543 4010 -509
rect 4044 -543 4078 -509
rect 4112 -543 4161 -509
rect 3961 -581 4161 -543
rect 4219 -509 4419 -493
rect 4219 -543 4268 -509
rect 4302 -543 4336 -509
rect 4370 -543 4419 -509
rect 4219 -581 4419 -543
rect 4724 -509 4924 -493
rect 4724 -543 4773 -509
rect 4807 -543 4841 -509
rect 4875 -543 4924 -509
rect 4724 -581 4924 -543
rect 4982 -509 5182 -493
rect 4982 -543 5031 -509
rect 5065 -543 5099 -509
rect 5133 -543 5182 -509
rect 4982 -581 5182 -543
rect 5240 -509 5440 -493
rect 5240 -543 5289 -509
rect 5323 -543 5357 -509
rect 5391 -543 5440 -509
rect 5240 -581 5440 -543
rect 5745 -509 5945 -493
rect 5745 -543 5794 -509
rect 5828 -543 5862 -509
rect 5896 -543 5945 -509
rect 5745 -581 5945 -543
rect 6003 -509 6203 -493
rect 6003 -543 6052 -509
rect 6086 -543 6120 -509
rect 6154 -543 6203 -509
rect 6003 -581 6203 -543
rect 6508 -509 6708 -493
rect 6508 -543 6557 -509
rect 6591 -543 6625 -509
rect 6659 -543 6708 -509
rect 6508 -581 6708 -543
rect -84 -807 116 -781
rect 421 -807 621 -781
rect 679 -807 879 -781
rect 1184 -807 1384 -781
rect 1442 -807 1642 -781
rect 1700 -807 1900 -781
rect 2205 -807 2405 -781
rect 2463 -807 2663 -781
rect 2969 -807 3169 -781
rect 3455 -807 3655 -781
rect 3961 -807 4161 -781
rect 4219 -807 4419 -781
rect 4724 -807 4924 -781
rect 4982 -807 5182 -781
rect 5240 -807 5440 -781
rect 5745 -807 5945 -781
rect 6003 -807 6203 -781
rect 6508 -807 6708 -781
rect -84 -1305 116 -1279
rect 421 -1305 621 -1279
rect 679 -1305 879 -1279
rect 1184 -1305 1384 -1279
rect 1442 -1305 1642 -1279
rect 1700 -1305 1900 -1279
rect 2205 -1305 2405 -1279
rect 2463 -1305 2663 -1279
rect 2969 -1305 3169 -1279
rect 3455 -1305 3655 -1279
rect 3961 -1305 4161 -1279
rect 4219 -1305 4419 -1279
rect 4724 -1305 4924 -1279
rect 4982 -1305 5182 -1279
rect 5240 -1305 5440 -1279
rect 5745 -1305 5945 -1279
rect 6003 -1305 6203 -1279
rect 6508 -1305 6708 -1279
rect -84 -1543 116 -1505
rect -84 -1577 -35 -1543
rect -1 -1577 33 -1543
rect 67 -1577 116 -1543
rect -84 -1593 116 -1577
rect 421 -1543 621 -1505
rect 421 -1577 470 -1543
rect 504 -1577 538 -1543
rect 572 -1577 621 -1543
rect 421 -1593 621 -1577
rect 679 -1543 879 -1505
rect 679 -1577 728 -1543
rect 762 -1577 796 -1543
rect 830 -1577 879 -1543
rect 679 -1593 879 -1577
rect 1184 -1543 1384 -1505
rect 1184 -1577 1233 -1543
rect 1267 -1577 1301 -1543
rect 1335 -1577 1384 -1543
rect 1184 -1593 1384 -1577
rect 1442 -1543 1642 -1505
rect 1442 -1577 1491 -1543
rect 1525 -1577 1559 -1543
rect 1593 -1577 1642 -1543
rect 1442 -1593 1642 -1577
rect 1700 -1543 1900 -1505
rect 1700 -1577 1749 -1543
rect 1783 -1577 1817 -1543
rect 1851 -1577 1900 -1543
rect 1700 -1593 1900 -1577
rect 2205 -1543 2405 -1505
rect 2205 -1577 2254 -1543
rect 2288 -1577 2322 -1543
rect 2356 -1577 2405 -1543
rect 2205 -1593 2405 -1577
rect 2463 -1543 2663 -1505
rect 2463 -1577 2512 -1543
rect 2546 -1577 2580 -1543
rect 2614 -1577 2663 -1543
rect 2463 -1593 2663 -1577
rect 2969 -1543 3169 -1505
rect 2969 -1577 3018 -1543
rect 3052 -1577 3086 -1543
rect 3120 -1577 3169 -1543
rect 2969 -1593 3169 -1577
rect 3455 -1543 3655 -1505
rect 3455 -1577 3504 -1543
rect 3538 -1577 3572 -1543
rect 3606 -1577 3655 -1543
rect 3455 -1593 3655 -1577
rect 3961 -1543 4161 -1505
rect 3961 -1577 4010 -1543
rect 4044 -1577 4078 -1543
rect 4112 -1577 4161 -1543
rect 3961 -1593 4161 -1577
rect 4219 -1543 4419 -1505
rect 4219 -1577 4268 -1543
rect 4302 -1577 4336 -1543
rect 4370 -1577 4419 -1543
rect 4219 -1593 4419 -1577
rect 4724 -1543 4924 -1505
rect 4724 -1577 4773 -1543
rect 4807 -1577 4841 -1543
rect 4875 -1577 4924 -1543
rect 4724 -1593 4924 -1577
rect 4982 -1543 5182 -1505
rect 4982 -1577 5031 -1543
rect 5065 -1577 5099 -1543
rect 5133 -1577 5182 -1543
rect 4982 -1593 5182 -1577
rect 5240 -1543 5440 -1505
rect 5240 -1577 5289 -1543
rect 5323 -1577 5357 -1543
rect 5391 -1577 5440 -1543
rect 5240 -1593 5440 -1577
rect 5745 -1543 5945 -1505
rect 5745 -1577 5794 -1543
rect 5828 -1577 5862 -1543
rect 5896 -1577 5945 -1543
rect 5745 -1593 5945 -1577
rect 6003 -1543 6203 -1505
rect 6003 -1577 6052 -1543
rect 6086 -1577 6120 -1543
rect 6154 -1577 6203 -1543
rect 6003 -1593 6203 -1577
rect 6508 -1543 6708 -1505
rect 6508 -1577 6557 -1543
rect 6591 -1577 6625 -1543
rect 6659 -1577 6708 -1543
rect 6508 -1593 6708 -1577
rect -84 -1906 116 -1890
rect -84 -1940 -35 -1906
rect -1 -1940 33 -1906
rect 67 -1940 116 -1906
rect -84 -1978 116 -1940
rect 421 -1906 621 -1890
rect 421 -1940 470 -1906
rect 504 -1940 538 -1906
rect 572 -1940 621 -1906
rect 421 -1978 621 -1940
rect 679 -1906 879 -1890
rect 679 -1940 728 -1906
rect 762 -1940 796 -1906
rect 830 -1940 879 -1906
rect 679 -1978 879 -1940
rect 1184 -1906 1384 -1890
rect 1184 -1940 1233 -1906
rect 1267 -1940 1301 -1906
rect 1335 -1940 1384 -1906
rect 1184 -1978 1384 -1940
rect 1442 -1906 1642 -1890
rect 1442 -1940 1491 -1906
rect 1525 -1940 1559 -1906
rect 1593 -1940 1642 -1906
rect 1442 -1978 1642 -1940
rect 1700 -1906 1900 -1890
rect 1700 -1940 1749 -1906
rect 1783 -1940 1817 -1906
rect 1851 -1940 1900 -1906
rect 1700 -1978 1900 -1940
rect 2205 -1906 2405 -1890
rect 2205 -1940 2254 -1906
rect 2288 -1940 2322 -1906
rect 2356 -1940 2405 -1906
rect 2205 -1978 2405 -1940
rect 2463 -1906 2663 -1890
rect 2463 -1940 2512 -1906
rect 2546 -1940 2580 -1906
rect 2614 -1940 2663 -1906
rect 2463 -1978 2663 -1940
rect 2969 -1906 3169 -1890
rect 2969 -1940 3018 -1906
rect 3052 -1940 3086 -1906
rect 3120 -1940 3169 -1906
rect 2969 -1978 3169 -1940
rect 3455 -1906 3655 -1890
rect 3455 -1940 3504 -1906
rect 3538 -1940 3572 -1906
rect 3606 -1940 3655 -1906
rect 3455 -1978 3655 -1940
rect 3961 -1906 4161 -1890
rect 3961 -1940 4010 -1906
rect 4044 -1940 4078 -1906
rect 4112 -1940 4161 -1906
rect 3961 -1978 4161 -1940
rect 4219 -1906 4419 -1890
rect 4219 -1940 4268 -1906
rect 4302 -1940 4336 -1906
rect 4370 -1940 4419 -1906
rect 4219 -1978 4419 -1940
rect 4724 -1906 4924 -1890
rect 4724 -1940 4773 -1906
rect 4807 -1940 4841 -1906
rect 4875 -1940 4924 -1906
rect 4724 -1978 4924 -1940
rect 4982 -1906 5182 -1890
rect 4982 -1940 5031 -1906
rect 5065 -1940 5099 -1906
rect 5133 -1940 5182 -1906
rect 4982 -1978 5182 -1940
rect 5240 -1906 5440 -1890
rect 5240 -1940 5289 -1906
rect 5323 -1940 5357 -1906
rect 5391 -1940 5440 -1906
rect 5240 -1978 5440 -1940
rect 5745 -1906 5945 -1890
rect 5745 -1940 5794 -1906
rect 5828 -1940 5862 -1906
rect 5896 -1940 5945 -1906
rect 5745 -1978 5945 -1940
rect 6003 -1906 6203 -1890
rect 6003 -1940 6052 -1906
rect 6086 -1940 6120 -1906
rect 6154 -1940 6203 -1906
rect 6003 -1978 6203 -1940
rect 6508 -1906 6708 -1890
rect 6508 -1940 6557 -1906
rect 6591 -1940 6625 -1906
rect 6659 -1940 6708 -1906
rect 6508 -1978 6708 -1940
rect -84 -2204 116 -2178
rect 421 -2204 621 -2178
rect 679 -2204 879 -2178
rect 1184 -2204 1384 -2178
rect 1442 -2204 1642 -2178
rect 1700 -2204 1900 -2178
rect 2205 -2204 2405 -2178
rect 2463 -2204 2663 -2178
rect 2969 -2204 3169 -2178
rect 3455 -2204 3655 -2178
rect 3961 -2204 4161 -2178
rect 4219 -2204 4419 -2178
rect 4724 -2204 4924 -2178
rect 4982 -2204 5182 -2178
rect 5240 -2204 5440 -2178
rect 5745 -2204 5945 -2178
rect 6003 -2204 6203 -2178
rect 6508 -2204 6708 -2178
rect -84 -2704 116 -2678
rect 421 -2704 621 -2678
rect 679 -2704 879 -2678
rect 1184 -2704 1384 -2678
rect 1442 -2704 1642 -2678
rect 1700 -2704 1900 -2678
rect 2205 -2704 2405 -2678
rect 2463 -2704 2663 -2678
rect 2969 -2704 3169 -2678
rect 3455 -2704 3655 -2678
rect 3961 -2704 4161 -2678
rect 4219 -2704 4419 -2678
rect 4724 -2704 4924 -2678
rect 4982 -2704 5182 -2678
rect 5240 -2704 5440 -2678
rect 5745 -2704 5945 -2678
rect 6003 -2704 6203 -2678
rect 6508 -2704 6708 -2678
rect -84 -2942 116 -2904
rect -84 -2976 -35 -2942
rect -1 -2976 33 -2942
rect 67 -2976 116 -2942
rect -84 -2992 116 -2976
rect 421 -2942 621 -2904
rect 421 -2976 470 -2942
rect 504 -2976 538 -2942
rect 572 -2976 621 -2942
rect 421 -2992 621 -2976
rect 679 -2942 879 -2904
rect 679 -2976 728 -2942
rect 762 -2976 796 -2942
rect 830 -2976 879 -2942
rect 679 -2992 879 -2976
rect 1184 -2942 1384 -2904
rect 1184 -2976 1233 -2942
rect 1267 -2976 1301 -2942
rect 1335 -2976 1384 -2942
rect 1184 -2992 1384 -2976
rect 1442 -2942 1642 -2904
rect 1442 -2976 1491 -2942
rect 1525 -2976 1559 -2942
rect 1593 -2976 1642 -2942
rect 1442 -2992 1642 -2976
rect 1700 -2942 1900 -2904
rect 1700 -2976 1749 -2942
rect 1783 -2976 1817 -2942
rect 1851 -2976 1900 -2942
rect 1700 -2992 1900 -2976
rect 2205 -2942 2405 -2904
rect 2205 -2976 2254 -2942
rect 2288 -2976 2322 -2942
rect 2356 -2976 2405 -2942
rect 2205 -2992 2405 -2976
rect 2463 -2942 2663 -2904
rect 2463 -2976 2512 -2942
rect 2546 -2976 2580 -2942
rect 2614 -2976 2663 -2942
rect 2463 -2992 2663 -2976
rect 2969 -2942 3169 -2904
rect 2969 -2976 3018 -2942
rect 3052 -2976 3086 -2942
rect 3120 -2976 3169 -2942
rect 2969 -2992 3169 -2976
rect 3455 -2942 3655 -2904
rect 3455 -2976 3504 -2942
rect 3538 -2976 3572 -2942
rect 3606 -2976 3655 -2942
rect 3455 -2992 3655 -2976
rect 3961 -2942 4161 -2904
rect 3961 -2976 4010 -2942
rect 4044 -2976 4078 -2942
rect 4112 -2976 4161 -2942
rect 3961 -2992 4161 -2976
rect 4219 -2942 4419 -2904
rect 4219 -2976 4268 -2942
rect 4302 -2976 4336 -2942
rect 4370 -2976 4419 -2942
rect 4219 -2992 4419 -2976
rect 4724 -2942 4924 -2904
rect 4724 -2976 4773 -2942
rect 4807 -2976 4841 -2942
rect 4875 -2976 4924 -2942
rect 4724 -2992 4924 -2976
rect 4982 -2942 5182 -2904
rect 4982 -2976 5031 -2942
rect 5065 -2976 5099 -2942
rect 5133 -2976 5182 -2942
rect 4982 -2992 5182 -2976
rect 5240 -2942 5440 -2904
rect 5240 -2976 5289 -2942
rect 5323 -2976 5357 -2942
rect 5391 -2976 5440 -2942
rect 5240 -2992 5440 -2976
rect 5745 -2942 5945 -2904
rect 5745 -2976 5794 -2942
rect 5828 -2976 5862 -2942
rect 5896 -2976 5945 -2942
rect 5745 -2992 5945 -2976
rect 6003 -2942 6203 -2904
rect 6003 -2976 6052 -2942
rect 6086 -2976 6120 -2942
rect 6154 -2976 6203 -2942
rect 6003 -2992 6203 -2976
rect 6508 -2942 6708 -2904
rect 6508 -2976 6557 -2942
rect 6591 -2976 6625 -2942
rect 6659 -2976 6708 -2942
rect 6508 -2992 6708 -2976
<< polycont >>
rect -35 856 -1 890
rect 33 856 67 890
rect 470 856 504 890
rect 538 856 572 890
rect 728 856 762 890
rect 796 856 830 890
rect 1233 856 1267 890
rect 1301 856 1335 890
rect 1491 856 1525 890
rect 1559 856 1593 890
rect 1749 856 1783 890
rect 1817 856 1851 890
rect 2254 856 2288 890
rect 2322 856 2356 890
rect 2512 856 2546 890
rect 2580 856 2614 890
rect 3018 856 3052 890
rect 3086 856 3120 890
rect 3504 856 3538 890
rect 3572 856 3606 890
rect 4010 856 4044 890
rect 4078 856 4112 890
rect 4268 856 4302 890
rect 4336 856 4370 890
rect 4773 856 4807 890
rect 4841 856 4875 890
rect 5031 856 5065 890
rect 5099 856 5133 890
rect 5289 856 5323 890
rect 5357 856 5391 890
rect 5794 856 5828 890
rect 5862 856 5896 890
rect 6052 856 6086 890
rect 6120 856 6154 890
rect 6557 856 6591 890
rect 6625 856 6659 890
rect -35 -180 -1 -146
rect 33 -180 67 -146
rect 470 -180 504 -146
rect 538 -180 572 -146
rect 728 -180 762 -146
rect 796 -180 830 -146
rect 1233 -180 1267 -146
rect 1301 -180 1335 -146
rect 1491 -180 1525 -146
rect 1559 -180 1593 -146
rect 1749 -180 1783 -146
rect 1817 -180 1851 -146
rect 2254 -180 2288 -146
rect 2322 -180 2356 -146
rect 2512 -180 2546 -146
rect 2580 -180 2614 -146
rect 3018 -180 3052 -146
rect 3086 -180 3120 -146
rect 3504 -180 3538 -146
rect 3572 -180 3606 -146
rect 4010 -180 4044 -146
rect 4078 -180 4112 -146
rect 4268 -180 4302 -146
rect 4336 -180 4370 -146
rect 4773 -180 4807 -146
rect 4841 -180 4875 -146
rect 5031 -180 5065 -146
rect 5099 -180 5133 -146
rect 5289 -180 5323 -146
rect 5357 -180 5391 -146
rect 5794 -180 5828 -146
rect 5862 -180 5896 -146
rect 6052 -180 6086 -146
rect 6120 -180 6154 -146
rect 6557 -180 6591 -146
rect 6625 -180 6659 -146
rect -35 -543 -1 -509
rect 33 -543 67 -509
rect 470 -543 504 -509
rect 538 -543 572 -509
rect 728 -543 762 -509
rect 796 -543 830 -509
rect 1233 -543 1267 -509
rect 1301 -543 1335 -509
rect 1491 -543 1525 -509
rect 1559 -543 1593 -509
rect 1749 -543 1783 -509
rect 1817 -543 1851 -509
rect 2254 -543 2288 -509
rect 2322 -543 2356 -509
rect 2512 -543 2546 -509
rect 2580 -543 2614 -509
rect 3018 -543 3052 -509
rect 3086 -543 3120 -509
rect 3504 -543 3538 -509
rect 3572 -543 3606 -509
rect 4010 -543 4044 -509
rect 4078 -543 4112 -509
rect 4268 -543 4302 -509
rect 4336 -543 4370 -509
rect 4773 -543 4807 -509
rect 4841 -543 4875 -509
rect 5031 -543 5065 -509
rect 5099 -543 5133 -509
rect 5289 -543 5323 -509
rect 5357 -543 5391 -509
rect 5794 -543 5828 -509
rect 5862 -543 5896 -509
rect 6052 -543 6086 -509
rect 6120 -543 6154 -509
rect 6557 -543 6591 -509
rect 6625 -543 6659 -509
rect -35 -1577 -1 -1543
rect 33 -1577 67 -1543
rect 470 -1577 504 -1543
rect 538 -1577 572 -1543
rect 728 -1577 762 -1543
rect 796 -1577 830 -1543
rect 1233 -1577 1267 -1543
rect 1301 -1577 1335 -1543
rect 1491 -1577 1525 -1543
rect 1559 -1577 1593 -1543
rect 1749 -1577 1783 -1543
rect 1817 -1577 1851 -1543
rect 2254 -1577 2288 -1543
rect 2322 -1577 2356 -1543
rect 2512 -1577 2546 -1543
rect 2580 -1577 2614 -1543
rect 3018 -1577 3052 -1543
rect 3086 -1577 3120 -1543
rect 3504 -1577 3538 -1543
rect 3572 -1577 3606 -1543
rect 4010 -1577 4044 -1543
rect 4078 -1577 4112 -1543
rect 4268 -1577 4302 -1543
rect 4336 -1577 4370 -1543
rect 4773 -1577 4807 -1543
rect 4841 -1577 4875 -1543
rect 5031 -1577 5065 -1543
rect 5099 -1577 5133 -1543
rect 5289 -1577 5323 -1543
rect 5357 -1577 5391 -1543
rect 5794 -1577 5828 -1543
rect 5862 -1577 5896 -1543
rect 6052 -1577 6086 -1543
rect 6120 -1577 6154 -1543
rect 6557 -1577 6591 -1543
rect 6625 -1577 6659 -1543
rect -35 -1940 -1 -1906
rect 33 -1940 67 -1906
rect 470 -1940 504 -1906
rect 538 -1940 572 -1906
rect 728 -1940 762 -1906
rect 796 -1940 830 -1906
rect 1233 -1940 1267 -1906
rect 1301 -1940 1335 -1906
rect 1491 -1940 1525 -1906
rect 1559 -1940 1593 -1906
rect 1749 -1940 1783 -1906
rect 1817 -1940 1851 -1906
rect 2254 -1940 2288 -1906
rect 2322 -1940 2356 -1906
rect 2512 -1940 2546 -1906
rect 2580 -1940 2614 -1906
rect 3018 -1940 3052 -1906
rect 3086 -1940 3120 -1906
rect 3504 -1940 3538 -1906
rect 3572 -1940 3606 -1906
rect 4010 -1940 4044 -1906
rect 4078 -1940 4112 -1906
rect 4268 -1940 4302 -1906
rect 4336 -1940 4370 -1906
rect 4773 -1940 4807 -1906
rect 4841 -1940 4875 -1906
rect 5031 -1940 5065 -1906
rect 5099 -1940 5133 -1906
rect 5289 -1940 5323 -1906
rect 5357 -1940 5391 -1906
rect 5794 -1940 5828 -1906
rect 5862 -1940 5896 -1906
rect 6052 -1940 6086 -1906
rect 6120 -1940 6154 -1906
rect 6557 -1940 6591 -1906
rect 6625 -1940 6659 -1906
rect -35 -2976 -1 -2942
rect 33 -2976 67 -2942
rect 470 -2976 504 -2942
rect 538 -2976 572 -2942
rect 728 -2976 762 -2942
rect 796 -2976 830 -2942
rect 1233 -2976 1267 -2942
rect 1301 -2976 1335 -2942
rect 1491 -2976 1525 -2942
rect 1559 -2976 1593 -2942
rect 1749 -2976 1783 -2942
rect 1817 -2976 1851 -2942
rect 2254 -2976 2288 -2942
rect 2322 -2976 2356 -2942
rect 2512 -2976 2546 -2942
rect 2580 -2976 2614 -2942
rect 3018 -2976 3052 -2942
rect 3086 -2976 3120 -2942
rect 3504 -2976 3538 -2942
rect 3572 -2976 3606 -2942
rect 4010 -2976 4044 -2942
rect 4078 -2976 4112 -2942
rect 4268 -2976 4302 -2942
rect 4336 -2976 4370 -2942
rect 4773 -2976 4807 -2942
rect 4841 -2976 4875 -2942
rect 5031 -2976 5065 -2942
rect 5099 -2976 5133 -2942
rect 5289 -2976 5323 -2942
rect 5357 -2976 5391 -2942
rect 5794 -2976 5828 -2942
rect 5862 -2976 5896 -2942
rect 6052 -2976 6086 -2942
rect 6120 -2976 6154 -2942
rect 6557 -2976 6591 -2942
rect 6625 -2976 6659 -2942
<< locali >>
rect -244 955 -80 989
rect -25 955 -8 989
rect 43 955 64 989
rect 111 955 136 989
rect 179 955 208 989
rect 247 955 280 989
rect 315 955 349 989
rect 386 955 417 989
rect 458 955 485 989
rect 530 955 553 989
rect 602 955 621 989
rect 674 955 689 989
rect 746 955 757 989
rect 818 955 825 989
rect 890 955 893 989
rect 927 955 928 989
rect 995 955 1000 989
rect 1063 955 1072 989
rect 1131 955 1144 989
rect 1199 955 1216 989
rect 1267 955 1288 989
rect 1335 955 1360 989
rect 1403 955 1432 989
rect 1471 955 1504 989
rect 1539 955 1573 989
rect 1610 955 1641 989
rect 1682 955 1709 989
rect 1754 955 1777 989
rect 1826 955 1845 989
rect 1898 955 1913 989
rect 1970 955 1981 989
rect 2042 955 2049 989
rect 2114 955 2117 989
rect 2151 955 2152 989
rect 2219 955 2224 989
rect 2287 955 2296 989
rect 2355 955 2368 989
rect 2423 955 2440 989
rect 2491 955 2512 989
rect 2559 955 2584 989
rect 2627 955 2656 989
rect 2695 955 2728 989
rect 2763 955 2797 989
rect 2834 955 2865 989
rect 2906 955 2933 989
rect 2978 955 3001 989
rect 3050 955 3069 989
rect 3122 955 3137 989
rect 3194 955 3430 989
rect 3487 955 3502 989
rect 3555 955 3574 989
rect 3623 955 3646 989
rect 3691 955 3718 989
rect 3759 955 3790 989
rect 3827 955 3861 989
rect 3896 955 3929 989
rect 3968 955 3997 989
rect 4040 955 4065 989
rect 4112 955 4133 989
rect 4184 955 4201 989
rect 4256 955 4269 989
rect 4328 955 4337 989
rect 4400 955 4405 989
rect 4472 955 4473 989
rect 4507 955 4510 989
rect 4575 955 4582 989
rect 4643 955 4654 989
rect 4711 955 4726 989
rect 4779 955 4798 989
rect 4847 955 4870 989
rect 4915 955 4942 989
rect 4983 955 5014 989
rect 5051 955 5085 989
rect 5120 955 5153 989
rect 5192 955 5221 989
rect 5264 955 5289 989
rect 5336 955 5357 989
rect 5408 955 5425 989
rect 5480 955 5493 989
rect 5552 955 5561 989
rect 5624 955 5629 989
rect 5696 955 5697 989
rect 5731 955 5734 989
rect 5799 955 5806 989
rect 5867 955 5878 989
rect 5935 955 5950 989
rect 6003 955 6022 989
rect 6071 955 6094 989
rect 6139 955 6166 989
rect 6207 955 6238 989
rect 6275 955 6309 989
rect 6344 955 6377 989
rect 6416 955 6445 989
rect 6488 955 6513 989
rect 6560 955 6581 989
rect 6632 955 6649 989
rect 6704 955 6868 989
rect -244 882 -210 955
rect -84 856 -37 890
rect -1 856 33 890
rect 69 856 116 890
rect 421 856 468 890
rect 504 856 538 890
rect 574 856 621 890
rect 679 856 726 890
rect 762 856 796 890
rect 832 856 879 890
rect 1184 856 1231 890
rect 1267 856 1301 890
rect 1337 856 1384 890
rect 1442 856 1489 890
rect 1525 856 1559 890
rect 1595 856 1642 890
rect 1700 856 1747 890
rect 1783 856 1817 890
rect 1853 856 1900 890
rect 2205 856 2252 890
rect 2288 856 2322 890
rect 2358 856 2405 890
rect 2463 856 2510 890
rect 2546 856 2580 890
rect 2616 856 2663 890
rect 2969 856 3016 890
rect 3052 856 3086 890
rect 3122 856 3169 890
rect 3295 882 3329 955
rect 3455 856 3502 890
rect 3538 856 3572 890
rect 3608 856 3655 890
rect 3961 856 4008 890
rect 4044 856 4078 890
rect 4114 856 4161 890
rect 4219 856 4266 890
rect 4302 856 4336 890
rect 4372 856 4419 890
rect 4724 856 4771 890
rect 4807 856 4841 890
rect 4877 856 4924 890
rect 4982 856 5029 890
rect 5065 856 5099 890
rect 5135 856 5182 890
rect 5240 856 5287 890
rect 5323 856 5357 890
rect 5393 856 5440 890
rect 5745 856 5792 890
rect 5828 856 5862 890
rect 5898 856 5945 890
rect 6003 856 6050 890
rect 6086 856 6120 890
rect 6156 856 6203 890
rect 6508 856 6555 890
rect 6591 856 6625 890
rect 6661 856 6708 890
rect 6834 882 6868 955
rect -244 810 -210 814
rect -244 738 -210 746
rect -244 666 -210 678
rect -130 803 -96 822
rect -130 735 -96 737
rect -130 699 -96 701
rect -130 614 -96 633
rect 128 803 162 822
rect 128 735 162 737
rect 128 699 162 701
rect 128 614 162 633
rect 375 803 409 822
rect 375 735 409 737
rect 375 699 409 701
rect 375 614 409 633
rect 633 803 667 822
rect 633 735 667 737
rect 633 699 667 701
rect 633 614 667 633
rect 891 803 925 822
rect 891 735 925 737
rect 891 699 925 701
rect 891 614 925 633
rect 1138 803 1172 822
rect 1138 735 1172 737
rect 1138 699 1172 701
rect 1138 614 1172 633
rect 1396 803 1430 822
rect 1396 735 1430 737
rect 1396 699 1430 701
rect 1396 614 1430 633
rect 1654 803 1688 822
rect 1654 735 1688 737
rect 1654 699 1688 701
rect 1654 614 1688 633
rect 1912 803 1946 822
rect 1912 735 1946 737
rect 1912 699 1946 701
rect 1912 614 1946 633
rect 2159 803 2193 822
rect 2159 735 2193 737
rect 2159 699 2193 701
rect 2159 614 2193 633
rect 2417 803 2451 822
rect 2417 735 2451 737
rect 2417 699 2451 701
rect 2417 614 2451 633
rect 2675 803 2709 822
rect 2675 735 2709 737
rect 2675 699 2709 701
rect 2675 614 2709 633
rect 2923 803 2957 822
rect 2923 735 2957 737
rect 2923 699 2957 701
rect 2923 614 2957 633
rect 3181 803 3215 822
rect 3181 735 3215 737
rect 3181 699 3215 701
rect 3181 614 3215 633
rect 3295 810 3329 814
rect 3295 738 3329 746
rect 3295 666 3329 678
rect -244 594 -210 610
rect -244 522 -210 542
rect -244 450 -210 474
rect -244 378 -210 406
rect 3409 803 3443 822
rect 3409 735 3443 737
rect 3409 699 3443 701
rect 3409 614 3443 633
rect 3667 803 3701 822
rect 3667 735 3701 737
rect 3667 699 3701 701
rect 3667 614 3701 633
rect 3915 803 3949 822
rect 3915 735 3949 737
rect 3915 699 3949 701
rect 3915 614 3949 633
rect 4173 803 4207 822
rect 4173 735 4207 737
rect 4173 699 4207 701
rect 4173 614 4207 633
rect 4431 803 4465 822
rect 4431 735 4465 737
rect 4431 699 4465 701
rect 4431 614 4465 633
rect 4678 803 4712 822
rect 4678 735 4712 737
rect 4678 699 4712 701
rect 4678 614 4712 633
rect 4936 803 4970 822
rect 4936 735 4970 737
rect 4936 699 4970 701
rect 4936 614 4970 633
rect 5194 803 5228 822
rect 5194 735 5228 737
rect 5194 699 5228 701
rect 5194 614 5228 633
rect 5452 803 5486 822
rect 5452 735 5486 737
rect 5452 699 5486 701
rect 5452 614 5486 633
rect 5699 803 5733 822
rect 5699 735 5733 737
rect 5699 699 5733 701
rect 5699 614 5733 633
rect 5957 803 5991 822
rect 5957 735 5991 737
rect 5957 699 5991 701
rect 5957 614 5991 633
rect 6215 803 6249 822
rect 6215 735 6249 737
rect 6215 699 6249 701
rect 6215 614 6249 633
rect 6462 803 6496 822
rect 6462 735 6496 737
rect 6462 699 6496 701
rect 6462 614 6496 633
rect 6720 803 6754 822
rect 6720 735 6754 737
rect 6720 699 6754 701
rect 6720 614 6754 633
rect 6834 810 6868 814
rect 6834 738 6868 746
rect 6834 666 6868 678
rect 3295 594 3329 610
rect 3295 522 3329 542
rect 3295 450 3329 474
rect 3295 378 3329 406
rect 6834 594 6868 610
rect 6834 522 6868 542
rect 6834 450 6868 474
rect 6834 378 6868 406
rect -210 338 -59 372
rect -25 338 9 372
rect 43 338 77 372
rect 111 338 145 372
rect 179 338 213 372
rect 247 338 281 372
rect 315 338 349 372
rect 383 338 417 372
rect 451 338 485 372
rect 519 338 553 372
rect 587 338 621 372
rect 655 338 689 372
rect 723 338 757 372
rect 791 338 825 372
rect 859 338 893 372
rect 927 338 961 372
rect 995 338 1029 372
rect 1063 338 1097 372
rect 1131 338 1165 372
rect 1199 338 1233 372
rect 1267 338 1301 372
rect 1335 338 1369 372
rect 1403 338 1437 372
rect 1471 338 1505 372
rect 1539 338 1573 372
rect 1607 338 1641 372
rect 1675 338 1709 372
rect 1743 338 1777 372
rect 1811 338 1845 372
rect 1879 338 1913 372
rect 1947 338 1981 372
rect 2015 338 2049 372
rect 2083 338 2117 372
rect 2151 338 2185 372
rect 2219 338 2253 372
rect 2287 338 2321 372
rect 2355 338 2389 372
rect 2423 338 2457 372
rect 2491 338 2525 372
rect 2559 338 2593 372
rect 2627 338 2661 372
rect 2695 338 2729 372
rect 2763 338 2797 372
rect 2831 338 2865 372
rect 2899 338 2933 372
rect 2967 338 3001 372
rect 3035 338 3069 372
rect 3103 338 3137 372
rect 3171 338 3295 372
rect 3329 338 3453 372
rect 3487 338 3521 372
rect 3555 338 3589 372
rect 3623 338 3657 372
rect 3691 338 3725 372
rect 3759 338 3793 372
rect 3827 338 3861 372
rect 3895 338 3929 372
rect 3963 338 3997 372
rect 4031 338 4065 372
rect 4099 338 4133 372
rect 4167 338 4201 372
rect 4235 338 4269 372
rect 4303 338 4337 372
rect 4371 338 4405 372
rect 4439 338 4473 372
rect 4507 338 4541 372
rect 4575 338 4609 372
rect 4643 338 4677 372
rect 4711 338 4745 372
rect 4779 338 4813 372
rect 4847 338 4881 372
rect 4915 338 4949 372
rect 4983 338 5017 372
rect 5051 338 5085 372
rect 5119 338 5153 372
rect 5187 338 5221 372
rect 5255 338 5289 372
rect 5323 338 5357 372
rect 5391 338 5425 372
rect 5459 338 5493 372
rect 5527 338 5561 372
rect 5595 338 5629 372
rect 5663 338 5697 372
rect 5731 338 5765 372
rect 5799 338 5833 372
rect 5867 338 5901 372
rect 5935 338 5969 372
rect 6003 338 6037 372
rect 6071 338 6105 372
rect 6139 338 6173 372
rect 6207 338 6241 372
rect 6275 338 6309 372
rect 6343 338 6377 372
rect 6411 338 6445 372
rect 6479 338 6513 372
rect 6547 338 6581 372
rect 6615 338 6649 372
rect 6683 338 6834 372
rect -244 306 -210 338
rect -244 236 -210 270
rect -244 168 -210 200
rect -244 100 -210 128
rect 3295 306 3329 338
rect 3295 236 3329 270
rect 3295 168 3329 200
rect 3295 100 3329 128
rect -244 32 -210 56
rect -244 -36 -210 -16
rect -244 -104 -210 -88
rect -130 77 -96 96
rect -130 9 -96 11
rect -130 -27 -96 -25
rect -130 -112 -96 -93
rect 128 77 162 96
rect 128 9 162 11
rect 128 -27 162 -25
rect 128 -112 162 -93
rect 375 77 409 96
rect 375 9 409 11
rect 375 -27 409 -25
rect 375 -112 409 -93
rect 633 77 667 96
rect 633 9 667 11
rect 633 -27 667 -25
rect 633 -112 667 -93
rect 891 77 925 96
rect 891 9 925 11
rect 891 -27 925 -25
rect 891 -112 925 -93
rect 1138 77 1172 96
rect 1138 9 1172 11
rect 1138 -27 1172 -25
rect 1138 -112 1172 -93
rect 1396 77 1430 96
rect 1396 9 1430 11
rect 1396 -27 1430 -25
rect 1396 -112 1430 -93
rect 1654 77 1688 96
rect 1654 9 1688 11
rect 1654 -27 1688 -25
rect 1654 -112 1688 -93
rect 1912 77 1946 96
rect 1912 9 1946 11
rect 1912 -27 1946 -25
rect 1912 -112 1946 -93
rect 2159 77 2193 96
rect 2159 9 2193 11
rect 2159 -27 2193 -25
rect 2159 -112 2193 -93
rect 2417 77 2451 96
rect 2417 9 2451 11
rect 2417 -27 2451 -25
rect 2417 -112 2451 -93
rect 2675 77 2709 96
rect 2675 9 2709 11
rect 2675 -27 2709 -25
rect 2675 -112 2709 -93
rect 2923 77 2957 96
rect 2923 9 2957 11
rect 2923 -27 2957 -25
rect 2923 -112 2957 -93
rect 3181 77 3215 96
rect 3181 9 3215 11
rect 3181 -27 3215 -25
rect 3181 -112 3215 -93
rect 6834 306 6868 338
rect 6834 236 6868 270
rect 6834 168 6868 200
rect 6834 100 6868 128
rect 3295 32 3329 56
rect 3295 -36 3329 -16
rect 3295 -104 3329 -88
rect 3409 77 3443 96
rect 3409 9 3443 11
rect 3409 -27 3443 -25
rect 3409 -112 3443 -93
rect 3667 77 3701 96
rect 3667 9 3701 11
rect 3667 -27 3701 -25
rect 3667 -112 3701 -93
rect 3915 77 3949 96
rect 3915 9 3949 11
rect 3915 -27 3949 -25
rect 3915 -112 3949 -93
rect 4173 77 4207 96
rect 4173 9 4207 11
rect 4173 -27 4207 -25
rect 4173 -112 4207 -93
rect 4431 77 4465 96
rect 4431 9 4465 11
rect 4431 -27 4465 -25
rect 4431 -112 4465 -93
rect 4678 77 4712 96
rect 4678 9 4712 11
rect 4678 -27 4712 -25
rect 4678 -112 4712 -93
rect 4936 77 4970 96
rect 4936 9 4970 11
rect 4936 -27 4970 -25
rect 4936 -112 4970 -93
rect 5194 77 5228 96
rect 5194 9 5228 11
rect 5194 -27 5228 -25
rect 5194 -112 5228 -93
rect 5452 77 5486 96
rect 5452 9 5486 11
rect 5452 -27 5486 -25
rect 5452 -112 5486 -93
rect 5699 77 5733 96
rect 5699 9 5733 11
rect 5699 -27 5733 -25
rect 5699 -112 5733 -93
rect 5957 77 5991 96
rect 5957 9 5991 11
rect 5957 -27 5991 -25
rect 5957 -112 5991 -93
rect 6215 77 6249 96
rect 6215 9 6249 11
rect 6215 -27 6249 -25
rect 6215 -112 6249 -93
rect 6462 77 6496 96
rect 6462 9 6496 11
rect 6462 -27 6496 -25
rect 6462 -112 6496 -93
rect 6720 77 6754 96
rect 6720 9 6754 11
rect 6720 -27 6754 -25
rect 6720 -112 6754 -93
rect 6834 32 6868 56
rect 6834 -36 6868 -16
rect 6834 -104 6868 -88
rect -244 -172 -210 -160
rect -84 -180 -37 -146
rect -1 -180 33 -146
rect 69 -180 116 -146
rect 421 -180 468 -146
rect 504 -180 538 -146
rect 574 -180 621 -146
rect 679 -180 726 -146
rect 762 -180 796 -146
rect 832 -180 879 -146
rect 1184 -180 1231 -146
rect 1267 -180 1301 -146
rect 1337 -180 1384 -146
rect 1442 -180 1489 -146
rect 1525 -180 1559 -146
rect 1595 -180 1642 -146
rect 1700 -180 1747 -146
rect 1783 -180 1817 -146
rect 1853 -180 1900 -146
rect 2205 -180 2252 -146
rect 2288 -180 2322 -146
rect 2358 -180 2405 -146
rect 2463 -180 2510 -146
rect 2546 -180 2580 -146
rect 2616 -180 2663 -146
rect 2969 -180 3016 -146
rect 3052 -180 3086 -146
rect 3122 -180 3169 -146
rect 3295 -172 3329 -160
rect -244 -240 -210 -232
rect -244 -308 -210 -304
rect -244 -414 -210 -410
rect -244 -486 -210 -478
rect 3455 -180 3502 -146
rect 3538 -180 3572 -146
rect 3608 -180 3655 -146
rect 3961 -180 4008 -146
rect 4044 -180 4078 -146
rect 4114 -180 4161 -146
rect 4219 -180 4266 -146
rect 4302 -180 4336 -146
rect 4372 -180 4419 -146
rect 4724 -180 4771 -146
rect 4807 -180 4841 -146
rect 4877 -180 4924 -146
rect 4982 -180 5029 -146
rect 5065 -180 5099 -146
rect 5135 -180 5182 -146
rect 5240 -180 5287 -146
rect 5323 -180 5357 -146
rect 5393 -180 5440 -146
rect 5745 -180 5792 -146
rect 5828 -180 5862 -146
rect 5898 -180 5945 -146
rect 6003 -180 6050 -146
rect 6086 -180 6120 -146
rect 6156 -180 6203 -146
rect 6508 -180 6555 -146
rect 6591 -180 6625 -146
rect 6661 -180 6708 -146
rect 6834 -172 6868 -160
rect 3295 -240 3329 -232
rect 3295 -308 3329 -304
rect 3295 -414 3329 -410
rect 3295 -486 3329 -478
rect -84 -543 -37 -509
rect -1 -543 33 -509
rect 69 -543 116 -509
rect 421 -543 468 -509
rect 504 -543 538 -509
rect 574 -543 621 -509
rect 679 -543 726 -509
rect 762 -543 796 -509
rect 832 -543 879 -509
rect 1184 -543 1231 -509
rect 1267 -543 1301 -509
rect 1337 -543 1384 -509
rect 1442 -543 1489 -509
rect 1525 -543 1559 -509
rect 1595 -543 1642 -509
rect 1700 -543 1747 -509
rect 1783 -543 1817 -509
rect 1853 -543 1900 -509
rect 2205 -543 2252 -509
rect 2288 -543 2322 -509
rect 2358 -543 2405 -509
rect 2463 -543 2510 -509
rect 2546 -543 2580 -509
rect 2616 -543 2663 -509
rect 2969 -543 3016 -509
rect 3052 -543 3086 -509
rect 3122 -543 3169 -509
rect 6834 -240 6868 -232
rect 6834 -308 6868 -304
rect 6834 -414 6868 -410
rect 6834 -486 6868 -478
rect -244 -558 -210 -546
rect 3455 -543 3502 -509
rect 3538 -543 3572 -509
rect 3608 -543 3655 -509
rect 3961 -543 4008 -509
rect 4044 -543 4078 -509
rect 4114 -543 4161 -509
rect 4219 -543 4266 -509
rect 4302 -543 4336 -509
rect 4372 -543 4419 -509
rect 4724 -543 4771 -509
rect 4807 -543 4841 -509
rect 4877 -543 4924 -509
rect 4982 -543 5029 -509
rect 5065 -543 5099 -509
rect 5135 -543 5182 -509
rect 5240 -543 5287 -509
rect 5323 -543 5357 -509
rect 5393 -543 5440 -509
rect 5745 -543 5792 -509
rect 5828 -543 5862 -509
rect 5898 -543 5945 -509
rect 6003 -543 6050 -509
rect 6086 -543 6120 -509
rect 6156 -543 6203 -509
rect 6508 -543 6555 -509
rect 6591 -543 6625 -509
rect 6661 -543 6708 -509
rect 3295 -558 3329 -546
rect -244 -630 -210 -614
rect -244 -702 -210 -682
rect -244 -774 -210 -750
rect -130 -596 -96 -577
rect -130 -664 -96 -662
rect -130 -700 -96 -698
rect -130 -785 -96 -766
rect 128 -596 162 -577
rect 128 -664 162 -662
rect 128 -700 162 -698
rect 128 -785 162 -766
rect 375 -596 409 -577
rect 375 -664 409 -662
rect 375 -700 409 -698
rect 375 -785 409 -766
rect 633 -596 667 -577
rect 633 -664 667 -662
rect 633 -700 667 -698
rect 633 -785 667 -766
rect 891 -596 925 -577
rect 891 -664 925 -662
rect 891 -700 925 -698
rect 891 -785 925 -766
rect 1138 -596 1172 -577
rect 1138 -664 1172 -662
rect 1138 -700 1172 -698
rect 1138 -785 1172 -766
rect 1396 -596 1430 -577
rect 1396 -664 1430 -662
rect 1396 -700 1430 -698
rect 1396 -785 1430 -766
rect 1654 -596 1688 -577
rect 1654 -664 1688 -662
rect 1654 -700 1688 -698
rect 1654 -785 1688 -766
rect 1912 -596 1946 -577
rect 1912 -664 1946 -662
rect 1912 -700 1946 -698
rect 1912 -785 1946 -766
rect 2159 -596 2193 -577
rect 2159 -664 2193 -662
rect 2159 -700 2193 -698
rect 2159 -785 2193 -766
rect 2417 -596 2451 -577
rect 2417 -664 2451 -662
rect 2417 -700 2451 -698
rect 2417 -785 2451 -766
rect 2675 -596 2709 -577
rect 2675 -664 2709 -662
rect 2675 -700 2709 -698
rect 2675 -785 2709 -766
rect 2923 -596 2957 -577
rect 2923 -664 2957 -662
rect 2923 -700 2957 -698
rect 2923 -785 2957 -766
rect 3181 -596 3215 -577
rect 3181 -664 3215 -662
rect 3181 -700 3215 -698
rect 3181 -785 3215 -766
rect 6834 -558 6868 -546
rect 3295 -630 3329 -614
rect 3295 -702 3329 -682
rect 3295 -774 3329 -750
rect -244 -846 -210 -818
rect -244 -918 -210 -886
rect -244 -990 -210 -952
rect -244 -1026 -210 -1024
rect 3409 -596 3443 -577
rect 3409 -664 3443 -662
rect 3409 -700 3443 -698
rect 3409 -785 3443 -766
rect 3667 -596 3701 -577
rect 3667 -664 3701 -662
rect 3667 -700 3701 -698
rect 3667 -785 3701 -766
rect 3915 -596 3949 -577
rect 3915 -664 3949 -662
rect 3915 -700 3949 -698
rect 3915 -785 3949 -766
rect 4173 -596 4207 -577
rect 4173 -664 4207 -662
rect 4173 -700 4207 -698
rect 4173 -785 4207 -766
rect 4431 -596 4465 -577
rect 4431 -664 4465 -662
rect 4431 -700 4465 -698
rect 4431 -785 4465 -766
rect 4678 -596 4712 -577
rect 4678 -664 4712 -662
rect 4678 -700 4712 -698
rect 4678 -785 4712 -766
rect 4936 -596 4970 -577
rect 4936 -664 4970 -662
rect 4936 -700 4970 -698
rect 4936 -785 4970 -766
rect 5194 -596 5228 -577
rect 5194 -664 5228 -662
rect 5194 -700 5228 -698
rect 5194 -785 5228 -766
rect 5452 -596 5486 -577
rect 5452 -664 5486 -662
rect 5452 -700 5486 -698
rect 5452 -785 5486 -766
rect 5699 -596 5733 -577
rect 5699 -664 5733 -662
rect 5699 -700 5733 -698
rect 5699 -785 5733 -766
rect 5957 -596 5991 -577
rect 5957 -664 5991 -662
rect 5957 -700 5991 -698
rect 5957 -785 5991 -766
rect 6215 -596 6249 -577
rect 6215 -664 6249 -662
rect 6215 -700 6249 -698
rect 6215 -785 6249 -766
rect 6462 -596 6496 -577
rect 6462 -664 6496 -662
rect 6462 -700 6496 -698
rect 6462 -785 6496 -766
rect 6720 -596 6754 -577
rect 6720 -664 6754 -662
rect 6720 -700 6754 -698
rect 6720 -785 6754 -766
rect 6834 -630 6868 -614
rect 6834 -702 6868 -682
rect 6834 -774 6868 -750
rect 3295 -846 3329 -818
rect 3295 -918 3329 -886
rect 3295 -990 3329 -952
rect 3295 -1026 3329 -1024
rect 6834 -846 6868 -818
rect 6834 -918 6868 -886
rect 6834 -990 6868 -952
rect 6834 -1026 6868 -1024
rect -244 -1060 -59 -1026
rect -25 -1060 9 -1026
rect 43 -1060 77 -1026
rect 111 -1060 145 -1026
rect 179 -1060 213 -1026
rect 247 -1060 281 -1026
rect 315 -1060 349 -1026
rect 383 -1060 417 -1026
rect 451 -1060 485 -1026
rect 519 -1060 553 -1026
rect 587 -1060 621 -1026
rect 655 -1060 689 -1026
rect 723 -1060 757 -1026
rect 791 -1060 825 -1026
rect 859 -1060 893 -1026
rect 927 -1060 961 -1026
rect 995 -1060 1029 -1026
rect 1063 -1060 1097 -1026
rect 1131 -1060 1165 -1026
rect 1199 -1060 1233 -1026
rect 1267 -1060 1301 -1026
rect 1335 -1060 1369 -1026
rect 1403 -1060 1437 -1026
rect 1471 -1060 1505 -1026
rect 1539 -1060 1573 -1026
rect 1607 -1060 1641 -1026
rect 1675 -1060 1709 -1026
rect 1743 -1060 1777 -1026
rect 1811 -1060 1845 -1026
rect 1879 -1060 1913 -1026
rect 1947 -1060 1981 -1026
rect 2015 -1060 2049 -1026
rect 2083 -1060 2117 -1026
rect 2151 -1060 2185 -1026
rect 2219 -1060 2253 -1026
rect 2287 -1060 2321 -1026
rect 2355 -1060 2389 -1026
rect 2423 -1060 2457 -1026
rect 2491 -1060 2525 -1026
rect 2559 -1060 2593 -1026
rect 2627 -1060 2661 -1026
rect 2695 -1060 2729 -1026
rect 2763 -1060 2797 -1026
rect 2831 -1060 2865 -1026
rect 2899 -1060 2933 -1026
rect 2967 -1060 3001 -1026
rect 3035 -1060 3069 -1026
rect 3103 -1060 3137 -1026
rect 3171 -1060 3453 -1026
rect 3487 -1060 3521 -1026
rect 3555 -1060 3589 -1026
rect 3623 -1060 3657 -1026
rect 3691 -1060 3725 -1026
rect 3759 -1060 3793 -1026
rect 3827 -1060 3861 -1026
rect 3895 -1060 3929 -1026
rect 3963 -1060 3997 -1026
rect 4031 -1060 4065 -1026
rect 4099 -1060 4133 -1026
rect 4167 -1060 4201 -1026
rect 4235 -1060 4269 -1026
rect 4303 -1060 4337 -1026
rect 4371 -1060 4405 -1026
rect 4439 -1060 4473 -1026
rect 4507 -1060 4541 -1026
rect 4575 -1060 4609 -1026
rect 4643 -1060 4677 -1026
rect 4711 -1060 4745 -1026
rect 4779 -1060 4813 -1026
rect 4847 -1060 4881 -1026
rect 4915 -1060 4949 -1026
rect 4983 -1060 5017 -1026
rect 5051 -1060 5085 -1026
rect 5119 -1060 5153 -1026
rect 5187 -1060 5221 -1026
rect 5255 -1060 5289 -1026
rect 5323 -1060 5357 -1026
rect 5391 -1060 5425 -1026
rect 5459 -1060 5493 -1026
rect 5527 -1060 5561 -1026
rect 5595 -1060 5629 -1026
rect 5663 -1060 5697 -1026
rect 5731 -1060 5765 -1026
rect 5799 -1060 5833 -1026
rect 5867 -1060 5901 -1026
rect 5935 -1060 5969 -1026
rect 6003 -1060 6037 -1026
rect 6071 -1060 6105 -1026
rect 6139 -1060 6173 -1026
rect 6207 -1060 6241 -1026
rect 6275 -1060 6309 -1026
rect 6343 -1060 6377 -1026
rect 6411 -1060 6445 -1026
rect 6479 -1060 6513 -1026
rect 6547 -1060 6581 -1026
rect 6615 -1060 6649 -1026
rect 6683 -1060 6868 -1026
rect -244 -1062 -210 -1060
rect -244 -1134 -210 -1096
rect -244 -1200 -210 -1168
rect -244 -1268 -210 -1240
rect 3295 -1062 3329 -1060
rect 3295 -1134 3329 -1096
rect 3295 -1200 3329 -1168
rect 3295 -1268 3329 -1240
rect -244 -1336 -210 -1312
rect -244 -1404 -210 -1384
rect -244 -1472 -210 -1456
rect -130 -1320 -96 -1301
rect -130 -1388 -96 -1386
rect -130 -1424 -96 -1422
rect -130 -1509 -96 -1490
rect 128 -1320 162 -1301
rect 128 -1388 162 -1386
rect 128 -1424 162 -1422
rect 128 -1509 162 -1490
rect 375 -1320 409 -1301
rect 375 -1388 409 -1386
rect 375 -1424 409 -1422
rect 375 -1509 409 -1490
rect 633 -1320 667 -1301
rect 633 -1388 667 -1386
rect 633 -1424 667 -1422
rect 633 -1509 667 -1490
rect 891 -1320 925 -1301
rect 891 -1388 925 -1386
rect 891 -1424 925 -1422
rect 891 -1509 925 -1490
rect 1138 -1320 1172 -1301
rect 1138 -1388 1172 -1386
rect 1138 -1424 1172 -1422
rect 1138 -1509 1172 -1490
rect 1396 -1320 1430 -1301
rect 1396 -1388 1430 -1386
rect 1396 -1424 1430 -1422
rect 1396 -1509 1430 -1490
rect 1654 -1320 1688 -1301
rect 1654 -1388 1688 -1386
rect 1654 -1424 1688 -1422
rect 1654 -1509 1688 -1490
rect 1912 -1320 1946 -1301
rect 1912 -1388 1946 -1386
rect 1912 -1424 1946 -1422
rect 1912 -1509 1946 -1490
rect 2159 -1320 2193 -1301
rect 2159 -1388 2193 -1386
rect 2159 -1424 2193 -1422
rect 2159 -1509 2193 -1490
rect 2417 -1320 2451 -1301
rect 2417 -1388 2451 -1386
rect 2417 -1424 2451 -1422
rect 2417 -1509 2451 -1490
rect 2675 -1320 2709 -1301
rect 2675 -1388 2709 -1386
rect 2675 -1424 2709 -1422
rect 2675 -1509 2709 -1490
rect 2923 -1320 2957 -1301
rect 2923 -1388 2957 -1386
rect 2923 -1424 2957 -1422
rect 2923 -1509 2957 -1490
rect 3181 -1320 3215 -1301
rect 3181 -1388 3215 -1386
rect 3181 -1424 3215 -1422
rect 3181 -1509 3215 -1490
rect 6834 -1062 6868 -1060
rect 6834 -1134 6868 -1096
rect 6834 -1200 6868 -1168
rect 6834 -1268 6868 -1240
rect 3295 -1336 3329 -1312
rect 3295 -1404 3329 -1384
rect 3295 -1472 3329 -1456
rect -244 -1540 -210 -1528
rect 3409 -1320 3443 -1301
rect 3409 -1388 3443 -1386
rect 3409 -1424 3443 -1422
rect 3409 -1509 3443 -1490
rect 3667 -1320 3701 -1301
rect 3667 -1388 3701 -1386
rect 3667 -1424 3701 -1422
rect 3667 -1509 3701 -1490
rect 3915 -1320 3949 -1301
rect 3915 -1388 3949 -1386
rect 3915 -1424 3949 -1422
rect 3915 -1509 3949 -1490
rect 4173 -1320 4207 -1301
rect 4173 -1388 4207 -1386
rect 4173 -1424 4207 -1422
rect 4173 -1509 4207 -1490
rect 4431 -1320 4465 -1301
rect 4431 -1388 4465 -1386
rect 4431 -1424 4465 -1422
rect 4431 -1509 4465 -1490
rect 4678 -1320 4712 -1301
rect 4678 -1388 4712 -1386
rect 4678 -1424 4712 -1422
rect 4678 -1509 4712 -1490
rect 4936 -1320 4970 -1301
rect 4936 -1388 4970 -1386
rect 4936 -1424 4970 -1422
rect 4936 -1509 4970 -1490
rect 5194 -1320 5228 -1301
rect 5194 -1388 5228 -1386
rect 5194 -1424 5228 -1422
rect 5194 -1509 5228 -1490
rect 5452 -1320 5486 -1301
rect 5452 -1388 5486 -1386
rect 5452 -1424 5486 -1422
rect 5452 -1509 5486 -1490
rect 5699 -1320 5733 -1301
rect 5699 -1388 5733 -1386
rect 5699 -1424 5733 -1422
rect 5699 -1509 5733 -1490
rect 5957 -1320 5991 -1301
rect 5957 -1388 5991 -1386
rect 5957 -1424 5991 -1422
rect 5957 -1509 5991 -1490
rect 6215 -1320 6249 -1301
rect 6215 -1388 6249 -1386
rect 6215 -1424 6249 -1422
rect 6215 -1509 6249 -1490
rect 6462 -1320 6496 -1301
rect 6462 -1388 6496 -1386
rect 6462 -1424 6496 -1422
rect 6462 -1509 6496 -1490
rect 6720 -1320 6754 -1301
rect 6720 -1388 6754 -1386
rect 6720 -1424 6754 -1422
rect 6720 -1509 6754 -1490
rect 6834 -1336 6868 -1312
rect 6834 -1404 6868 -1384
rect 6834 -1472 6868 -1456
rect 3295 -1540 3329 -1528
rect -84 -1577 -37 -1543
rect -1 -1577 33 -1543
rect 69 -1577 116 -1543
rect 421 -1577 468 -1543
rect 504 -1577 538 -1543
rect 574 -1577 621 -1543
rect 679 -1577 726 -1543
rect 762 -1577 796 -1543
rect 832 -1577 879 -1543
rect 1184 -1577 1231 -1543
rect 1267 -1577 1301 -1543
rect 1337 -1577 1384 -1543
rect 1442 -1577 1489 -1543
rect 1525 -1577 1559 -1543
rect 1595 -1577 1642 -1543
rect 1700 -1577 1747 -1543
rect 1783 -1577 1817 -1543
rect 1853 -1577 1900 -1543
rect 2205 -1577 2252 -1543
rect 2288 -1577 2322 -1543
rect 2358 -1577 2405 -1543
rect 2463 -1577 2510 -1543
rect 2546 -1577 2580 -1543
rect 2616 -1577 2663 -1543
rect 2969 -1577 3016 -1543
rect 3052 -1577 3086 -1543
rect 3122 -1577 3169 -1543
rect 6834 -1540 6868 -1528
rect -244 -1608 -210 -1600
rect -244 -1676 -210 -1672
rect -244 -1782 -210 -1778
rect -244 -1854 -210 -1846
rect 3455 -1577 3502 -1543
rect 3538 -1577 3572 -1543
rect 3608 -1577 3655 -1543
rect 3961 -1577 4008 -1543
rect 4044 -1577 4078 -1543
rect 4114 -1577 4161 -1543
rect 4219 -1577 4266 -1543
rect 4302 -1577 4336 -1543
rect 4372 -1577 4419 -1543
rect 4724 -1577 4771 -1543
rect 4807 -1577 4841 -1543
rect 4877 -1577 4924 -1543
rect 4982 -1577 5029 -1543
rect 5065 -1577 5099 -1543
rect 5135 -1577 5182 -1543
rect 5240 -1577 5287 -1543
rect 5323 -1577 5357 -1543
rect 5393 -1577 5440 -1543
rect 5745 -1577 5792 -1543
rect 5828 -1577 5862 -1543
rect 5898 -1577 5945 -1543
rect 6003 -1577 6050 -1543
rect 6086 -1577 6120 -1543
rect 6156 -1577 6203 -1543
rect 6508 -1577 6555 -1543
rect 6591 -1577 6625 -1543
rect 6661 -1577 6708 -1543
rect 3295 -1608 3329 -1600
rect 3295 -1676 3329 -1672
rect 3295 -1782 3329 -1778
rect 3295 -1854 3329 -1846
rect -244 -1926 -210 -1914
rect -84 -1940 -37 -1906
rect -1 -1940 33 -1906
rect 69 -1940 116 -1906
rect 421 -1940 468 -1906
rect 504 -1940 538 -1906
rect 574 -1940 621 -1906
rect 679 -1940 726 -1906
rect 762 -1940 796 -1906
rect 832 -1940 879 -1906
rect 1184 -1940 1231 -1906
rect 1267 -1940 1301 -1906
rect 1337 -1940 1384 -1906
rect 1442 -1940 1489 -1906
rect 1525 -1940 1559 -1906
rect 1595 -1940 1642 -1906
rect 1700 -1940 1747 -1906
rect 1783 -1940 1817 -1906
rect 1853 -1940 1900 -1906
rect 2205 -1940 2252 -1906
rect 2288 -1940 2322 -1906
rect 2358 -1940 2405 -1906
rect 2463 -1940 2510 -1906
rect 2546 -1940 2580 -1906
rect 2616 -1940 2663 -1906
rect 2969 -1940 3016 -1906
rect 3052 -1940 3086 -1906
rect 3122 -1940 3169 -1906
rect 6834 -1608 6868 -1600
rect 6834 -1676 6868 -1672
rect 6834 -1782 6868 -1778
rect 6834 -1854 6868 -1846
rect 3295 -1926 3329 -1914
rect 3455 -1940 3502 -1906
rect 3538 -1940 3572 -1906
rect 3608 -1940 3655 -1906
rect 3961 -1940 4008 -1906
rect 4044 -1940 4078 -1906
rect 4114 -1940 4161 -1906
rect 4219 -1940 4266 -1906
rect 4302 -1940 4336 -1906
rect 4372 -1940 4419 -1906
rect 4724 -1940 4771 -1906
rect 4807 -1940 4841 -1906
rect 4877 -1940 4924 -1906
rect 4982 -1940 5029 -1906
rect 5065 -1940 5099 -1906
rect 5135 -1940 5182 -1906
rect 5240 -1940 5287 -1906
rect 5323 -1940 5357 -1906
rect 5393 -1940 5440 -1906
rect 5745 -1940 5792 -1906
rect 5828 -1940 5862 -1906
rect 5898 -1940 5945 -1906
rect 6003 -1940 6050 -1906
rect 6086 -1940 6120 -1906
rect 6156 -1940 6203 -1906
rect 6508 -1940 6555 -1906
rect 6591 -1940 6625 -1906
rect 6661 -1940 6708 -1906
rect 6834 -1926 6868 -1914
rect -244 -1998 -210 -1982
rect -244 -2070 -210 -2050
rect -244 -2142 -210 -2118
rect -130 -1993 -96 -1974
rect -130 -2061 -96 -2059
rect -130 -2097 -96 -2095
rect -130 -2182 -96 -2163
rect 128 -1993 162 -1974
rect 128 -2061 162 -2059
rect 128 -2097 162 -2095
rect 128 -2182 162 -2163
rect 375 -1993 409 -1974
rect 375 -2061 409 -2059
rect 375 -2097 409 -2095
rect 375 -2182 409 -2163
rect 633 -1993 667 -1974
rect 633 -2061 667 -2059
rect 633 -2097 667 -2095
rect 633 -2182 667 -2163
rect 891 -1993 925 -1974
rect 891 -2061 925 -2059
rect 891 -2097 925 -2095
rect 891 -2182 925 -2163
rect 1138 -1993 1172 -1974
rect 1138 -2061 1172 -2059
rect 1138 -2097 1172 -2095
rect 1138 -2182 1172 -2163
rect 1396 -1993 1430 -1974
rect 1396 -2061 1430 -2059
rect 1396 -2097 1430 -2095
rect 1396 -2182 1430 -2163
rect 1654 -1993 1688 -1974
rect 1654 -2061 1688 -2059
rect 1654 -2097 1688 -2095
rect 1654 -2182 1688 -2163
rect 1912 -1993 1946 -1974
rect 1912 -2061 1946 -2059
rect 1912 -2097 1946 -2095
rect 1912 -2182 1946 -2163
rect 2159 -1993 2193 -1974
rect 2159 -2061 2193 -2059
rect 2159 -2097 2193 -2095
rect 2159 -2182 2193 -2163
rect 2417 -1993 2451 -1974
rect 2417 -2061 2451 -2059
rect 2417 -2097 2451 -2095
rect 2417 -2182 2451 -2163
rect 2675 -1993 2709 -1974
rect 2675 -2061 2709 -2059
rect 2675 -2097 2709 -2095
rect 2675 -2182 2709 -2163
rect 2923 -1993 2957 -1974
rect 2923 -2061 2957 -2059
rect 2923 -2097 2957 -2095
rect 2923 -2182 2957 -2163
rect 3181 -1993 3215 -1974
rect 3181 -2061 3215 -2059
rect 3181 -2097 3215 -2095
rect 3181 -2182 3215 -2163
rect 3295 -1998 3329 -1982
rect 3295 -2070 3329 -2050
rect 3295 -2142 3329 -2118
rect -244 -2214 -210 -2186
rect -244 -2286 -210 -2254
rect -244 -2356 -210 -2322
rect -244 -2424 -210 -2392
rect 3409 -1993 3443 -1974
rect 3409 -2061 3443 -2059
rect 3409 -2097 3443 -2095
rect 3409 -2182 3443 -2163
rect 3667 -1993 3701 -1974
rect 3667 -2061 3701 -2059
rect 3667 -2097 3701 -2095
rect 3667 -2182 3701 -2163
rect 3915 -1993 3949 -1974
rect 3915 -2061 3949 -2059
rect 3915 -2097 3949 -2095
rect 3915 -2182 3949 -2163
rect 4173 -1993 4207 -1974
rect 4173 -2061 4207 -2059
rect 4173 -2097 4207 -2095
rect 4173 -2182 4207 -2163
rect 4431 -1993 4465 -1974
rect 4431 -2061 4465 -2059
rect 4431 -2097 4465 -2095
rect 4431 -2182 4465 -2163
rect 4678 -1993 4712 -1974
rect 4678 -2061 4712 -2059
rect 4678 -2097 4712 -2095
rect 4678 -2182 4712 -2163
rect 4936 -1993 4970 -1974
rect 4936 -2061 4970 -2059
rect 4936 -2097 4970 -2095
rect 4936 -2182 4970 -2163
rect 5194 -1993 5228 -1974
rect 5194 -2061 5228 -2059
rect 5194 -2097 5228 -2095
rect 5194 -2182 5228 -2163
rect 5452 -1993 5486 -1974
rect 5452 -2061 5486 -2059
rect 5452 -2097 5486 -2095
rect 5452 -2182 5486 -2163
rect 5699 -1993 5733 -1974
rect 5699 -2061 5733 -2059
rect 5699 -2097 5733 -2095
rect 5699 -2182 5733 -2163
rect 5957 -1993 5991 -1974
rect 5957 -2061 5991 -2059
rect 5957 -2097 5991 -2095
rect 5957 -2182 5991 -2163
rect 6215 -1993 6249 -1974
rect 6215 -2061 6249 -2059
rect 6215 -2097 6249 -2095
rect 6215 -2182 6249 -2163
rect 6462 -1993 6496 -1974
rect 6462 -2061 6496 -2059
rect 6462 -2097 6496 -2095
rect 6462 -2182 6496 -2163
rect 6720 -1993 6754 -1974
rect 6720 -2061 6754 -2059
rect 6720 -2097 6754 -2095
rect 6720 -2182 6754 -2163
rect 6834 -1998 6868 -1982
rect 6834 -2070 6868 -2050
rect 6834 -2142 6868 -2118
rect 3295 -2214 3329 -2186
rect 3295 -2286 3329 -2254
rect 3295 -2356 3329 -2322
rect 3295 -2424 3329 -2392
rect 6834 -2214 6868 -2186
rect 6834 -2286 6868 -2254
rect 6834 -2356 6868 -2322
rect 6834 -2424 6868 -2392
rect -210 -2458 -59 -2424
rect -25 -2458 9 -2424
rect 43 -2458 77 -2424
rect 111 -2458 145 -2424
rect 179 -2458 213 -2424
rect 247 -2458 281 -2424
rect 315 -2458 349 -2424
rect 383 -2458 417 -2424
rect 451 -2458 485 -2424
rect 519 -2458 553 -2424
rect 587 -2458 621 -2424
rect 655 -2458 689 -2424
rect 723 -2458 757 -2424
rect 791 -2458 825 -2424
rect 859 -2458 893 -2424
rect 927 -2458 961 -2424
rect 995 -2458 1029 -2424
rect 1063 -2458 1097 -2424
rect 1131 -2458 1165 -2424
rect 1199 -2458 1233 -2424
rect 1267 -2458 1301 -2424
rect 1335 -2458 1369 -2424
rect 1403 -2458 1437 -2424
rect 1471 -2458 1505 -2424
rect 1539 -2458 1573 -2424
rect 1607 -2458 1641 -2424
rect 1675 -2458 1709 -2424
rect 1743 -2458 1777 -2424
rect 1811 -2458 1845 -2424
rect 1879 -2458 1913 -2424
rect 1947 -2458 1981 -2424
rect 2015 -2458 2049 -2424
rect 2083 -2458 2117 -2424
rect 2151 -2458 2185 -2424
rect 2219 -2458 2253 -2424
rect 2287 -2458 2321 -2424
rect 2355 -2458 2389 -2424
rect 2423 -2458 2457 -2424
rect 2491 -2458 2525 -2424
rect 2559 -2458 2593 -2424
rect 2627 -2458 2661 -2424
rect 2695 -2458 2729 -2424
rect 2763 -2458 2797 -2424
rect 2831 -2458 2865 -2424
rect 2899 -2458 2933 -2424
rect 2967 -2458 3001 -2424
rect 3035 -2458 3069 -2424
rect 3103 -2458 3137 -2424
rect 3171 -2458 3295 -2424
rect 3329 -2458 3453 -2424
rect 3487 -2458 3521 -2424
rect 3555 -2458 3589 -2424
rect 3623 -2458 3657 -2424
rect 3691 -2458 3725 -2424
rect 3759 -2458 3793 -2424
rect 3827 -2458 3861 -2424
rect 3895 -2458 3929 -2424
rect 3963 -2458 3997 -2424
rect 4031 -2458 4065 -2424
rect 4099 -2458 4133 -2424
rect 4167 -2458 4201 -2424
rect 4235 -2458 4269 -2424
rect 4303 -2458 4337 -2424
rect 4371 -2458 4405 -2424
rect 4439 -2458 4473 -2424
rect 4507 -2458 4541 -2424
rect 4575 -2458 4609 -2424
rect 4643 -2458 4677 -2424
rect 4711 -2458 4745 -2424
rect 4779 -2458 4813 -2424
rect 4847 -2458 4881 -2424
rect 4915 -2458 4949 -2424
rect 4983 -2458 5017 -2424
rect 5051 -2458 5085 -2424
rect 5119 -2458 5153 -2424
rect 5187 -2458 5221 -2424
rect 5255 -2458 5289 -2424
rect 5323 -2458 5357 -2424
rect 5391 -2458 5425 -2424
rect 5459 -2458 5493 -2424
rect 5527 -2458 5561 -2424
rect 5595 -2458 5629 -2424
rect 5663 -2458 5697 -2424
rect 5731 -2458 5765 -2424
rect 5799 -2458 5833 -2424
rect 5867 -2458 5901 -2424
rect 5935 -2458 5969 -2424
rect 6003 -2458 6037 -2424
rect 6071 -2458 6105 -2424
rect 6139 -2458 6173 -2424
rect 6207 -2458 6241 -2424
rect 6275 -2458 6309 -2424
rect 6343 -2458 6377 -2424
rect 6411 -2458 6445 -2424
rect 6479 -2458 6513 -2424
rect 6547 -2458 6581 -2424
rect 6615 -2458 6649 -2424
rect 6683 -2458 6834 -2424
rect -244 -2492 -210 -2464
rect -244 -2560 -210 -2536
rect -244 -2628 -210 -2608
rect -244 -2696 -210 -2680
rect 3295 -2492 3329 -2464
rect 3295 -2560 3329 -2536
rect 3295 -2628 3329 -2608
rect 3295 -2696 3329 -2680
rect -244 -2764 -210 -2752
rect -244 -2832 -210 -2824
rect -244 -2900 -210 -2896
rect -130 -2719 -96 -2700
rect -130 -2787 -96 -2785
rect -130 -2823 -96 -2821
rect -130 -2908 -96 -2889
rect 128 -2719 162 -2700
rect 128 -2787 162 -2785
rect 128 -2823 162 -2821
rect 128 -2908 162 -2889
rect 375 -2719 409 -2700
rect 375 -2787 409 -2785
rect 375 -2823 409 -2821
rect 375 -2908 409 -2889
rect 633 -2719 667 -2700
rect 633 -2787 667 -2785
rect 633 -2823 667 -2821
rect 633 -2908 667 -2889
rect 891 -2719 925 -2700
rect 891 -2787 925 -2785
rect 891 -2823 925 -2821
rect 891 -2908 925 -2889
rect 1138 -2719 1172 -2700
rect 1138 -2787 1172 -2785
rect 1138 -2823 1172 -2821
rect 1138 -2908 1172 -2889
rect 1396 -2719 1430 -2700
rect 1396 -2787 1430 -2785
rect 1396 -2823 1430 -2821
rect 1396 -2908 1430 -2889
rect 1654 -2719 1688 -2700
rect 1654 -2787 1688 -2785
rect 1654 -2823 1688 -2821
rect 1654 -2908 1688 -2889
rect 1912 -2719 1946 -2700
rect 1912 -2787 1946 -2785
rect 1912 -2823 1946 -2821
rect 1912 -2908 1946 -2889
rect 2159 -2719 2193 -2700
rect 2159 -2787 2193 -2785
rect 2159 -2823 2193 -2821
rect 2159 -2908 2193 -2889
rect 2417 -2719 2451 -2700
rect 2417 -2787 2451 -2785
rect 2417 -2823 2451 -2821
rect 2417 -2908 2451 -2889
rect 2675 -2719 2709 -2700
rect 2675 -2787 2709 -2785
rect 2675 -2823 2709 -2821
rect 2675 -2908 2709 -2889
rect 2923 -2719 2957 -2700
rect 2923 -2787 2957 -2785
rect 2923 -2823 2957 -2821
rect 2923 -2908 2957 -2889
rect 3181 -2719 3215 -2700
rect 3181 -2787 3215 -2785
rect 3181 -2823 3215 -2821
rect 3181 -2908 3215 -2889
rect 6834 -2492 6868 -2464
rect 6834 -2560 6868 -2536
rect 6834 -2628 6868 -2608
rect 6834 -2696 6868 -2680
rect 3295 -2764 3329 -2752
rect 3295 -2832 3329 -2824
rect 3295 -2900 3329 -2896
rect 3409 -2719 3443 -2700
rect 3409 -2787 3443 -2785
rect 3409 -2823 3443 -2821
rect 3409 -2908 3443 -2889
rect 3667 -2719 3701 -2700
rect 3667 -2787 3701 -2785
rect 3667 -2823 3701 -2821
rect 3667 -2908 3701 -2889
rect 3915 -2719 3949 -2700
rect 3915 -2787 3949 -2785
rect 3915 -2823 3949 -2821
rect 3915 -2908 3949 -2889
rect 4173 -2719 4207 -2700
rect 4173 -2787 4207 -2785
rect 4173 -2823 4207 -2821
rect 4173 -2908 4207 -2889
rect 4431 -2719 4465 -2700
rect 4431 -2787 4465 -2785
rect 4431 -2823 4465 -2821
rect 4431 -2908 4465 -2889
rect 4678 -2719 4712 -2700
rect 4678 -2787 4712 -2785
rect 4678 -2823 4712 -2821
rect 4678 -2908 4712 -2889
rect 4936 -2719 4970 -2700
rect 4936 -2787 4970 -2785
rect 4936 -2823 4970 -2821
rect 4936 -2908 4970 -2889
rect 5194 -2719 5228 -2700
rect 5194 -2787 5228 -2785
rect 5194 -2823 5228 -2821
rect 5194 -2908 5228 -2889
rect 5452 -2719 5486 -2700
rect 5452 -2787 5486 -2785
rect 5452 -2823 5486 -2821
rect 5452 -2908 5486 -2889
rect 5699 -2719 5733 -2700
rect 5699 -2787 5733 -2785
rect 5699 -2823 5733 -2821
rect 5699 -2908 5733 -2889
rect 5957 -2719 5991 -2700
rect 5957 -2787 5991 -2785
rect 5957 -2823 5991 -2821
rect 5957 -2908 5991 -2889
rect 6215 -2719 6249 -2700
rect 6215 -2787 6249 -2785
rect 6215 -2823 6249 -2821
rect 6215 -2908 6249 -2889
rect 6462 -2719 6496 -2700
rect 6462 -2787 6496 -2785
rect 6462 -2823 6496 -2821
rect 6462 -2908 6496 -2889
rect 6720 -2719 6754 -2700
rect 6720 -2787 6754 -2785
rect 6720 -2823 6754 -2821
rect 6720 -2908 6754 -2889
rect 6834 -2764 6868 -2752
rect 6834 -2832 6868 -2824
rect 6834 -2900 6868 -2896
rect -244 -3041 -210 -2968
rect -84 -2976 -37 -2942
rect -1 -2976 33 -2942
rect 69 -2976 116 -2942
rect 421 -2976 468 -2942
rect 504 -2976 538 -2942
rect 574 -2976 621 -2942
rect 679 -2976 726 -2942
rect 762 -2976 796 -2942
rect 832 -2976 879 -2942
rect 1184 -2976 1231 -2942
rect 1267 -2976 1301 -2942
rect 1337 -2976 1384 -2942
rect 1442 -2976 1489 -2942
rect 1525 -2976 1559 -2942
rect 1595 -2976 1642 -2942
rect 1700 -2976 1747 -2942
rect 1783 -2976 1817 -2942
rect 1853 -2976 1900 -2942
rect 2205 -2976 2252 -2942
rect 2288 -2976 2322 -2942
rect 2358 -2976 2405 -2942
rect 2463 -2976 2510 -2942
rect 2546 -2976 2580 -2942
rect 2616 -2976 2663 -2942
rect 2969 -2976 3016 -2942
rect 3052 -2976 3086 -2942
rect 3122 -2976 3169 -2942
rect 3295 -3041 3329 -2968
rect 3455 -2976 3502 -2942
rect 3538 -2976 3572 -2942
rect 3608 -2976 3655 -2942
rect 3961 -2976 4008 -2942
rect 4044 -2976 4078 -2942
rect 4114 -2976 4161 -2942
rect 4219 -2976 4266 -2942
rect 4302 -2976 4336 -2942
rect 4372 -2976 4419 -2942
rect 4724 -2976 4771 -2942
rect 4807 -2976 4841 -2942
rect 4877 -2976 4924 -2942
rect 4982 -2976 5029 -2942
rect 5065 -2976 5099 -2942
rect 5135 -2976 5182 -2942
rect 5240 -2976 5287 -2942
rect 5323 -2976 5357 -2942
rect 5393 -2976 5440 -2942
rect 5745 -2976 5792 -2942
rect 5828 -2976 5862 -2942
rect 5898 -2976 5945 -2942
rect 6003 -2976 6050 -2942
rect 6086 -2976 6120 -2942
rect 6156 -2976 6203 -2942
rect 6508 -2976 6555 -2942
rect 6591 -2976 6625 -2942
rect 6661 -2976 6708 -2942
rect 6834 -3041 6868 -2968
rect -244 -3075 -80 -3041
rect -25 -3075 -8 -3041
rect 43 -3075 64 -3041
rect 111 -3075 136 -3041
rect 179 -3075 208 -3041
rect 247 -3075 280 -3041
rect 315 -3075 349 -3041
rect 386 -3075 417 -3041
rect 458 -3075 485 -3041
rect 530 -3075 553 -3041
rect 602 -3075 621 -3041
rect 674 -3075 689 -3041
rect 746 -3075 757 -3041
rect 818 -3075 825 -3041
rect 890 -3075 893 -3041
rect 927 -3075 928 -3041
rect 995 -3075 1000 -3041
rect 1063 -3075 1072 -3041
rect 1131 -3075 1144 -3041
rect 1199 -3075 1216 -3041
rect 1267 -3075 1288 -3041
rect 1335 -3075 1360 -3041
rect 1403 -3075 1432 -3041
rect 1471 -3075 1504 -3041
rect 1539 -3075 1573 -3041
rect 1610 -3075 1641 -3041
rect 1682 -3075 1709 -3041
rect 1754 -3075 1777 -3041
rect 1826 -3075 1845 -3041
rect 1898 -3075 1913 -3041
rect 1970 -3075 1981 -3041
rect 2042 -3075 2049 -3041
rect 2114 -3075 2117 -3041
rect 2151 -3075 2152 -3041
rect 2219 -3075 2224 -3041
rect 2287 -3075 2296 -3041
rect 2355 -3075 2368 -3041
rect 2423 -3075 2440 -3041
rect 2491 -3075 2512 -3041
rect 2559 -3075 2584 -3041
rect 2627 -3075 2656 -3041
rect 2695 -3075 2728 -3041
rect 2763 -3075 2797 -3041
rect 2834 -3075 2865 -3041
rect 2906 -3075 2933 -3041
rect 2978 -3075 3001 -3041
rect 3050 -3075 3069 -3041
rect 3122 -3075 3137 -3041
rect 3194 -3075 3430 -3041
rect 3487 -3075 3502 -3041
rect 3555 -3075 3574 -3041
rect 3623 -3075 3646 -3041
rect 3691 -3075 3718 -3041
rect 3759 -3075 3790 -3041
rect 3827 -3075 3861 -3041
rect 3896 -3075 3929 -3041
rect 3968 -3075 3997 -3041
rect 4040 -3075 4065 -3041
rect 4112 -3075 4133 -3041
rect 4184 -3075 4201 -3041
rect 4256 -3075 4269 -3041
rect 4328 -3075 4337 -3041
rect 4400 -3075 4405 -3041
rect 4472 -3075 4473 -3041
rect 4507 -3075 4510 -3041
rect 4575 -3075 4582 -3041
rect 4643 -3075 4654 -3041
rect 4711 -3075 4726 -3041
rect 4779 -3075 4798 -3041
rect 4847 -3075 4870 -3041
rect 4915 -3075 4942 -3041
rect 4983 -3075 5014 -3041
rect 5051 -3075 5085 -3041
rect 5120 -3075 5153 -3041
rect 5192 -3075 5221 -3041
rect 5264 -3075 5289 -3041
rect 5336 -3075 5357 -3041
rect 5408 -3075 5425 -3041
rect 5480 -3075 5493 -3041
rect 5552 -3075 5561 -3041
rect 5624 -3075 5629 -3041
rect 5696 -3075 5697 -3041
rect 5731 -3075 5734 -3041
rect 5799 -3075 5806 -3041
rect 5867 -3075 5878 -3041
rect 5935 -3075 5950 -3041
rect 6003 -3075 6022 -3041
rect 6071 -3075 6094 -3041
rect 6139 -3075 6166 -3041
rect 6207 -3075 6238 -3041
rect 6275 -3075 6309 -3041
rect 6344 -3075 6377 -3041
rect 6416 -3075 6445 -3041
rect 6488 -3075 6513 -3041
rect 6560 -3075 6581 -3041
rect 6632 -3075 6649 -3041
rect 6704 -3075 6868 -3041
<< viali >>
rect -80 955 -59 989
rect -59 955 -46 989
rect -8 955 9 989
rect 9 955 26 989
rect 64 955 77 989
rect 77 955 98 989
rect 136 955 145 989
rect 145 955 170 989
rect 208 955 213 989
rect 213 955 242 989
rect 280 955 281 989
rect 281 955 314 989
rect 352 955 383 989
rect 383 955 386 989
rect 424 955 451 989
rect 451 955 458 989
rect 496 955 519 989
rect 519 955 530 989
rect 568 955 587 989
rect 587 955 602 989
rect 640 955 655 989
rect 655 955 674 989
rect 712 955 723 989
rect 723 955 746 989
rect 784 955 791 989
rect 791 955 818 989
rect 856 955 859 989
rect 859 955 890 989
rect 928 955 961 989
rect 961 955 962 989
rect 1000 955 1029 989
rect 1029 955 1034 989
rect 1072 955 1097 989
rect 1097 955 1106 989
rect 1144 955 1165 989
rect 1165 955 1178 989
rect 1216 955 1233 989
rect 1233 955 1250 989
rect 1288 955 1301 989
rect 1301 955 1322 989
rect 1360 955 1369 989
rect 1369 955 1394 989
rect 1432 955 1437 989
rect 1437 955 1466 989
rect 1504 955 1505 989
rect 1505 955 1538 989
rect 1576 955 1607 989
rect 1607 955 1610 989
rect 1648 955 1675 989
rect 1675 955 1682 989
rect 1720 955 1743 989
rect 1743 955 1754 989
rect 1792 955 1811 989
rect 1811 955 1826 989
rect 1864 955 1879 989
rect 1879 955 1898 989
rect 1936 955 1947 989
rect 1947 955 1970 989
rect 2008 955 2015 989
rect 2015 955 2042 989
rect 2080 955 2083 989
rect 2083 955 2114 989
rect 2152 955 2185 989
rect 2185 955 2186 989
rect 2224 955 2253 989
rect 2253 955 2258 989
rect 2296 955 2321 989
rect 2321 955 2330 989
rect 2368 955 2389 989
rect 2389 955 2402 989
rect 2440 955 2457 989
rect 2457 955 2474 989
rect 2512 955 2525 989
rect 2525 955 2546 989
rect 2584 955 2593 989
rect 2593 955 2618 989
rect 2656 955 2661 989
rect 2661 955 2690 989
rect 2728 955 2729 989
rect 2729 955 2762 989
rect 2800 955 2831 989
rect 2831 955 2834 989
rect 2872 955 2899 989
rect 2899 955 2906 989
rect 2944 955 2967 989
rect 2967 955 2978 989
rect 3016 955 3035 989
rect 3035 955 3050 989
rect 3088 955 3103 989
rect 3103 955 3122 989
rect 3160 955 3171 989
rect 3171 955 3194 989
rect 3430 955 3453 989
rect 3453 955 3464 989
rect 3502 955 3521 989
rect 3521 955 3536 989
rect 3574 955 3589 989
rect 3589 955 3608 989
rect 3646 955 3657 989
rect 3657 955 3680 989
rect 3718 955 3725 989
rect 3725 955 3752 989
rect 3790 955 3793 989
rect 3793 955 3824 989
rect 3862 955 3895 989
rect 3895 955 3896 989
rect 3934 955 3963 989
rect 3963 955 3968 989
rect 4006 955 4031 989
rect 4031 955 4040 989
rect 4078 955 4099 989
rect 4099 955 4112 989
rect 4150 955 4167 989
rect 4167 955 4184 989
rect 4222 955 4235 989
rect 4235 955 4256 989
rect 4294 955 4303 989
rect 4303 955 4328 989
rect 4366 955 4371 989
rect 4371 955 4400 989
rect 4438 955 4439 989
rect 4439 955 4472 989
rect 4510 955 4541 989
rect 4541 955 4544 989
rect 4582 955 4609 989
rect 4609 955 4616 989
rect 4654 955 4677 989
rect 4677 955 4688 989
rect 4726 955 4745 989
rect 4745 955 4760 989
rect 4798 955 4813 989
rect 4813 955 4832 989
rect 4870 955 4881 989
rect 4881 955 4904 989
rect 4942 955 4949 989
rect 4949 955 4976 989
rect 5014 955 5017 989
rect 5017 955 5048 989
rect 5086 955 5119 989
rect 5119 955 5120 989
rect 5158 955 5187 989
rect 5187 955 5192 989
rect 5230 955 5255 989
rect 5255 955 5264 989
rect 5302 955 5323 989
rect 5323 955 5336 989
rect 5374 955 5391 989
rect 5391 955 5408 989
rect 5446 955 5459 989
rect 5459 955 5480 989
rect 5518 955 5527 989
rect 5527 955 5552 989
rect 5590 955 5595 989
rect 5595 955 5624 989
rect 5662 955 5663 989
rect 5663 955 5696 989
rect 5734 955 5765 989
rect 5765 955 5768 989
rect 5806 955 5833 989
rect 5833 955 5840 989
rect 5878 955 5901 989
rect 5901 955 5912 989
rect 5950 955 5969 989
rect 5969 955 5984 989
rect 6022 955 6037 989
rect 6037 955 6056 989
rect 6094 955 6105 989
rect 6105 955 6128 989
rect 6166 955 6173 989
rect 6173 955 6200 989
rect 6238 955 6241 989
rect 6241 955 6272 989
rect 6310 955 6343 989
rect 6343 955 6344 989
rect 6382 955 6411 989
rect 6411 955 6416 989
rect 6454 955 6479 989
rect 6479 955 6488 989
rect 6526 955 6547 989
rect 6547 955 6560 989
rect 6598 955 6615 989
rect 6615 955 6632 989
rect 6670 955 6683 989
rect 6683 955 6704 989
rect -244 848 -210 882
rect -37 856 -35 890
rect -35 856 -3 890
rect 35 856 67 890
rect 67 856 69 890
rect 468 856 470 890
rect 470 856 502 890
rect 540 856 572 890
rect 572 856 574 890
rect 726 856 728 890
rect 728 856 760 890
rect 798 856 830 890
rect 830 856 832 890
rect 1231 856 1233 890
rect 1233 856 1265 890
rect 1303 856 1335 890
rect 1335 856 1337 890
rect 1489 856 1491 890
rect 1491 856 1523 890
rect 1561 856 1593 890
rect 1593 856 1595 890
rect 1747 856 1749 890
rect 1749 856 1781 890
rect 1819 856 1851 890
rect 1851 856 1853 890
rect 2252 856 2254 890
rect 2254 856 2286 890
rect 2324 856 2356 890
rect 2356 856 2358 890
rect 2510 856 2512 890
rect 2512 856 2544 890
rect 2582 856 2614 890
rect 2614 856 2616 890
rect 3016 856 3018 890
rect 3018 856 3050 890
rect 3088 856 3120 890
rect 3120 856 3122 890
rect 3295 848 3329 882
rect 3502 856 3504 890
rect 3504 856 3536 890
rect 3574 856 3606 890
rect 3606 856 3608 890
rect 4008 856 4010 890
rect 4010 856 4042 890
rect 4080 856 4112 890
rect 4112 856 4114 890
rect 4266 856 4268 890
rect 4268 856 4300 890
rect 4338 856 4370 890
rect 4370 856 4372 890
rect 4771 856 4773 890
rect 4773 856 4805 890
rect 4843 856 4875 890
rect 4875 856 4877 890
rect 5029 856 5031 890
rect 5031 856 5063 890
rect 5101 856 5133 890
rect 5133 856 5135 890
rect 5287 856 5289 890
rect 5289 856 5321 890
rect 5359 856 5391 890
rect 5391 856 5393 890
rect 5792 856 5794 890
rect 5794 856 5826 890
rect 5864 856 5896 890
rect 5896 856 5898 890
rect 6050 856 6052 890
rect 6052 856 6084 890
rect 6122 856 6154 890
rect 6154 856 6156 890
rect 6555 856 6557 890
rect 6557 856 6589 890
rect 6627 856 6659 890
rect 6659 856 6661 890
rect -244 780 -210 810
rect -244 776 -210 780
rect -244 712 -210 738
rect -244 704 -210 712
rect -244 644 -210 666
rect -244 632 -210 644
rect -130 769 -96 771
rect -130 737 -96 769
rect -130 667 -96 699
rect -130 665 -96 667
rect 128 769 162 771
rect 128 737 162 769
rect 128 667 162 699
rect 128 665 162 667
rect 375 769 409 771
rect 375 737 409 769
rect 375 667 409 699
rect 375 665 409 667
rect 633 769 667 771
rect 633 737 667 769
rect 633 667 667 699
rect 633 665 667 667
rect 891 769 925 771
rect 891 737 925 769
rect 891 667 925 699
rect 891 665 925 667
rect 1138 769 1172 771
rect 1138 737 1172 769
rect 1138 667 1172 699
rect 1138 665 1172 667
rect 1396 769 1430 771
rect 1396 737 1430 769
rect 1396 667 1430 699
rect 1396 665 1430 667
rect 1654 769 1688 771
rect 1654 737 1688 769
rect 1654 667 1688 699
rect 1654 665 1688 667
rect 1912 769 1946 771
rect 1912 737 1946 769
rect 1912 667 1946 699
rect 1912 665 1946 667
rect 2159 769 2193 771
rect 2159 737 2193 769
rect 2159 667 2193 699
rect 2159 665 2193 667
rect 2417 769 2451 771
rect 2417 737 2451 769
rect 2417 667 2451 699
rect 2417 665 2451 667
rect 2675 769 2709 771
rect 2675 737 2709 769
rect 2675 667 2709 699
rect 2675 665 2709 667
rect 2923 769 2957 771
rect 2923 737 2957 769
rect 2923 667 2957 699
rect 2923 665 2957 667
rect 3181 769 3215 771
rect 3181 737 3215 769
rect 3181 667 3215 699
rect 3181 665 3215 667
rect 6834 848 6868 882
rect 3295 780 3329 810
rect 3295 776 3329 780
rect 3295 712 3329 738
rect 3295 704 3329 712
rect 3295 644 3329 666
rect 3295 632 3329 644
rect -244 576 -210 594
rect -244 560 -210 576
rect -244 508 -210 522
rect -244 488 -210 508
rect -244 440 -210 450
rect -244 416 -210 440
rect -244 372 -210 378
rect 3409 769 3443 771
rect 3409 737 3443 769
rect 3409 667 3443 699
rect 3409 665 3443 667
rect 3667 769 3701 771
rect 3667 737 3701 769
rect 3667 667 3701 699
rect 3667 665 3701 667
rect 3915 769 3949 771
rect 3915 737 3949 769
rect 3915 667 3949 699
rect 3915 665 3949 667
rect 4173 769 4207 771
rect 4173 737 4207 769
rect 4173 667 4207 699
rect 4173 665 4207 667
rect 4431 769 4465 771
rect 4431 737 4465 769
rect 4431 667 4465 699
rect 4431 665 4465 667
rect 4678 769 4712 771
rect 4678 737 4712 769
rect 4678 667 4712 699
rect 4678 665 4712 667
rect 4936 769 4970 771
rect 4936 737 4970 769
rect 4936 667 4970 699
rect 4936 665 4970 667
rect 5194 769 5228 771
rect 5194 737 5228 769
rect 5194 667 5228 699
rect 5194 665 5228 667
rect 5452 769 5486 771
rect 5452 737 5486 769
rect 5452 667 5486 699
rect 5452 665 5486 667
rect 5699 769 5733 771
rect 5699 737 5733 769
rect 5699 667 5733 699
rect 5699 665 5733 667
rect 5957 769 5991 771
rect 5957 737 5991 769
rect 5957 667 5991 699
rect 5957 665 5991 667
rect 6215 769 6249 771
rect 6215 737 6249 769
rect 6215 667 6249 699
rect 6215 665 6249 667
rect 6462 769 6496 771
rect 6462 737 6496 769
rect 6462 667 6496 699
rect 6462 665 6496 667
rect 6720 769 6754 771
rect 6720 737 6754 769
rect 6720 667 6754 699
rect 6720 665 6754 667
rect 6834 780 6868 810
rect 6834 776 6868 780
rect 6834 712 6868 738
rect 6834 704 6868 712
rect 6834 644 6868 666
rect 6834 632 6868 644
rect 3295 576 3329 594
rect 3295 560 3329 576
rect 3295 508 3329 522
rect 3295 488 3329 508
rect 3295 440 3329 450
rect 3295 416 3329 440
rect 3295 372 3329 378
rect 6834 576 6868 594
rect 6834 560 6868 576
rect 6834 508 6868 522
rect 6834 488 6868 508
rect 6834 440 6868 450
rect 6834 416 6868 440
rect 6834 372 6868 378
rect -244 344 -210 372
rect 3295 344 3329 372
rect 6834 344 6868 372
rect -244 304 -210 306
rect -244 272 -210 304
rect -244 202 -210 234
rect -244 200 -210 202
rect -244 134 -210 162
rect -244 128 -210 134
rect 3295 304 3329 306
rect 3295 272 3329 304
rect 3295 202 3329 234
rect 3295 200 3329 202
rect 3295 134 3329 162
rect 3295 128 3329 134
rect -244 66 -210 90
rect -244 56 -210 66
rect -244 -2 -210 18
rect -244 -16 -210 -2
rect -244 -70 -210 -54
rect -244 -88 -210 -70
rect -130 43 -96 45
rect -130 11 -96 43
rect -130 -59 -96 -27
rect -130 -61 -96 -59
rect 128 43 162 45
rect 128 11 162 43
rect 128 -59 162 -27
rect 128 -61 162 -59
rect 375 43 409 45
rect 375 11 409 43
rect 375 -59 409 -27
rect 375 -61 409 -59
rect 633 43 667 45
rect 633 11 667 43
rect 633 -59 667 -27
rect 633 -61 667 -59
rect 891 43 925 45
rect 891 11 925 43
rect 891 -59 925 -27
rect 891 -61 925 -59
rect 1138 43 1172 45
rect 1138 11 1172 43
rect 1138 -59 1172 -27
rect 1138 -61 1172 -59
rect 1396 43 1430 45
rect 1396 11 1430 43
rect 1396 -59 1430 -27
rect 1396 -61 1430 -59
rect 1654 43 1688 45
rect 1654 11 1688 43
rect 1654 -59 1688 -27
rect 1654 -61 1688 -59
rect 1912 43 1946 45
rect 1912 11 1946 43
rect 1912 -59 1946 -27
rect 1912 -61 1946 -59
rect 2159 43 2193 45
rect 2159 11 2193 43
rect 2159 -59 2193 -27
rect 2159 -61 2193 -59
rect 2417 43 2451 45
rect 2417 11 2451 43
rect 2417 -59 2451 -27
rect 2417 -61 2451 -59
rect 2675 43 2709 45
rect 2675 11 2709 43
rect 2675 -59 2709 -27
rect 2675 -61 2709 -59
rect 2923 43 2957 45
rect 2923 11 2957 43
rect 2923 -59 2957 -27
rect 2923 -61 2957 -59
rect 3181 43 3215 45
rect 3181 11 3215 43
rect 3181 -59 3215 -27
rect 3181 -61 3215 -59
rect 6834 304 6868 306
rect 6834 272 6868 304
rect 6834 202 6868 234
rect 6834 200 6868 202
rect 6834 134 6868 162
rect 6834 128 6868 134
rect 3295 66 3329 90
rect 3295 56 3329 66
rect 3295 -2 3329 18
rect 3295 -16 3329 -2
rect 3295 -70 3329 -54
rect 3295 -88 3329 -70
rect -244 -138 -210 -126
rect -244 -160 -210 -138
rect 3409 43 3443 45
rect 3409 11 3443 43
rect 3409 -59 3443 -27
rect 3409 -61 3443 -59
rect 3667 43 3701 45
rect 3667 11 3701 43
rect 3667 -59 3701 -27
rect 3667 -61 3701 -59
rect 3915 43 3949 45
rect 3915 11 3949 43
rect 3915 -59 3949 -27
rect 3915 -61 3949 -59
rect 4173 43 4207 45
rect 4173 11 4207 43
rect 4173 -59 4207 -27
rect 4173 -61 4207 -59
rect 4431 43 4465 45
rect 4431 11 4465 43
rect 4431 -59 4465 -27
rect 4431 -61 4465 -59
rect 4678 43 4712 45
rect 4678 11 4712 43
rect 4678 -59 4712 -27
rect 4678 -61 4712 -59
rect 4936 43 4970 45
rect 4936 11 4970 43
rect 4936 -59 4970 -27
rect 4936 -61 4970 -59
rect 5194 43 5228 45
rect 5194 11 5228 43
rect 5194 -59 5228 -27
rect 5194 -61 5228 -59
rect 5452 43 5486 45
rect 5452 11 5486 43
rect 5452 -59 5486 -27
rect 5452 -61 5486 -59
rect 5699 43 5733 45
rect 5699 11 5733 43
rect 5699 -59 5733 -27
rect 5699 -61 5733 -59
rect 5957 43 5991 45
rect 5957 11 5991 43
rect 5957 -59 5991 -27
rect 5957 -61 5991 -59
rect 6215 43 6249 45
rect 6215 11 6249 43
rect 6215 -59 6249 -27
rect 6215 -61 6249 -59
rect 6462 43 6496 45
rect 6462 11 6496 43
rect 6462 -59 6496 -27
rect 6462 -61 6496 -59
rect 6720 43 6754 45
rect 6720 11 6754 43
rect 6720 -59 6754 -27
rect 6720 -61 6754 -59
rect 6834 66 6868 90
rect 6834 56 6868 66
rect 6834 -2 6868 18
rect 6834 -16 6868 -2
rect 6834 -70 6868 -54
rect 6834 -88 6868 -70
rect 3295 -138 3329 -126
rect -37 -180 -35 -146
rect -35 -180 -3 -146
rect 35 -180 67 -146
rect 67 -180 69 -146
rect 468 -180 470 -146
rect 470 -180 502 -146
rect 540 -180 572 -146
rect 572 -180 574 -146
rect 726 -180 728 -146
rect 728 -180 760 -146
rect 798 -180 830 -146
rect 830 -180 832 -146
rect 1231 -180 1233 -146
rect 1233 -180 1265 -146
rect 1303 -180 1335 -146
rect 1335 -180 1337 -146
rect 1489 -180 1491 -146
rect 1491 -180 1523 -146
rect 1561 -180 1593 -146
rect 1593 -180 1595 -146
rect 1747 -180 1749 -146
rect 1749 -180 1781 -146
rect 1819 -180 1851 -146
rect 1851 -180 1853 -146
rect 2252 -180 2254 -146
rect 2254 -180 2286 -146
rect 2324 -180 2356 -146
rect 2356 -180 2358 -146
rect 2510 -180 2512 -146
rect 2512 -180 2544 -146
rect 2582 -180 2614 -146
rect 2614 -180 2616 -146
rect 3016 -180 3018 -146
rect 3018 -180 3050 -146
rect 3088 -180 3120 -146
rect 3120 -180 3122 -146
rect 3295 -160 3329 -138
rect 6834 -138 6868 -126
rect -244 -206 -210 -198
rect -244 -232 -210 -206
rect -244 -274 -210 -270
rect -244 -304 -210 -274
rect -244 -376 -210 -342
rect -244 -444 -210 -414
rect -244 -448 -210 -444
rect -244 -512 -210 -486
rect 3502 -180 3504 -146
rect 3504 -180 3536 -146
rect 3574 -180 3606 -146
rect 3606 -180 3608 -146
rect 4008 -180 4010 -146
rect 4010 -180 4042 -146
rect 4080 -180 4112 -146
rect 4112 -180 4114 -146
rect 4266 -180 4268 -146
rect 4268 -180 4300 -146
rect 4338 -180 4370 -146
rect 4370 -180 4372 -146
rect 4771 -180 4773 -146
rect 4773 -180 4805 -146
rect 4843 -180 4875 -146
rect 4875 -180 4877 -146
rect 5029 -180 5031 -146
rect 5031 -180 5063 -146
rect 5101 -180 5133 -146
rect 5133 -180 5135 -146
rect 5287 -180 5289 -146
rect 5289 -180 5321 -146
rect 5359 -180 5391 -146
rect 5391 -180 5393 -146
rect 5792 -180 5794 -146
rect 5794 -180 5826 -146
rect 5864 -180 5896 -146
rect 5896 -180 5898 -146
rect 6050 -180 6052 -146
rect 6052 -180 6084 -146
rect 6122 -180 6154 -146
rect 6154 -180 6156 -146
rect 6555 -180 6557 -146
rect 6557 -180 6589 -146
rect 6627 -180 6659 -146
rect 6659 -180 6661 -146
rect 6834 -160 6868 -138
rect 3295 -206 3329 -198
rect 3295 -232 3329 -206
rect 3295 -274 3329 -270
rect 3295 -304 3329 -274
rect 3295 -376 3329 -342
rect 3295 -444 3329 -414
rect 3295 -448 3329 -444
rect -244 -520 -210 -512
rect -37 -543 -35 -509
rect -35 -543 -3 -509
rect 35 -543 67 -509
rect 67 -543 69 -509
rect 468 -543 470 -509
rect 470 -543 502 -509
rect 540 -543 572 -509
rect 572 -543 574 -509
rect 726 -543 728 -509
rect 728 -543 760 -509
rect 798 -543 830 -509
rect 830 -543 832 -509
rect 1231 -543 1233 -509
rect 1233 -543 1265 -509
rect 1303 -543 1335 -509
rect 1335 -543 1337 -509
rect 1489 -543 1491 -509
rect 1491 -543 1523 -509
rect 1561 -543 1593 -509
rect 1593 -543 1595 -509
rect 1747 -543 1749 -509
rect 1749 -543 1781 -509
rect 1819 -543 1851 -509
rect 1851 -543 1853 -509
rect 2252 -543 2254 -509
rect 2254 -543 2286 -509
rect 2324 -543 2356 -509
rect 2356 -543 2358 -509
rect 2510 -543 2512 -509
rect 2512 -543 2544 -509
rect 2582 -543 2614 -509
rect 2614 -543 2616 -509
rect 3016 -543 3018 -509
rect 3018 -543 3050 -509
rect 3088 -543 3120 -509
rect 3120 -543 3122 -509
rect 3295 -512 3329 -486
rect 6834 -206 6868 -198
rect 6834 -232 6868 -206
rect 6834 -274 6868 -270
rect 6834 -304 6868 -274
rect 6834 -376 6868 -342
rect 6834 -444 6868 -414
rect 6834 -448 6868 -444
rect 3295 -520 3329 -512
rect -244 -580 -210 -558
rect 3502 -543 3504 -509
rect 3504 -543 3536 -509
rect 3574 -543 3606 -509
rect 3606 -543 3608 -509
rect 4008 -543 4010 -509
rect 4010 -543 4042 -509
rect 4080 -543 4112 -509
rect 4112 -543 4114 -509
rect 4266 -543 4268 -509
rect 4268 -543 4300 -509
rect 4338 -543 4370 -509
rect 4370 -543 4372 -509
rect 4771 -543 4773 -509
rect 4773 -543 4805 -509
rect 4843 -543 4875 -509
rect 4875 -543 4877 -509
rect 5029 -543 5031 -509
rect 5031 -543 5063 -509
rect 5101 -543 5133 -509
rect 5133 -543 5135 -509
rect 5287 -543 5289 -509
rect 5289 -543 5321 -509
rect 5359 -543 5391 -509
rect 5391 -543 5393 -509
rect 5792 -543 5794 -509
rect 5794 -543 5826 -509
rect 5864 -543 5896 -509
rect 5896 -543 5898 -509
rect 6050 -543 6052 -509
rect 6052 -543 6084 -509
rect 6122 -543 6154 -509
rect 6154 -543 6156 -509
rect 6555 -543 6557 -509
rect 6557 -543 6589 -509
rect 6627 -543 6659 -509
rect 6659 -543 6661 -509
rect 6834 -512 6868 -486
rect 6834 -520 6868 -512
rect -244 -592 -210 -580
rect -244 -648 -210 -630
rect -244 -664 -210 -648
rect -244 -716 -210 -702
rect -244 -736 -210 -716
rect -244 -784 -210 -774
rect -244 -808 -210 -784
rect -130 -630 -96 -628
rect -130 -662 -96 -630
rect -130 -732 -96 -700
rect -130 -734 -96 -732
rect 128 -630 162 -628
rect 128 -662 162 -630
rect 128 -732 162 -700
rect 128 -734 162 -732
rect 375 -630 409 -628
rect 375 -662 409 -630
rect 375 -732 409 -700
rect 375 -734 409 -732
rect 633 -630 667 -628
rect 633 -662 667 -630
rect 633 -732 667 -700
rect 633 -734 667 -732
rect 891 -630 925 -628
rect 891 -662 925 -630
rect 891 -732 925 -700
rect 891 -734 925 -732
rect 1138 -630 1172 -628
rect 1138 -662 1172 -630
rect 1138 -732 1172 -700
rect 1138 -734 1172 -732
rect 1396 -630 1430 -628
rect 1396 -662 1430 -630
rect 1396 -732 1430 -700
rect 1396 -734 1430 -732
rect 1654 -630 1688 -628
rect 1654 -662 1688 -630
rect 1654 -732 1688 -700
rect 1654 -734 1688 -732
rect 1912 -630 1946 -628
rect 1912 -662 1946 -630
rect 1912 -732 1946 -700
rect 1912 -734 1946 -732
rect 2159 -630 2193 -628
rect 2159 -662 2193 -630
rect 2159 -732 2193 -700
rect 2159 -734 2193 -732
rect 2417 -630 2451 -628
rect 2417 -662 2451 -630
rect 2417 -732 2451 -700
rect 2417 -734 2451 -732
rect 2675 -630 2709 -628
rect 2675 -662 2709 -630
rect 2675 -732 2709 -700
rect 2675 -734 2709 -732
rect 2923 -630 2957 -628
rect 2923 -662 2957 -630
rect 2923 -732 2957 -700
rect 2923 -734 2957 -732
rect 3181 -630 3215 -628
rect 3181 -662 3215 -630
rect 3181 -732 3215 -700
rect 3181 -734 3215 -732
rect 3295 -580 3329 -558
rect 3295 -592 3329 -580
rect 3295 -648 3329 -630
rect 3295 -664 3329 -648
rect 3295 -716 3329 -702
rect 3295 -736 3329 -716
rect 3295 -784 3329 -774
rect -244 -852 -210 -846
rect -244 -880 -210 -852
rect -244 -952 -210 -918
rect -244 -1024 -210 -990
rect 3295 -808 3329 -784
rect 3409 -630 3443 -628
rect 3409 -662 3443 -630
rect 3409 -732 3443 -700
rect 3409 -734 3443 -732
rect 3667 -630 3701 -628
rect 3667 -662 3701 -630
rect 3667 -732 3701 -700
rect 3667 -734 3701 -732
rect 3915 -630 3949 -628
rect 3915 -662 3949 -630
rect 3915 -732 3949 -700
rect 3915 -734 3949 -732
rect 4173 -630 4207 -628
rect 4173 -662 4207 -630
rect 4173 -732 4207 -700
rect 4173 -734 4207 -732
rect 4431 -630 4465 -628
rect 4431 -662 4465 -630
rect 4431 -732 4465 -700
rect 4431 -734 4465 -732
rect 4678 -630 4712 -628
rect 4678 -662 4712 -630
rect 4678 -732 4712 -700
rect 4678 -734 4712 -732
rect 4936 -630 4970 -628
rect 4936 -662 4970 -630
rect 4936 -732 4970 -700
rect 4936 -734 4970 -732
rect 5194 -630 5228 -628
rect 5194 -662 5228 -630
rect 5194 -732 5228 -700
rect 5194 -734 5228 -732
rect 5452 -630 5486 -628
rect 5452 -662 5486 -630
rect 5452 -732 5486 -700
rect 5452 -734 5486 -732
rect 5699 -630 5733 -628
rect 5699 -662 5733 -630
rect 5699 -732 5733 -700
rect 5699 -734 5733 -732
rect 5957 -630 5991 -628
rect 5957 -662 5991 -630
rect 5957 -732 5991 -700
rect 5957 -734 5991 -732
rect 6215 -630 6249 -628
rect 6215 -662 6249 -630
rect 6215 -732 6249 -700
rect 6215 -734 6249 -732
rect 6462 -630 6496 -628
rect 6462 -662 6496 -630
rect 6462 -732 6496 -700
rect 6462 -734 6496 -732
rect 6720 -630 6754 -628
rect 6720 -662 6754 -630
rect 6720 -732 6754 -700
rect 6720 -734 6754 -732
rect 6834 -580 6868 -558
rect 6834 -592 6868 -580
rect 6834 -648 6868 -630
rect 6834 -664 6868 -648
rect 6834 -716 6868 -702
rect 6834 -736 6868 -716
rect 6834 -784 6868 -774
rect 3295 -852 3329 -846
rect 3295 -880 3329 -852
rect 3295 -952 3329 -918
rect 3295 -1024 3329 -990
rect 6834 -808 6868 -784
rect 6834 -852 6868 -846
rect 6834 -880 6868 -852
rect 6834 -952 6868 -918
rect 6834 -1024 6868 -990
rect -244 -1096 -210 -1062
rect -244 -1168 -210 -1134
rect -244 -1234 -210 -1206
rect -244 -1240 -210 -1234
rect -244 -1302 -210 -1278
rect 3295 -1096 3329 -1062
rect 3295 -1168 3329 -1134
rect 3295 -1234 3329 -1206
rect 3295 -1240 3329 -1234
rect -244 -1312 -210 -1302
rect -244 -1370 -210 -1350
rect -244 -1384 -210 -1370
rect -244 -1438 -210 -1422
rect -244 -1456 -210 -1438
rect -244 -1506 -210 -1494
rect -244 -1528 -210 -1506
rect -130 -1354 -96 -1352
rect -130 -1386 -96 -1354
rect -130 -1456 -96 -1424
rect -130 -1458 -96 -1456
rect 128 -1354 162 -1352
rect 128 -1386 162 -1354
rect 128 -1456 162 -1424
rect 128 -1458 162 -1456
rect 375 -1354 409 -1352
rect 375 -1386 409 -1354
rect 375 -1456 409 -1424
rect 375 -1458 409 -1456
rect 633 -1354 667 -1352
rect 633 -1386 667 -1354
rect 633 -1456 667 -1424
rect 633 -1458 667 -1456
rect 891 -1354 925 -1352
rect 891 -1386 925 -1354
rect 891 -1456 925 -1424
rect 891 -1458 925 -1456
rect 1138 -1354 1172 -1352
rect 1138 -1386 1172 -1354
rect 1138 -1456 1172 -1424
rect 1138 -1458 1172 -1456
rect 1396 -1354 1430 -1352
rect 1396 -1386 1430 -1354
rect 1396 -1456 1430 -1424
rect 1396 -1458 1430 -1456
rect 1654 -1354 1688 -1352
rect 1654 -1386 1688 -1354
rect 1654 -1456 1688 -1424
rect 1654 -1458 1688 -1456
rect 1912 -1354 1946 -1352
rect 1912 -1386 1946 -1354
rect 1912 -1456 1946 -1424
rect 1912 -1458 1946 -1456
rect 2159 -1354 2193 -1352
rect 2159 -1386 2193 -1354
rect 2159 -1456 2193 -1424
rect 2159 -1458 2193 -1456
rect 2417 -1354 2451 -1352
rect 2417 -1386 2451 -1354
rect 2417 -1456 2451 -1424
rect 2417 -1458 2451 -1456
rect 2675 -1354 2709 -1352
rect 2675 -1386 2709 -1354
rect 2675 -1456 2709 -1424
rect 2675 -1458 2709 -1456
rect 2923 -1354 2957 -1352
rect 2923 -1386 2957 -1354
rect 2923 -1456 2957 -1424
rect 2923 -1458 2957 -1456
rect 3181 -1354 3215 -1352
rect 3181 -1386 3215 -1354
rect 3181 -1456 3215 -1424
rect 3181 -1458 3215 -1456
rect 3295 -1302 3329 -1278
rect 6834 -1096 6868 -1062
rect 6834 -1168 6868 -1134
rect 6834 -1234 6868 -1206
rect 6834 -1240 6868 -1234
rect 3295 -1312 3329 -1302
rect 3295 -1370 3329 -1350
rect 3295 -1384 3329 -1370
rect 3295 -1438 3329 -1422
rect 3295 -1456 3329 -1438
rect 3295 -1506 3329 -1494
rect 3295 -1528 3329 -1506
rect 3409 -1354 3443 -1352
rect 3409 -1386 3443 -1354
rect 3409 -1456 3443 -1424
rect 3409 -1458 3443 -1456
rect 3667 -1354 3701 -1352
rect 3667 -1386 3701 -1354
rect 3667 -1456 3701 -1424
rect 3667 -1458 3701 -1456
rect 3915 -1354 3949 -1352
rect 3915 -1386 3949 -1354
rect 3915 -1456 3949 -1424
rect 3915 -1458 3949 -1456
rect 4173 -1354 4207 -1352
rect 4173 -1386 4207 -1354
rect 4173 -1456 4207 -1424
rect 4173 -1458 4207 -1456
rect 4431 -1354 4465 -1352
rect 4431 -1386 4465 -1354
rect 4431 -1456 4465 -1424
rect 4431 -1458 4465 -1456
rect 4678 -1354 4712 -1352
rect 4678 -1386 4712 -1354
rect 4678 -1456 4712 -1424
rect 4678 -1458 4712 -1456
rect 4936 -1354 4970 -1352
rect 4936 -1386 4970 -1354
rect 4936 -1456 4970 -1424
rect 4936 -1458 4970 -1456
rect 5194 -1354 5228 -1352
rect 5194 -1386 5228 -1354
rect 5194 -1456 5228 -1424
rect 5194 -1458 5228 -1456
rect 5452 -1354 5486 -1352
rect 5452 -1386 5486 -1354
rect 5452 -1456 5486 -1424
rect 5452 -1458 5486 -1456
rect 5699 -1354 5733 -1352
rect 5699 -1386 5733 -1354
rect 5699 -1456 5733 -1424
rect 5699 -1458 5733 -1456
rect 5957 -1354 5991 -1352
rect 5957 -1386 5991 -1354
rect 5957 -1456 5991 -1424
rect 5957 -1458 5991 -1456
rect 6215 -1354 6249 -1352
rect 6215 -1386 6249 -1354
rect 6215 -1456 6249 -1424
rect 6215 -1458 6249 -1456
rect 6462 -1354 6496 -1352
rect 6462 -1386 6496 -1354
rect 6462 -1456 6496 -1424
rect 6462 -1458 6496 -1456
rect 6720 -1354 6754 -1352
rect 6720 -1386 6754 -1354
rect 6720 -1456 6754 -1424
rect 6720 -1458 6754 -1456
rect 6834 -1302 6868 -1278
rect 6834 -1312 6868 -1302
rect 6834 -1370 6868 -1350
rect 6834 -1384 6868 -1370
rect 6834 -1438 6868 -1422
rect 6834 -1456 6868 -1438
rect 6834 -1506 6868 -1494
rect -244 -1574 -210 -1566
rect -244 -1600 -210 -1574
rect -37 -1577 -35 -1543
rect -35 -1577 -3 -1543
rect 35 -1577 67 -1543
rect 67 -1577 69 -1543
rect 468 -1577 470 -1543
rect 470 -1577 502 -1543
rect 540 -1577 572 -1543
rect 572 -1577 574 -1543
rect 726 -1577 728 -1543
rect 728 -1577 760 -1543
rect 798 -1577 830 -1543
rect 830 -1577 832 -1543
rect 1231 -1577 1233 -1543
rect 1233 -1577 1265 -1543
rect 1303 -1577 1335 -1543
rect 1335 -1577 1337 -1543
rect 1489 -1577 1491 -1543
rect 1491 -1577 1523 -1543
rect 1561 -1577 1593 -1543
rect 1593 -1577 1595 -1543
rect 1747 -1577 1749 -1543
rect 1749 -1577 1781 -1543
rect 1819 -1577 1851 -1543
rect 1851 -1577 1853 -1543
rect 2252 -1577 2254 -1543
rect 2254 -1577 2286 -1543
rect 2324 -1577 2356 -1543
rect 2356 -1577 2358 -1543
rect 2510 -1577 2512 -1543
rect 2512 -1577 2544 -1543
rect 2582 -1577 2614 -1543
rect 2614 -1577 2616 -1543
rect 3016 -1577 3018 -1543
rect 3018 -1577 3050 -1543
rect 3088 -1577 3120 -1543
rect 3120 -1577 3122 -1543
rect 6834 -1528 6868 -1506
rect 3295 -1574 3329 -1566
rect -244 -1642 -210 -1638
rect -244 -1672 -210 -1642
rect -244 -1744 -210 -1710
rect -244 -1812 -210 -1782
rect -244 -1816 -210 -1812
rect -244 -1880 -210 -1854
rect -244 -1888 -210 -1880
rect 3295 -1600 3329 -1574
rect 3502 -1577 3504 -1543
rect 3504 -1577 3536 -1543
rect 3574 -1577 3606 -1543
rect 3606 -1577 3608 -1543
rect 4008 -1577 4010 -1543
rect 4010 -1577 4042 -1543
rect 4080 -1577 4112 -1543
rect 4112 -1577 4114 -1543
rect 4266 -1577 4268 -1543
rect 4268 -1577 4300 -1543
rect 4338 -1577 4370 -1543
rect 4370 -1577 4372 -1543
rect 4771 -1577 4773 -1543
rect 4773 -1577 4805 -1543
rect 4843 -1577 4875 -1543
rect 4875 -1577 4877 -1543
rect 5029 -1577 5031 -1543
rect 5031 -1577 5063 -1543
rect 5101 -1577 5133 -1543
rect 5133 -1577 5135 -1543
rect 5287 -1577 5289 -1543
rect 5289 -1577 5321 -1543
rect 5359 -1577 5391 -1543
rect 5391 -1577 5393 -1543
rect 5792 -1577 5794 -1543
rect 5794 -1577 5826 -1543
rect 5864 -1577 5896 -1543
rect 5896 -1577 5898 -1543
rect 6050 -1577 6052 -1543
rect 6052 -1577 6084 -1543
rect 6122 -1577 6154 -1543
rect 6154 -1577 6156 -1543
rect 6555 -1577 6557 -1543
rect 6557 -1577 6589 -1543
rect 6627 -1577 6659 -1543
rect 6659 -1577 6661 -1543
rect 6834 -1574 6868 -1566
rect 3295 -1642 3329 -1638
rect 3295 -1672 3329 -1642
rect 3295 -1744 3329 -1710
rect 3295 -1812 3329 -1782
rect 3295 -1816 3329 -1812
rect 3295 -1880 3329 -1854
rect 3295 -1888 3329 -1880
rect -244 -1948 -210 -1926
rect -37 -1940 -35 -1906
rect -35 -1940 -3 -1906
rect 35 -1940 67 -1906
rect 67 -1940 69 -1906
rect 468 -1940 470 -1906
rect 470 -1940 502 -1906
rect 540 -1940 572 -1906
rect 572 -1940 574 -1906
rect 726 -1940 728 -1906
rect 728 -1940 760 -1906
rect 798 -1940 830 -1906
rect 830 -1940 832 -1906
rect 1231 -1940 1233 -1906
rect 1233 -1940 1265 -1906
rect 1303 -1940 1335 -1906
rect 1335 -1940 1337 -1906
rect 1489 -1940 1491 -1906
rect 1491 -1940 1523 -1906
rect 1561 -1940 1593 -1906
rect 1593 -1940 1595 -1906
rect 1747 -1940 1749 -1906
rect 1749 -1940 1781 -1906
rect 1819 -1940 1851 -1906
rect 1851 -1940 1853 -1906
rect 2252 -1940 2254 -1906
rect 2254 -1940 2286 -1906
rect 2324 -1940 2356 -1906
rect 2356 -1940 2358 -1906
rect 2510 -1940 2512 -1906
rect 2512 -1940 2544 -1906
rect 2582 -1940 2614 -1906
rect 2614 -1940 2616 -1906
rect 3016 -1940 3018 -1906
rect 3018 -1940 3050 -1906
rect 3088 -1940 3120 -1906
rect 3120 -1940 3122 -1906
rect 6834 -1600 6868 -1574
rect 6834 -1642 6868 -1638
rect 6834 -1672 6868 -1642
rect 6834 -1744 6868 -1710
rect 6834 -1812 6868 -1782
rect 6834 -1816 6868 -1812
rect 6834 -1880 6868 -1854
rect 6834 -1888 6868 -1880
rect -244 -1960 -210 -1948
rect 3295 -1948 3329 -1926
rect 3502 -1940 3504 -1906
rect 3504 -1940 3536 -1906
rect 3574 -1940 3606 -1906
rect 3606 -1940 3608 -1906
rect 4008 -1940 4010 -1906
rect 4010 -1940 4042 -1906
rect 4080 -1940 4112 -1906
rect 4112 -1940 4114 -1906
rect 4266 -1940 4268 -1906
rect 4268 -1940 4300 -1906
rect 4338 -1940 4370 -1906
rect 4370 -1940 4372 -1906
rect 4771 -1940 4773 -1906
rect 4773 -1940 4805 -1906
rect 4843 -1940 4875 -1906
rect 4875 -1940 4877 -1906
rect 5029 -1940 5031 -1906
rect 5031 -1940 5063 -1906
rect 5101 -1940 5133 -1906
rect 5133 -1940 5135 -1906
rect 5287 -1940 5289 -1906
rect 5289 -1940 5321 -1906
rect 5359 -1940 5391 -1906
rect 5391 -1940 5393 -1906
rect 5792 -1940 5794 -1906
rect 5794 -1940 5826 -1906
rect 5864 -1940 5896 -1906
rect 5896 -1940 5898 -1906
rect 6050 -1940 6052 -1906
rect 6052 -1940 6084 -1906
rect 6122 -1940 6154 -1906
rect 6154 -1940 6156 -1906
rect 6555 -1940 6557 -1906
rect 6557 -1940 6589 -1906
rect 6627 -1940 6659 -1906
rect 6659 -1940 6661 -1906
rect 3295 -1960 3329 -1948
rect -244 -2016 -210 -1998
rect -244 -2032 -210 -2016
rect -244 -2084 -210 -2070
rect -244 -2104 -210 -2084
rect -244 -2152 -210 -2142
rect -244 -2176 -210 -2152
rect -130 -2027 -96 -2025
rect -130 -2059 -96 -2027
rect -130 -2129 -96 -2097
rect -130 -2131 -96 -2129
rect 128 -2027 162 -2025
rect 128 -2059 162 -2027
rect 128 -2129 162 -2097
rect 128 -2131 162 -2129
rect 375 -2027 409 -2025
rect 375 -2059 409 -2027
rect 375 -2129 409 -2097
rect 375 -2131 409 -2129
rect 633 -2027 667 -2025
rect 633 -2059 667 -2027
rect 633 -2129 667 -2097
rect 633 -2131 667 -2129
rect 891 -2027 925 -2025
rect 891 -2059 925 -2027
rect 891 -2129 925 -2097
rect 891 -2131 925 -2129
rect 1138 -2027 1172 -2025
rect 1138 -2059 1172 -2027
rect 1138 -2129 1172 -2097
rect 1138 -2131 1172 -2129
rect 1396 -2027 1430 -2025
rect 1396 -2059 1430 -2027
rect 1396 -2129 1430 -2097
rect 1396 -2131 1430 -2129
rect 1654 -2027 1688 -2025
rect 1654 -2059 1688 -2027
rect 1654 -2129 1688 -2097
rect 1654 -2131 1688 -2129
rect 1912 -2027 1946 -2025
rect 1912 -2059 1946 -2027
rect 1912 -2129 1946 -2097
rect 1912 -2131 1946 -2129
rect 2159 -2027 2193 -2025
rect 2159 -2059 2193 -2027
rect 2159 -2129 2193 -2097
rect 2159 -2131 2193 -2129
rect 2417 -2027 2451 -2025
rect 2417 -2059 2451 -2027
rect 2417 -2129 2451 -2097
rect 2417 -2131 2451 -2129
rect 2675 -2027 2709 -2025
rect 2675 -2059 2709 -2027
rect 2675 -2129 2709 -2097
rect 2675 -2131 2709 -2129
rect 2923 -2027 2957 -2025
rect 2923 -2059 2957 -2027
rect 2923 -2129 2957 -2097
rect 2923 -2131 2957 -2129
rect 3181 -2027 3215 -2025
rect 3181 -2059 3215 -2027
rect 3181 -2129 3215 -2097
rect 3181 -2131 3215 -2129
rect 6834 -1948 6868 -1926
rect 6834 -1960 6868 -1948
rect 3295 -2016 3329 -1998
rect 3295 -2032 3329 -2016
rect 3295 -2084 3329 -2070
rect 3295 -2104 3329 -2084
rect 3295 -2152 3329 -2142
rect 3295 -2176 3329 -2152
rect -244 -2220 -210 -2214
rect -244 -2248 -210 -2220
rect -244 -2288 -210 -2286
rect -244 -2320 -210 -2288
rect -244 -2390 -210 -2358
rect -244 -2392 -210 -2390
rect 3409 -2027 3443 -2025
rect 3409 -2059 3443 -2027
rect 3409 -2129 3443 -2097
rect 3409 -2131 3443 -2129
rect 3667 -2027 3701 -2025
rect 3667 -2059 3701 -2027
rect 3667 -2129 3701 -2097
rect 3667 -2131 3701 -2129
rect 3915 -2027 3949 -2025
rect 3915 -2059 3949 -2027
rect 3915 -2129 3949 -2097
rect 3915 -2131 3949 -2129
rect 4173 -2027 4207 -2025
rect 4173 -2059 4207 -2027
rect 4173 -2129 4207 -2097
rect 4173 -2131 4207 -2129
rect 4431 -2027 4465 -2025
rect 4431 -2059 4465 -2027
rect 4431 -2129 4465 -2097
rect 4431 -2131 4465 -2129
rect 4678 -2027 4712 -2025
rect 4678 -2059 4712 -2027
rect 4678 -2129 4712 -2097
rect 4678 -2131 4712 -2129
rect 4936 -2027 4970 -2025
rect 4936 -2059 4970 -2027
rect 4936 -2129 4970 -2097
rect 4936 -2131 4970 -2129
rect 5194 -2027 5228 -2025
rect 5194 -2059 5228 -2027
rect 5194 -2129 5228 -2097
rect 5194 -2131 5228 -2129
rect 5452 -2027 5486 -2025
rect 5452 -2059 5486 -2027
rect 5452 -2129 5486 -2097
rect 5452 -2131 5486 -2129
rect 5699 -2027 5733 -2025
rect 5699 -2059 5733 -2027
rect 5699 -2129 5733 -2097
rect 5699 -2131 5733 -2129
rect 5957 -2027 5991 -2025
rect 5957 -2059 5991 -2027
rect 5957 -2129 5991 -2097
rect 5957 -2131 5991 -2129
rect 6215 -2027 6249 -2025
rect 6215 -2059 6249 -2027
rect 6215 -2129 6249 -2097
rect 6215 -2131 6249 -2129
rect 6462 -2027 6496 -2025
rect 6462 -2059 6496 -2027
rect 6462 -2129 6496 -2097
rect 6462 -2131 6496 -2129
rect 6720 -2027 6754 -2025
rect 6720 -2059 6754 -2027
rect 6720 -2129 6754 -2097
rect 6720 -2131 6754 -2129
rect 6834 -2016 6868 -1998
rect 6834 -2032 6868 -2016
rect 6834 -2084 6868 -2070
rect 6834 -2104 6868 -2084
rect 6834 -2152 6868 -2142
rect 6834 -2176 6868 -2152
rect 3295 -2220 3329 -2214
rect 3295 -2248 3329 -2220
rect 3295 -2288 3329 -2286
rect 3295 -2320 3329 -2288
rect 3295 -2390 3329 -2358
rect 3295 -2392 3329 -2390
rect 6834 -2220 6868 -2214
rect 6834 -2248 6868 -2220
rect 6834 -2288 6868 -2286
rect 6834 -2320 6868 -2288
rect 6834 -2390 6868 -2358
rect 6834 -2392 6868 -2390
rect -244 -2458 -210 -2430
rect 3295 -2458 3329 -2430
rect 6834 -2458 6868 -2430
rect -244 -2464 -210 -2458
rect -244 -2526 -210 -2502
rect -244 -2536 -210 -2526
rect -244 -2594 -210 -2574
rect -244 -2608 -210 -2594
rect -244 -2662 -210 -2646
rect -244 -2680 -210 -2662
rect 3295 -2464 3329 -2458
rect 3295 -2526 3329 -2502
rect 3295 -2536 3329 -2526
rect 3295 -2594 3329 -2574
rect 3295 -2608 3329 -2594
rect 3295 -2662 3329 -2646
rect 3295 -2680 3329 -2662
rect -244 -2730 -210 -2718
rect -244 -2752 -210 -2730
rect -244 -2798 -210 -2790
rect -244 -2824 -210 -2798
rect -244 -2866 -210 -2862
rect -244 -2896 -210 -2866
rect -130 -2753 -96 -2751
rect -130 -2785 -96 -2753
rect -130 -2855 -96 -2823
rect -130 -2857 -96 -2855
rect 128 -2753 162 -2751
rect 128 -2785 162 -2753
rect 128 -2855 162 -2823
rect 128 -2857 162 -2855
rect 375 -2753 409 -2751
rect 375 -2785 409 -2753
rect 375 -2855 409 -2823
rect 375 -2857 409 -2855
rect 633 -2753 667 -2751
rect 633 -2785 667 -2753
rect 633 -2855 667 -2823
rect 633 -2857 667 -2855
rect 891 -2753 925 -2751
rect 891 -2785 925 -2753
rect 891 -2855 925 -2823
rect 891 -2857 925 -2855
rect 1138 -2753 1172 -2751
rect 1138 -2785 1172 -2753
rect 1138 -2855 1172 -2823
rect 1138 -2857 1172 -2855
rect 1396 -2753 1430 -2751
rect 1396 -2785 1430 -2753
rect 1396 -2855 1430 -2823
rect 1396 -2857 1430 -2855
rect 1654 -2753 1688 -2751
rect 1654 -2785 1688 -2753
rect 1654 -2855 1688 -2823
rect 1654 -2857 1688 -2855
rect 1912 -2753 1946 -2751
rect 1912 -2785 1946 -2753
rect 1912 -2855 1946 -2823
rect 1912 -2857 1946 -2855
rect 2159 -2753 2193 -2751
rect 2159 -2785 2193 -2753
rect 2159 -2855 2193 -2823
rect 2159 -2857 2193 -2855
rect 2417 -2753 2451 -2751
rect 2417 -2785 2451 -2753
rect 2417 -2855 2451 -2823
rect 2417 -2857 2451 -2855
rect 2675 -2753 2709 -2751
rect 2675 -2785 2709 -2753
rect 2675 -2855 2709 -2823
rect 2675 -2857 2709 -2855
rect 2923 -2753 2957 -2751
rect 2923 -2785 2957 -2753
rect 2923 -2855 2957 -2823
rect 2923 -2857 2957 -2855
rect 3181 -2753 3215 -2751
rect 3181 -2785 3215 -2753
rect 3181 -2855 3215 -2823
rect 3181 -2857 3215 -2855
rect 6834 -2464 6868 -2458
rect 6834 -2526 6868 -2502
rect 6834 -2536 6868 -2526
rect 6834 -2594 6868 -2574
rect 6834 -2608 6868 -2594
rect 6834 -2662 6868 -2646
rect 6834 -2680 6868 -2662
rect 3295 -2730 3329 -2718
rect 3295 -2752 3329 -2730
rect 3295 -2798 3329 -2790
rect 3295 -2824 3329 -2798
rect 3295 -2866 3329 -2862
rect 3295 -2896 3329 -2866
rect -244 -2968 -210 -2934
rect 3409 -2753 3443 -2751
rect 3409 -2785 3443 -2753
rect 3409 -2855 3443 -2823
rect 3409 -2857 3443 -2855
rect 3667 -2753 3701 -2751
rect 3667 -2785 3701 -2753
rect 3667 -2855 3701 -2823
rect 3667 -2857 3701 -2855
rect 3915 -2753 3949 -2751
rect 3915 -2785 3949 -2753
rect 3915 -2855 3949 -2823
rect 3915 -2857 3949 -2855
rect 4173 -2753 4207 -2751
rect 4173 -2785 4207 -2753
rect 4173 -2855 4207 -2823
rect 4173 -2857 4207 -2855
rect 4431 -2753 4465 -2751
rect 4431 -2785 4465 -2753
rect 4431 -2855 4465 -2823
rect 4431 -2857 4465 -2855
rect 4678 -2753 4712 -2751
rect 4678 -2785 4712 -2753
rect 4678 -2855 4712 -2823
rect 4678 -2857 4712 -2855
rect 4936 -2753 4970 -2751
rect 4936 -2785 4970 -2753
rect 4936 -2855 4970 -2823
rect 4936 -2857 4970 -2855
rect 5194 -2753 5228 -2751
rect 5194 -2785 5228 -2753
rect 5194 -2855 5228 -2823
rect 5194 -2857 5228 -2855
rect 5452 -2753 5486 -2751
rect 5452 -2785 5486 -2753
rect 5452 -2855 5486 -2823
rect 5452 -2857 5486 -2855
rect 5699 -2753 5733 -2751
rect 5699 -2785 5733 -2753
rect 5699 -2855 5733 -2823
rect 5699 -2857 5733 -2855
rect 5957 -2753 5991 -2751
rect 5957 -2785 5991 -2753
rect 5957 -2855 5991 -2823
rect 5957 -2857 5991 -2855
rect 6215 -2753 6249 -2751
rect 6215 -2785 6249 -2753
rect 6215 -2855 6249 -2823
rect 6215 -2857 6249 -2855
rect 6462 -2753 6496 -2751
rect 6462 -2785 6496 -2753
rect 6462 -2855 6496 -2823
rect 6462 -2857 6496 -2855
rect 6720 -2753 6754 -2751
rect 6720 -2785 6754 -2753
rect 6720 -2855 6754 -2823
rect 6720 -2857 6754 -2855
rect 6834 -2730 6868 -2718
rect 6834 -2752 6868 -2730
rect 6834 -2798 6868 -2790
rect 6834 -2824 6868 -2798
rect 6834 -2866 6868 -2862
rect 6834 -2896 6868 -2866
rect -37 -2976 -35 -2942
rect -35 -2976 -3 -2942
rect 35 -2976 67 -2942
rect 67 -2976 69 -2942
rect 468 -2976 470 -2942
rect 470 -2976 502 -2942
rect 540 -2976 572 -2942
rect 572 -2976 574 -2942
rect 726 -2976 728 -2942
rect 728 -2976 760 -2942
rect 798 -2976 830 -2942
rect 830 -2976 832 -2942
rect 1231 -2976 1233 -2942
rect 1233 -2976 1265 -2942
rect 1303 -2976 1335 -2942
rect 1335 -2976 1337 -2942
rect 1489 -2976 1491 -2942
rect 1491 -2976 1523 -2942
rect 1561 -2976 1593 -2942
rect 1593 -2976 1595 -2942
rect 1747 -2976 1749 -2942
rect 1749 -2976 1781 -2942
rect 1819 -2976 1851 -2942
rect 1851 -2976 1853 -2942
rect 2252 -2976 2254 -2942
rect 2254 -2976 2286 -2942
rect 2324 -2976 2356 -2942
rect 2356 -2976 2358 -2942
rect 2510 -2976 2512 -2942
rect 2512 -2976 2544 -2942
rect 2582 -2976 2614 -2942
rect 2614 -2976 2616 -2942
rect 3016 -2976 3018 -2942
rect 3018 -2976 3050 -2942
rect 3088 -2976 3120 -2942
rect 3120 -2976 3122 -2942
rect 3295 -2968 3329 -2934
rect 3502 -2976 3504 -2942
rect 3504 -2976 3536 -2942
rect 3574 -2976 3606 -2942
rect 3606 -2976 3608 -2942
rect 4008 -2976 4010 -2942
rect 4010 -2976 4042 -2942
rect 4080 -2976 4112 -2942
rect 4112 -2976 4114 -2942
rect 4266 -2976 4268 -2942
rect 4268 -2976 4300 -2942
rect 4338 -2976 4370 -2942
rect 4370 -2976 4372 -2942
rect 4771 -2976 4773 -2942
rect 4773 -2976 4805 -2942
rect 4843 -2976 4875 -2942
rect 4875 -2976 4877 -2942
rect 5029 -2976 5031 -2942
rect 5031 -2976 5063 -2942
rect 5101 -2976 5133 -2942
rect 5133 -2976 5135 -2942
rect 5287 -2976 5289 -2942
rect 5289 -2976 5321 -2942
rect 5359 -2976 5391 -2942
rect 5391 -2976 5393 -2942
rect 5792 -2976 5794 -2942
rect 5794 -2976 5826 -2942
rect 5864 -2976 5896 -2942
rect 5896 -2976 5898 -2942
rect 6050 -2976 6052 -2942
rect 6052 -2976 6084 -2942
rect 6122 -2976 6154 -2942
rect 6154 -2976 6156 -2942
rect 6555 -2976 6557 -2942
rect 6557 -2976 6589 -2942
rect 6627 -2976 6659 -2942
rect 6659 -2976 6661 -2942
rect 6834 -2968 6868 -2934
rect -80 -3075 -59 -3041
rect -59 -3075 -46 -3041
rect -8 -3075 9 -3041
rect 9 -3075 26 -3041
rect 64 -3075 77 -3041
rect 77 -3075 98 -3041
rect 136 -3075 145 -3041
rect 145 -3075 170 -3041
rect 208 -3075 213 -3041
rect 213 -3075 242 -3041
rect 280 -3075 281 -3041
rect 281 -3075 314 -3041
rect 352 -3075 383 -3041
rect 383 -3075 386 -3041
rect 424 -3075 451 -3041
rect 451 -3075 458 -3041
rect 496 -3075 519 -3041
rect 519 -3075 530 -3041
rect 568 -3075 587 -3041
rect 587 -3075 602 -3041
rect 640 -3075 655 -3041
rect 655 -3075 674 -3041
rect 712 -3075 723 -3041
rect 723 -3075 746 -3041
rect 784 -3075 791 -3041
rect 791 -3075 818 -3041
rect 856 -3075 859 -3041
rect 859 -3075 890 -3041
rect 928 -3075 961 -3041
rect 961 -3075 962 -3041
rect 1000 -3075 1029 -3041
rect 1029 -3075 1034 -3041
rect 1072 -3075 1097 -3041
rect 1097 -3075 1106 -3041
rect 1144 -3075 1165 -3041
rect 1165 -3075 1178 -3041
rect 1216 -3075 1233 -3041
rect 1233 -3075 1250 -3041
rect 1288 -3075 1301 -3041
rect 1301 -3075 1322 -3041
rect 1360 -3075 1369 -3041
rect 1369 -3075 1394 -3041
rect 1432 -3075 1437 -3041
rect 1437 -3075 1466 -3041
rect 1504 -3075 1505 -3041
rect 1505 -3075 1538 -3041
rect 1576 -3075 1607 -3041
rect 1607 -3075 1610 -3041
rect 1648 -3075 1675 -3041
rect 1675 -3075 1682 -3041
rect 1720 -3075 1743 -3041
rect 1743 -3075 1754 -3041
rect 1792 -3075 1811 -3041
rect 1811 -3075 1826 -3041
rect 1864 -3075 1879 -3041
rect 1879 -3075 1898 -3041
rect 1936 -3075 1947 -3041
rect 1947 -3075 1970 -3041
rect 2008 -3075 2015 -3041
rect 2015 -3075 2042 -3041
rect 2080 -3075 2083 -3041
rect 2083 -3075 2114 -3041
rect 2152 -3075 2185 -3041
rect 2185 -3075 2186 -3041
rect 2224 -3075 2253 -3041
rect 2253 -3075 2258 -3041
rect 2296 -3075 2321 -3041
rect 2321 -3075 2330 -3041
rect 2368 -3075 2389 -3041
rect 2389 -3075 2402 -3041
rect 2440 -3075 2457 -3041
rect 2457 -3075 2474 -3041
rect 2512 -3075 2525 -3041
rect 2525 -3075 2546 -3041
rect 2584 -3075 2593 -3041
rect 2593 -3075 2618 -3041
rect 2656 -3075 2661 -3041
rect 2661 -3075 2690 -3041
rect 2728 -3075 2729 -3041
rect 2729 -3075 2762 -3041
rect 2800 -3075 2831 -3041
rect 2831 -3075 2834 -3041
rect 2872 -3075 2899 -3041
rect 2899 -3075 2906 -3041
rect 2944 -3075 2967 -3041
rect 2967 -3075 2978 -3041
rect 3016 -3075 3035 -3041
rect 3035 -3075 3050 -3041
rect 3088 -3075 3103 -3041
rect 3103 -3075 3122 -3041
rect 3160 -3075 3171 -3041
rect 3171 -3075 3194 -3041
rect 3430 -3075 3453 -3041
rect 3453 -3075 3464 -3041
rect 3502 -3075 3521 -3041
rect 3521 -3075 3536 -3041
rect 3574 -3075 3589 -3041
rect 3589 -3075 3608 -3041
rect 3646 -3075 3657 -3041
rect 3657 -3075 3680 -3041
rect 3718 -3075 3725 -3041
rect 3725 -3075 3752 -3041
rect 3790 -3075 3793 -3041
rect 3793 -3075 3824 -3041
rect 3862 -3075 3895 -3041
rect 3895 -3075 3896 -3041
rect 3934 -3075 3963 -3041
rect 3963 -3075 3968 -3041
rect 4006 -3075 4031 -3041
rect 4031 -3075 4040 -3041
rect 4078 -3075 4099 -3041
rect 4099 -3075 4112 -3041
rect 4150 -3075 4167 -3041
rect 4167 -3075 4184 -3041
rect 4222 -3075 4235 -3041
rect 4235 -3075 4256 -3041
rect 4294 -3075 4303 -3041
rect 4303 -3075 4328 -3041
rect 4366 -3075 4371 -3041
rect 4371 -3075 4400 -3041
rect 4438 -3075 4439 -3041
rect 4439 -3075 4472 -3041
rect 4510 -3075 4541 -3041
rect 4541 -3075 4544 -3041
rect 4582 -3075 4609 -3041
rect 4609 -3075 4616 -3041
rect 4654 -3075 4677 -3041
rect 4677 -3075 4688 -3041
rect 4726 -3075 4745 -3041
rect 4745 -3075 4760 -3041
rect 4798 -3075 4813 -3041
rect 4813 -3075 4832 -3041
rect 4870 -3075 4881 -3041
rect 4881 -3075 4904 -3041
rect 4942 -3075 4949 -3041
rect 4949 -3075 4976 -3041
rect 5014 -3075 5017 -3041
rect 5017 -3075 5048 -3041
rect 5086 -3075 5119 -3041
rect 5119 -3075 5120 -3041
rect 5158 -3075 5187 -3041
rect 5187 -3075 5192 -3041
rect 5230 -3075 5255 -3041
rect 5255 -3075 5264 -3041
rect 5302 -3075 5323 -3041
rect 5323 -3075 5336 -3041
rect 5374 -3075 5391 -3041
rect 5391 -3075 5408 -3041
rect 5446 -3075 5459 -3041
rect 5459 -3075 5480 -3041
rect 5518 -3075 5527 -3041
rect 5527 -3075 5552 -3041
rect 5590 -3075 5595 -3041
rect 5595 -3075 5624 -3041
rect 5662 -3075 5663 -3041
rect 5663 -3075 5696 -3041
rect 5734 -3075 5765 -3041
rect 5765 -3075 5768 -3041
rect 5806 -3075 5833 -3041
rect 5833 -3075 5840 -3041
rect 5878 -3075 5901 -3041
rect 5901 -3075 5912 -3041
rect 5950 -3075 5969 -3041
rect 5969 -3075 5984 -3041
rect 6022 -3075 6037 -3041
rect 6037 -3075 6056 -3041
rect 6094 -3075 6105 -3041
rect 6105 -3075 6128 -3041
rect 6166 -3075 6173 -3041
rect 6173 -3075 6200 -3041
rect 6238 -3075 6241 -3041
rect 6241 -3075 6272 -3041
rect 6310 -3075 6343 -3041
rect 6343 -3075 6344 -3041
rect 6382 -3075 6411 -3041
rect 6411 -3075 6416 -3041
rect 6454 -3075 6479 -3041
rect 6479 -3075 6488 -3041
rect 6526 -3075 6547 -3041
rect 6547 -3075 6560 -3041
rect 6598 -3075 6615 -3041
rect 6615 -3075 6632 -3041
rect 6670 -3075 6683 -3041
rect 6683 -3075 6704 -3041
<< metal1 >>
rect -269 989 6893 1014
rect -269 955 -80 989
rect -46 955 -8 989
rect 26 955 64 989
rect 98 955 136 989
rect 170 955 208 989
rect 242 955 280 989
rect 314 955 352 989
rect 386 955 424 989
rect 458 955 496 989
rect 530 955 568 989
rect 602 955 640 989
rect 674 955 712 989
rect 746 955 784 989
rect 818 955 856 989
rect 890 955 928 989
rect 962 955 1000 989
rect 1034 955 1072 989
rect 1106 955 1144 989
rect 1178 955 1216 989
rect 1250 955 1288 989
rect 1322 955 1360 989
rect 1394 955 1432 989
rect 1466 955 1504 989
rect 1538 955 1576 989
rect 1610 955 1648 989
rect 1682 955 1720 989
rect 1754 955 1792 989
rect 1826 955 1864 989
rect 1898 955 1936 989
rect 1970 955 2008 989
rect 2042 955 2080 989
rect 2114 955 2152 989
rect 2186 955 2224 989
rect 2258 955 2296 989
rect 2330 955 2368 989
rect 2402 955 2440 989
rect 2474 955 2512 989
rect 2546 955 2584 989
rect 2618 955 2656 989
rect 2690 955 2728 989
rect 2762 955 2800 989
rect 2834 955 2872 989
rect 2906 955 2944 989
rect 2978 955 3016 989
rect 3050 955 3088 989
rect 3122 955 3160 989
rect 3194 955 3430 989
rect 3464 955 3502 989
rect 3536 955 3574 989
rect 3608 955 3646 989
rect 3680 955 3718 989
rect 3752 955 3790 989
rect 3824 955 3862 989
rect 3896 955 3934 989
rect 3968 955 4006 989
rect 4040 955 4078 989
rect 4112 955 4150 989
rect 4184 955 4222 989
rect 4256 955 4294 989
rect 4328 955 4366 989
rect 4400 955 4438 989
rect 4472 955 4510 989
rect 4544 955 4582 989
rect 4616 955 4654 989
rect 4688 955 4726 989
rect 4760 955 4798 989
rect 4832 955 4870 989
rect 4904 955 4942 989
rect 4976 955 5014 989
rect 5048 955 5086 989
rect 5120 955 5158 989
rect 5192 955 5230 989
rect 5264 955 5302 989
rect 5336 955 5374 989
rect 5408 955 5446 989
rect 5480 955 5518 989
rect 5552 955 5590 989
rect 5624 955 5662 989
rect 5696 955 5734 989
rect 5768 955 5806 989
rect 5840 955 5878 989
rect 5912 955 5950 989
rect 5984 955 6022 989
rect 6056 955 6094 989
rect 6128 955 6166 989
rect 6200 955 6238 989
rect 6272 955 6310 989
rect 6344 955 6382 989
rect 6416 955 6454 989
rect 6488 955 6526 989
rect 6560 955 6598 989
rect 6632 955 6670 989
rect 6704 955 6893 989
rect -269 890 6893 955
rect -269 882 -37 890
rect -269 848 -244 882
rect -210 856 -37 882
rect -3 856 35 890
rect 69 856 468 890
rect 502 856 540 890
rect 574 856 726 890
rect 760 856 798 890
rect 832 856 1231 890
rect 1265 856 1303 890
rect 1337 856 1489 890
rect 1523 856 1561 890
rect 1595 856 1747 890
rect 1781 856 1819 890
rect 1853 856 2252 890
rect 2286 856 2324 890
rect 2358 856 2510 890
rect 2544 856 2582 890
rect 2616 856 3016 890
rect 3050 856 3088 890
rect 3122 882 3502 890
rect 3122 856 3295 882
rect -210 850 3295 856
rect -210 848 168 850
rect -269 810 168 848
rect -269 776 -244 810
rect -210 776 168 810
rect -269 771 168 776
rect -269 738 -130 771
rect -269 704 -244 738
rect -210 737 -130 738
rect -96 737 128 771
rect 162 737 168 771
rect -210 704 168 737
rect -269 699 168 704
rect -269 666 -130 699
rect -269 632 -244 666
rect -210 665 -130 666
rect -96 665 128 699
rect 162 665 168 699
rect -210 632 168 665
rect -269 594 168 632
rect 369 771 415 850
rect 369 737 375 771
rect 409 737 415 771
rect 369 699 415 737
rect 369 665 375 699
rect 409 665 415 699
rect 369 618 415 665
rect 627 771 673 850
rect 627 737 633 771
rect 667 737 673 771
rect 627 699 673 737
rect 627 665 633 699
rect 667 665 673 699
rect 627 618 673 665
rect 885 771 931 850
rect 885 737 891 771
rect 925 737 931 771
rect 885 699 931 737
rect 885 665 891 699
rect 925 665 931 699
rect 885 618 931 665
rect 1132 771 1178 850
rect 1132 737 1138 771
rect 1172 737 1178 771
rect 1132 699 1178 737
rect 1132 665 1138 699
rect 1172 665 1178 699
rect 1132 618 1178 665
rect 1390 771 1436 850
rect 1390 737 1396 771
rect 1430 737 1436 771
rect 1390 699 1436 737
rect 1390 665 1396 699
rect 1430 665 1436 699
rect 1390 618 1436 665
rect 1648 771 1694 850
rect 1648 737 1654 771
rect 1688 737 1694 771
rect 1648 699 1694 737
rect 1648 665 1654 699
rect 1688 665 1694 699
rect 1648 618 1694 665
rect 1906 771 1952 850
rect 1906 737 1912 771
rect 1946 737 1952 771
rect 1906 699 1952 737
rect 1906 665 1912 699
rect 1946 665 1952 699
rect 1906 618 1952 665
rect 2153 771 2199 850
rect 2153 737 2159 771
rect 2193 737 2199 771
rect 2153 699 2199 737
rect 2153 665 2159 699
rect 2193 665 2199 699
rect 2153 618 2199 665
rect 2411 771 2457 850
rect 2411 737 2417 771
rect 2451 737 2457 771
rect 2411 699 2457 737
rect 2411 665 2417 699
rect 2451 665 2457 699
rect 2411 618 2457 665
rect 2669 771 2715 850
rect 2669 737 2675 771
rect 2709 737 2715 771
rect 2669 699 2715 737
rect 2669 665 2675 699
rect 2709 665 2715 699
rect 2669 618 2715 665
rect 2917 848 3295 850
rect 3329 856 3502 882
rect 3536 856 3574 890
rect 3608 856 4008 890
rect 4042 856 4080 890
rect 4114 856 4266 890
rect 4300 856 4338 890
rect 4372 856 4771 890
rect 4805 856 4843 890
rect 4877 856 5029 890
rect 5063 856 5101 890
rect 5135 856 5287 890
rect 5321 856 5359 890
rect 5393 856 5792 890
rect 5826 856 5864 890
rect 5898 856 6050 890
rect 6084 856 6122 890
rect 6156 856 6555 890
rect 6589 856 6627 890
rect 6661 882 6893 890
rect 6661 856 6834 882
rect 3329 850 6834 856
rect 3329 848 3707 850
rect 2917 810 3707 848
rect 2917 776 3295 810
rect 3329 776 3707 810
rect 2917 771 3707 776
rect 2917 737 2923 771
rect 2957 737 3181 771
rect 3215 738 3409 771
rect 3215 737 3295 738
rect 2917 704 3295 737
rect 3329 737 3409 738
rect 3443 737 3667 771
rect 3701 737 3707 771
rect 3329 704 3707 737
rect 2917 699 3707 704
rect 2917 665 2923 699
rect 2957 665 3181 699
rect 3215 666 3409 699
rect 3215 665 3295 666
rect 2917 632 3295 665
rect 3329 665 3409 666
rect 3443 665 3667 699
rect 3701 665 3707 699
rect 3329 632 3707 665
rect -269 560 -244 594
rect -210 560 168 594
rect 2917 594 3707 632
rect 3909 771 3955 850
rect 3909 737 3915 771
rect 3949 737 3955 771
rect 3909 699 3955 737
rect 3909 665 3915 699
rect 3949 665 3955 699
rect 3909 618 3955 665
rect 4167 771 4213 850
rect 4167 737 4173 771
rect 4207 737 4213 771
rect 4167 699 4213 737
rect 4167 665 4173 699
rect 4207 665 4213 699
rect 4167 618 4213 665
rect 4425 771 4471 850
rect 4425 737 4431 771
rect 4465 737 4471 771
rect 4425 699 4471 737
rect 4425 665 4431 699
rect 4465 665 4471 699
rect 4425 618 4471 665
rect 4672 771 4718 850
rect 4672 737 4678 771
rect 4712 737 4718 771
rect 4672 699 4718 737
rect 4672 665 4678 699
rect 4712 665 4718 699
rect 4672 618 4718 665
rect 4930 771 4976 850
rect 4930 737 4936 771
rect 4970 737 4976 771
rect 4930 699 4976 737
rect 4930 665 4936 699
rect 4970 665 4976 699
rect 4930 618 4976 665
rect 5188 771 5234 850
rect 5188 737 5194 771
rect 5228 737 5234 771
rect 5188 699 5234 737
rect 5188 665 5194 699
rect 5228 665 5234 699
rect 5188 618 5234 665
rect 5446 771 5492 850
rect 5446 737 5452 771
rect 5486 737 5492 771
rect 5446 699 5492 737
rect 5446 665 5452 699
rect 5486 665 5492 699
rect 5446 618 5492 665
rect 5693 771 5739 850
rect 5693 737 5699 771
rect 5733 737 5739 771
rect 5693 699 5739 737
rect 5693 665 5699 699
rect 5733 665 5739 699
rect 5693 618 5739 665
rect 5951 771 5997 850
rect 5951 737 5957 771
rect 5991 737 5997 771
rect 5951 699 5997 737
rect 5951 665 5957 699
rect 5991 665 5997 699
rect 5951 618 5997 665
rect 6209 771 6255 850
rect 6209 737 6215 771
rect 6249 737 6255 771
rect 6209 699 6255 737
rect 6209 665 6215 699
rect 6249 665 6255 699
rect 6209 618 6255 665
rect 6456 848 6834 850
rect 6868 848 6893 882
rect 6456 810 6893 848
rect 6456 776 6834 810
rect 6868 776 6893 810
rect 6456 771 6893 776
rect 6456 737 6462 771
rect 6496 737 6720 771
rect 6754 738 6893 771
rect 6754 737 6834 738
rect 6456 704 6834 737
rect 6868 704 6893 738
rect 6456 699 6893 704
rect 6456 665 6462 699
rect 6496 665 6720 699
rect 6754 666 6893 699
rect 6754 665 6834 666
rect 6456 632 6834 665
rect 6868 632 6893 666
rect 2917 560 3295 594
rect 3329 560 3707 594
rect 6456 594 6893 632
rect 6456 560 6834 594
rect 6868 560 6893 594
rect -269 522 168 560
rect -269 488 -244 522
rect -210 488 168 522
rect 1058 552 1254 560
rect 1058 500 1067 552
rect 1119 500 1131 552
rect 1183 500 1195 552
rect 1247 500 1254 552
rect 1058 490 1254 500
rect 1575 552 1771 560
rect 1575 500 1584 552
rect 1636 500 1648 552
rect 1700 500 1712 552
rect 1764 500 1771 552
rect 1575 490 1771 500
rect 2917 522 3707 560
rect -269 450 168 488
rect -269 416 -244 450
rect -210 416 168 450
rect -269 378 168 416
rect -269 344 -244 378
rect -210 344 168 378
rect -269 306 168 344
rect -269 272 -244 306
rect -210 272 168 306
rect -269 234 168 272
rect -269 200 -244 234
rect -210 200 168 234
rect -269 162 168 200
rect -269 128 -244 162
rect -210 128 168 162
rect -269 90 168 128
rect -269 56 -244 90
rect -210 56 168 90
rect -269 45 168 56
rect -269 18 -130 45
rect -269 -16 -244 18
rect -210 11 -130 18
rect -96 11 128 45
rect 162 11 168 45
rect -210 -16 168 11
rect -269 -27 168 -16
rect -269 -54 -130 -27
rect -269 -88 -244 -54
rect -210 -61 -130 -54
rect -96 -61 128 -27
rect 162 -61 168 -27
rect -210 -88 168 -61
rect -269 -126 168 -88
rect 369 436 931 444
rect 369 384 378 436
rect 430 384 442 436
rect 494 384 506 436
rect 558 384 744 436
rect 796 384 808 436
rect 860 384 872 436
rect 924 384 931 436
rect 369 374 931 384
rect 369 45 415 374
rect 551 211 747 219
rect 551 159 560 211
rect 612 159 624 211
rect 676 159 688 211
rect 740 159 747 211
rect 551 149 747 159
rect 369 11 375 45
rect 409 11 415 45
rect 369 -27 415 11
rect 369 -61 375 -27
rect 409 -61 415 -27
rect 369 -108 415 -61
rect 627 45 673 149
rect 627 11 633 45
rect 667 11 673 45
rect 627 -27 673 11
rect 627 -61 633 -27
rect 667 -61 673 -27
rect 627 -108 673 -61
rect 885 45 931 374
rect 885 11 891 45
rect 925 11 931 45
rect 885 -27 931 11
rect 885 -61 891 -27
rect 925 -61 931 -27
rect 885 -108 931 -61
rect 1132 45 1178 490
rect 1315 310 1511 318
rect 1315 258 1324 310
rect 1376 258 1388 310
rect 1440 258 1452 310
rect 1504 258 1511 310
rect 1315 248 1511 258
rect 1132 11 1138 45
rect 1172 11 1178 45
rect 1132 -27 1178 11
rect 1132 -61 1138 -27
rect 1172 -61 1178 -27
rect 1132 -108 1178 -61
rect 1390 45 1436 248
rect 1390 11 1396 45
rect 1430 11 1436 45
rect 1390 -27 1436 11
rect 1390 -61 1396 -27
rect 1430 -61 1436 -27
rect 1390 -108 1436 -61
rect 1648 45 1694 490
rect 2917 488 3295 522
rect 3329 488 3707 522
rect 4853 552 5049 560
rect 4853 500 4860 552
rect 4912 500 4924 552
rect 4976 500 4988 552
rect 5040 500 5049 552
rect 4853 490 5049 500
rect 5370 552 5566 560
rect 5370 500 5377 552
rect 5429 500 5441 552
rect 5493 500 5505 552
rect 5557 500 5566 552
rect 5370 490 5566 500
rect 6456 522 6893 560
rect 2917 450 3707 488
rect 2153 436 2715 444
rect 2153 384 2162 436
rect 2214 384 2226 436
rect 2278 384 2290 436
rect 2342 384 2528 436
rect 2580 384 2592 436
rect 2644 384 2656 436
rect 2708 384 2715 436
rect 2153 374 2715 384
rect 1832 310 2028 318
rect 1832 258 1841 310
rect 1893 258 1905 310
rect 1957 258 1969 310
rect 2021 258 2028 310
rect 1832 248 2028 258
rect 1648 11 1654 45
rect 1688 11 1694 45
rect 1648 -27 1694 11
rect 1648 -61 1654 -27
rect 1688 -61 1694 -27
rect 1648 -108 1694 -61
rect 1906 45 1952 248
rect 1906 11 1912 45
rect 1946 11 1952 45
rect 1906 -27 1952 11
rect 1906 -61 1912 -27
rect 1946 -61 1952 -27
rect 1906 -108 1952 -61
rect 2153 45 2199 374
rect 2336 211 2532 219
rect 2336 159 2345 211
rect 2397 159 2409 211
rect 2461 159 2473 211
rect 2525 159 2532 211
rect 2336 149 2532 159
rect 2153 11 2159 45
rect 2193 11 2199 45
rect 2153 -27 2199 11
rect 2153 -61 2159 -27
rect 2193 -61 2199 -27
rect 2153 -108 2199 -61
rect 2411 45 2457 149
rect 2411 11 2417 45
rect 2451 11 2457 45
rect 2411 -27 2457 11
rect 2411 -61 2417 -27
rect 2451 -61 2457 -27
rect 2411 -108 2457 -61
rect 2669 45 2715 374
rect 2669 11 2675 45
rect 2709 11 2715 45
rect 2669 -27 2715 11
rect 2669 -61 2675 -27
rect 2709 -61 2715 -27
rect 2669 -108 2715 -61
rect 2917 416 3295 450
rect 3329 416 3707 450
rect 2917 378 3707 416
rect 2917 344 3295 378
rect 3329 344 3707 378
rect 2917 306 3707 344
rect 2917 272 3295 306
rect 3329 272 3707 306
rect 2917 234 3707 272
rect 2917 200 3295 234
rect 3329 200 3707 234
rect 2917 162 3707 200
rect 2917 128 3295 162
rect 3329 128 3707 162
rect 2917 90 3707 128
rect 2917 56 3295 90
rect 3329 56 3707 90
rect 2917 45 3707 56
rect 2917 11 2923 45
rect 2957 11 3181 45
rect 3215 18 3409 45
rect 3215 11 3295 18
rect 2917 -16 3295 11
rect 3329 11 3409 18
rect 3443 11 3667 45
rect 3701 11 3707 45
rect 3329 -16 3707 11
rect 2917 -27 3707 -16
rect 2917 -61 2923 -27
rect 2957 -61 3181 -27
rect 3215 -54 3409 -27
rect 3215 -61 3295 -54
rect 2917 -88 3295 -61
rect 3329 -61 3409 -54
rect 3443 -61 3667 -27
rect 3701 -61 3707 -27
rect 3329 -88 3707 -61
rect -269 -160 -244 -126
rect -210 -146 168 -126
rect 2917 -126 3707 -88
rect 3909 436 4471 444
rect 3909 384 3916 436
rect 3968 384 3980 436
rect 4032 384 4044 436
rect 4096 384 4282 436
rect 4334 384 4346 436
rect 4398 384 4410 436
rect 4462 384 4471 436
rect 3909 374 4471 384
rect 3909 45 3955 374
rect 4092 211 4288 219
rect 4092 159 4099 211
rect 4151 159 4163 211
rect 4215 159 4227 211
rect 4279 159 4288 211
rect 4092 149 4288 159
rect 3909 11 3915 45
rect 3949 11 3955 45
rect 3909 -27 3955 11
rect 3909 -61 3915 -27
rect 3949 -61 3955 -27
rect 3909 -108 3955 -61
rect 4167 45 4213 149
rect 4167 11 4173 45
rect 4207 11 4213 45
rect 4167 -27 4213 11
rect 4167 -61 4173 -27
rect 4207 -61 4213 -27
rect 4167 -108 4213 -61
rect 4425 45 4471 374
rect 4596 310 4792 318
rect 4596 258 4603 310
rect 4655 258 4667 310
rect 4719 258 4731 310
rect 4783 258 4792 310
rect 4596 248 4792 258
rect 4425 11 4431 45
rect 4465 11 4471 45
rect 4425 -27 4471 11
rect 4425 -61 4431 -27
rect 4465 -61 4471 -27
rect 4425 -108 4471 -61
rect 4672 45 4718 248
rect 4672 11 4678 45
rect 4712 11 4718 45
rect 4672 -27 4718 11
rect 4672 -61 4678 -27
rect 4712 -61 4718 -27
rect 4672 -108 4718 -61
rect 4930 45 4976 490
rect 5113 310 5309 318
rect 5113 258 5120 310
rect 5172 258 5184 310
rect 5236 258 5248 310
rect 5300 258 5309 310
rect 5113 248 5309 258
rect 4930 11 4936 45
rect 4970 11 4976 45
rect 4930 -27 4976 11
rect 4930 -61 4936 -27
rect 4970 -61 4976 -27
rect 4930 -108 4976 -61
rect 5188 45 5234 248
rect 5188 11 5194 45
rect 5228 11 5234 45
rect 5188 -27 5234 11
rect 5188 -61 5194 -27
rect 5228 -61 5234 -27
rect 5188 -108 5234 -61
rect 5446 45 5492 490
rect 6456 488 6834 522
rect 6868 488 6893 522
rect 6456 450 6893 488
rect 5446 11 5452 45
rect 5486 11 5492 45
rect 5446 -27 5492 11
rect 5446 -61 5452 -27
rect 5486 -61 5492 -27
rect 5446 -108 5492 -61
rect 5693 436 6255 444
rect 5693 384 5700 436
rect 5752 384 5764 436
rect 5816 384 5828 436
rect 5880 384 6066 436
rect 6118 384 6130 436
rect 6182 384 6194 436
rect 6246 384 6255 436
rect 5693 374 6255 384
rect 5693 45 5739 374
rect 5877 211 6073 219
rect 5877 159 5884 211
rect 5936 159 5948 211
rect 6000 159 6012 211
rect 6064 159 6073 211
rect 5877 149 6073 159
rect 5693 11 5699 45
rect 5733 11 5739 45
rect 5693 -27 5739 11
rect 5693 -61 5699 -27
rect 5733 -61 5739 -27
rect 5693 -108 5739 -61
rect 5951 45 5997 149
rect 5951 11 5957 45
rect 5991 11 5997 45
rect 5951 -27 5997 11
rect 5951 -61 5957 -27
rect 5991 -61 5997 -27
rect 5951 -108 5997 -61
rect 6209 45 6255 374
rect 6209 11 6215 45
rect 6249 11 6255 45
rect 6209 -27 6255 11
rect 6209 -61 6215 -27
rect 6249 -61 6255 -27
rect 6209 -108 6255 -61
rect 6456 416 6834 450
rect 6868 416 6893 450
rect 6456 378 6893 416
rect 6456 344 6834 378
rect 6868 344 6893 378
rect 6456 306 6893 344
rect 6456 272 6834 306
rect 6868 272 6893 306
rect 6456 234 6893 272
rect 6456 200 6834 234
rect 6868 200 6893 234
rect 6456 162 6893 200
rect 6456 128 6834 162
rect 6868 128 6893 162
rect 6456 90 6893 128
rect 6456 56 6834 90
rect 6868 56 6893 90
rect 6456 45 6893 56
rect 6456 11 6462 45
rect 6496 11 6720 45
rect 6754 18 6893 45
rect 6754 11 6834 18
rect 6456 -16 6834 11
rect 6868 -16 6893 18
rect 6456 -27 6893 -16
rect 6456 -61 6462 -27
rect 6496 -61 6720 -27
rect 6754 -54 6893 -27
rect 6754 -61 6834 -54
rect 6456 -88 6834 -61
rect 6868 -88 6893 -54
rect -210 -160 -37 -146
rect -269 -180 -37 -160
rect -3 -180 35 -146
rect 69 -180 168 -146
rect -269 -198 168 -180
rect -269 -232 -244 -198
rect -210 -232 168 -198
rect -269 -270 168 -232
rect -269 -304 -244 -270
rect -210 -304 168 -270
rect -269 -342 168 -304
rect -269 -376 -244 -342
rect -210 -376 168 -342
rect -269 -414 168 -376
rect 425 -146 875 -140
rect 425 -180 468 -146
rect 502 -180 540 -146
rect 574 -164 726 -146
rect 425 -216 551 -180
rect 603 -216 615 -164
rect 667 -216 679 -164
rect 760 -180 798 -146
rect 832 -180 875 -146
rect 731 -216 875 -180
rect 425 -315 875 -216
rect 425 -367 551 -315
rect 603 -367 615 -315
rect 667 -367 679 -315
rect 731 -367 875 -315
rect 425 -380 875 -367
rect 964 -146 2121 -140
rect 964 -180 1231 -146
rect 1265 -180 1303 -146
rect 1337 -180 1489 -146
rect 1523 -180 1561 -146
rect 1595 -180 1747 -146
rect 1781 -180 1819 -146
rect 1853 -180 2121 -146
rect 964 -236 2121 -180
rect -269 -448 -244 -414
rect -210 -448 168 -414
rect -269 -486 168 -448
rect 964 -453 1099 -236
rect -269 -520 -244 -486
rect -210 -509 168 -486
rect -210 -520 -37 -509
rect -269 -543 -37 -520
rect -3 -543 35 -509
rect 69 -543 168 -509
rect -269 -558 168 -543
rect 425 -473 1099 -453
rect 425 -509 551 -473
rect 425 -543 468 -509
rect 502 -543 540 -509
rect 603 -525 615 -473
rect 667 -525 679 -473
rect 731 -509 1099 -473
rect 574 -543 726 -525
rect 760 -543 798 -509
rect 832 -543 1099 -509
rect 425 -549 1099 -543
rect 1188 -315 1896 -299
rect 1188 -367 1217 -315
rect 1269 -367 1281 -315
rect 1333 -367 1345 -315
rect 1397 -367 1446 -315
rect 1498 -367 1510 -315
rect 1562 -367 1574 -315
rect 1626 -367 1684 -315
rect 1736 -367 1748 -315
rect 1800 -367 1812 -315
rect 1864 -367 1896 -315
rect 1188 -509 1896 -367
rect 1188 -543 1231 -509
rect 1265 -543 1303 -509
rect 1337 -543 1489 -509
rect 1523 -543 1561 -509
rect 1595 -543 1747 -509
rect 1781 -543 1819 -509
rect 1853 -543 1896 -509
rect 1188 -549 1896 -543
rect 1988 -453 2121 -236
rect 2209 -146 2659 -140
rect 2209 -180 2252 -146
rect 2286 -180 2324 -146
rect 2358 -164 2510 -146
rect 2209 -216 2335 -180
rect 2387 -216 2399 -164
rect 2451 -216 2463 -164
rect 2544 -180 2582 -146
rect 2616 -180 2659 -146
rect 2515 -216 2659 -180
rect 2209 -315 2659 -216
rect 2209 -367 2335 -315
rect 2387 -367 2399 -315
rect 2451 -367 2463 -315
rect 2515 -367 2659 -315
rect 2209 -380 2659 -367
rect 2917 -146 3295 -126
rect 2917 -180 3016 -146
rect 3050 -180 3088 -146
rect 3122 -160 3295 -146
rect 3329 -146 3707 -126
rect 6456 -126 6893 -88
rect 3329 -160 3502 -146
rect 3122 -180 3502 -160
rect 3536 -180 3574 -146
rect 3608 -180 3707 -146
rect 2917 -198 3707 -180
rect 2917 -232 3295 -198
rect 3329 -232 3707 -198
rect 2917 -270 3707 -232
rect 2917 -304 3295 -270
rect 3329 -304 3707 -270
rect 2917 -342 3707 -304
rect 2917 -376 3295 -342
rect 3329 -376 3707 -342
rect 2917 -414 3707 -376
rect 3965 -146 4415 -140
rect 3965 -180 4008 -146
rect 4042 -180 4080 -146
rect 4114 -164 4266 -146
rect 3965 -216 4109 -180
rect 4161 -216 4173 -164
rect 4225 -216 4237 -164
rect 4300 -180 4338 -146
rect 4372 -180 4415 -146
rect 4289 -216 4415 -180
rect 3965 -315 4415 -216
rect 3965 -367 4109 -315
rect 4161 -367 4173 -315
rect 4225 -367 4237 -315
rect 4289 -367 4415 -315
rect 3965 -380 4415 -367
rect 4503 -146 5660 -140
rect 4503 -180 4771 -146
rect 4805 -180 4843 -146
rect 4877 -180 5029 -146
rect 5063 -180 5101 -146
rect 5135 -180 5287 -146
rect 5321 -180 5359 -146
rect 5393 -180 5660 -146
rect 4503 -236 5660 -180
rect 2917 -448 3295 -414
rect 3329 -448 3707 -414
rect 1988 -473 2659 -453
rect 1988 -509 2335 -473
rect 1988 -543 2252 -509
rect 2286 -543 2324 -509
rect 2387 -525 2399 -473
rect 2451 -525 2463 -473
rect 2515 -509 2659 -473
rect 2358 -543 2510 -525
rect 2544 -543 2582 -509
rect 2616 -543 2659 -509
rect 1988 -549 2659 -543
rect 2917 -486 3707 -448
rect 4503 -453 4636 -236
rect 2917 -509 3295 -486
rect 2917 -543 3016 -509
rect 3050 -543 3088 -509
rect 3122 -520 3295 -509
rect 3329 -509 3707 -486
rect 3329 -520 3502 -509
rect 3122 -543 3502 -520
rect 3536 -543 3574 -509
rect 3608 -543 3707 -509
rect -269 -592 -244 -558
rect -210 -592 168 -558
rect 2917 -558 3707 -543
rect 3965 -473 4636 -453
rect 3965 -509 4109 -473
rect 3965 -543 4008 -509
rect 4042 -543 4080 -509
rect 4161 -525 4173 -473
rect 4225 -525 4237 -473
rect 4289 -509 4636 -473
rect 4114 -543 4266 -525
rect 4300 -543 4338 -509
rect 4372 -543 4636 -509
rect 3965 -549 4636 -543
rect 4728 -315 5436 -299
rect 4728 -367 4760 -315
rect 4812 -367 4824 -315
rect 4876 -367 4888 -315
rect 4940 -367 4998 -315
rect 5050 -367 5062 -315
rect 5114 -367 5126 -315
rect 5178 -367 5227 -315
rect 5279 -367 5291 -315
rect 5343 -367 5355 -315
rect 5407 -367 5436 -315
rect 4728 -509 5436 -367
rect 4728 -543 4771 -509
rect 4805 -543 4843 -509
rect 4877 -543 5029 -509
rect 5063 -543 5101 -509
rect 5135 -543 5287 -509
rect 5321 -543 5359 -509
rect 5393 -543 5436 -509
rect 4728 -549 5436 -543
rect 5525 -453 5660 -236
rect 5749 -146 6199 -140
rect 5749 -180 5792 -146
rect 5826 -180 5864 -146
rect 5898 -164 6050 -146
rect 5749 -216 5893 -180
rect 5945 -216 5957 -164
rect 6009 -216 6021 -164
rect 6084 -180 6122 -146
rect 6156 -180 6199 -146
rect 6073 -216 6199 -180
rect 5749 -315 6199 -216
rect 5749 -367 5893 -315
rect 5945 -367 5957 -315
rect 6009 -367 6021 -315
rect 6073 -367 6199 -315
rect 5749 -380 6199 -367
rect 6456 -146 6834 -126
rect 6456 -180 6555 -146
rect 6589 -180 6627 -146
rect 6661 -160 6834 -146
rect 6868 -160 6893 -126
rect 6661 -180 6893 -160
rect 6456 -198 6893 -180
rect 6456 -232 6834 -198
rect 6868 -232 6893 -198
rect 6456 -270 6893 -232
rect 6456 -304 6834 -270
rect 6868 -304 6893 -270
rect 6456 -342 6893 -304
rect 6456 -376 6834 -342
rect 6868 -376 6893 -342
rect 6456 -414 6893 -376
rect 6456 -448 6834 -414
rect 6868 -448 6893 -414
rect 5525 -473 6199 -453
rect 5525 -509 5893 -473
rect 5525 -543 5792 -509
rect 5826 -543 5864 -509
rect 5945 -525 5957 -473
rect 6009 -525 6021 -473
rect 6073 -509 6199 -473
rect 5898 -543 6050 -525
rect 6084 -543 6122 -509
rect 6156 -543 6199 -509
rect 5525 -549 6199 -543
rect 6456 -486 6893 -448
rect 6456 -509 6834 -486
rect 6456 -543 6555 -509
rect 6589 -543 6627 -509
rect 6661 -520 6834 -509
rect 6868 -520 6893 -486
rect 6661 -543 6893 -520
rect -269 -628 168 -592
rect -269 -630 -130 -628
rect -269 -664 -244 -630
rect -210 -662 -130 -630
rect -96 -662 128 -628
rect 162 -662 168 -628
rect -210 -664 168 -662
rect -269 -700 168 -664
rect -269 -702 -130 -700
rect -269 -736 -244 -702
rect -210 -734 -130 -702
rect -96 -734 128 -700
rect 162 -734 168 -700
rect -210 -736 168 -734
rect -269 -774 168 -736
rect -269 -808 -244 -774
rect -210 -808 168 -774
rect -269 -846 168 -808
rect -269 -880 -244 -846
rect -210 -880 168 -846
rect -269 -918 168 -880
rect -269 -952 -244 -918
rect -210 -952 168 -918
rect -269 -990 168 -952
rect -269 -1024 -244 -990
rect -210 -1024 168 -990
rect -269 -1062 168 -1024
rect -269 -1096 -244 -1062
rect -210 -1096 168 -1062
rect 369 -628 415 -581
rect 369 -662 375 -628
rect 409 -662 415 -628
rect 369 -700 415 -662
rect 369 -734 375 -700
rect 409 -734 415 -700
rect 369 -1063 415 -734
rect 627 -628 673 -581
rect 627 -662 633 -628
rect 667 -662 673 -628
rect 627 -700 673 -662
rect 627 -734 633 -700
rect 667 -734 673 -700
rect 627 -799 673 -734
rect 885 -628 931 -581
rect 885 -662 891 -628
rect 925 -662 931 -628
rect 885 -700 931 -662
rect 885 -734 891 -700
rect 925 -734 931 -700
rect 553 -809 749 -799
rect 553 -861 560 -809
rect 612 -861 624 -809
rect 676 -861 688 -809
rect 740 -861 749 -809
rect 553 -869 749 -861
rect -269 -1134 168 -1096
rect 294 -1073 490 -1063
rect 294 -1125 301 -1073
rect 353 -1125 365 -1073
rect 417 -1125 429 -1073
rect 481 -1125 490 -1073
rect 294 -1133 490 -1125
rect -269 -1168 -244 -1134
rect -210 -1168 168 -1134
rect -269 -1206 168 -1168
rect -269 -1240 -244 -1206
rect -210 -1240 168 -1206
rect -269 -1278 168 -1240
rect -269 -1312 -244 -1278
rect -210 -1312 168 -1278
rect -269 -1350 168 -1312
rect -269 -1384 -244 -1350
rect -210 -1352 168 -1350
rect -210 -1384 -130 -1352
rect -269 -1386 -130 -1384
rect -96 -1386 128 -1352
rect 162 -1386 168 -1352
rect -269 -1422 168 -1386
rect -269 -1456 -244 -1422
rect -210 -1424 168 -1422
rect -210 -1456 -130 -1424
rect -269 -1458 -130 -1456
rect -96 -1458 128 -1424
rect 162 -1458 168 -1424
rect -269 -1494 168 -1458
rect -269 -1528 -244 -1494
rect -210 -1528 168 -1494
rect 369 -1352 415 -1133
rect 369 -1386 375 -1352
rect 409 -1386 415 -1352
rect 369 -1424 415 -1386
rect 369 -1458 375 -1424
rect 409 -1458 415 -1424
rect 369 -1505 415 -1458
rect 627 -1352 673 -869
rect 885 -1063 931 -734
rect 1132 -628 1178 -581
rect 1132 -662 1138 -628
rect 1172 -662 1178 -628
rect 1132 -700 1178 -662
rect 1132 -734 1138 -700
rect 1172 -734 1178 -700
rect 1132 -952 1178 -734
rect 1390 -628 1436 -581
rect 1390 -662 1396 -628
rect 1430 -662 1436 -628
rect 1390 -700 1436 -662
rect 1390 -734 1396 -700
rect 1430 -734 1436 -700
rect 1057 -962 1253 -952
rect 1057 -1014 1064 -962
rect 1116 -1014 1128 -962
rect 1180 -1014 1192 -962
rect 1244 -1014 1253 -962
rect 1057 -1022 1253 -1014
rect 813 -1073 1009 -1063
rect 813 -1125 820 -1073
rect 872 -1125 884 -1073
rect 936 -1125 948 -1073
rect 1000 -1125 1009 -1073
rect 813 -1133 1009 -1125
rect 627 -1386 633 -1352
rect 667 -1386 673 -1352
rect 627 -1424 673 -1386
rect 627 -1458 633 -1424
rect 667 -1458 673 -1424
rect 627 -1505 673 -1458
rect 885 -1352 931 -1133
rect 885 -1386 891 -1352
rect 925 -1386 931 -1352
rect 885 -1424 931 -1386
rect 885 -1458 891 -1424
rect 925 -1458 931 -1424
rect 885 -1505 931 -1458
rect 1132 -1352 1178 -1022
rect 1390 -1163 1436 -734
rect 1648 -628 1694 -581
rect 1648 -662 1654 -628
rect 1688 -662 1694 -628
rect 1648 -700 1694 -662
rect 1648 -734 1654 -700
rect 1688 -734 1694 -700
rect 1648 -952 1694 -734
rect 1906 -628 1952 -581
rect 1906 -662 1912 -628
rect 1946 -662 1952 -628
rect 1906 -700 1952 -662
rect 1906 -734 1912 -700
rect 1946 -734 1952 -700
rect 1574 -962 1770 -952
rect 1574 -1014 1581 -962
rect 1633 -1014 1645 -962
rect 1697 -1014 1709 -962
rect 1761 -1014 1770 -962
rect 1574 -1022 1770 -1014
rect 1314 -1173 1510 -1163
rect 1314 -1225 1321 -1173
rect 1373 -1225 1385 -1173
rect 1437 -1225 1449 -1173
rect 1501 -1225 1510 -1173
rect 1314 -1233 1510 -1225
rect 1132 -1386 1138 -1352
rect 1172 -1386 1178 -1352
rect 1132 -1424 1178 -1386
rect 1132 -1458 1138 -1424
rect 1172 -1458 1178 -1424
rect 1132 -1505 1178 -1458
rect 1390 -1352 1436 -1233
rect 1390 -1386 1396 -1352
rect 1430 -1386 1436 -1352
rect 1390 -1424 1436 -1386
rect 1390 -1458 1396 -1424
rect 1430 -1458 1436 -1424
rect 1390 -1505 1436 -1458
rect 1648 -1352 1694 -1022
rect 1906 -1163 1952 -734
rect 2153 -628 2199 -581
rect 2153 -662 2159 -628
rect 2193 -662 2199 -628
rect 2153 -700 2199 -662
rect 2153 -734 2159 -700
rect 2193 -734 2199 -700
rect 2153 -1063 2199 -734
rect 2411 -628 2457 -581
rect 2411 -662 2417 -628
rect 2451 -662 2457 -628
rect 2411 -700 2457 -662
rect 2411 -734 2417 -700
rect 2451 -734 2457 -700
rect 2411 -799 2457 -734
rect 2669 -628 2715 -581
rect 2669 -662 2675 -628
rect 2709 -662 2715 -628
rect 2669 -700 2715 -662
rect 2669 -734 2675 -700
rect 2709 -734 2715 -700
rect 2337 -809 2533 -799
rect 2337 -861 2344 -809
rect 2396 -861 2408 -809
rect 2460 -861 2472 -809
rect 2524 -861 2533 -809
rect 2337 -869 2533 -861
rect 2080 -1073 2276 -1063
rect 2080 -1125 2087 -1073
rect 2139 -1125 2151 -1073
rect 2203 -1125 2215 -1073
rect 2267 -1125 2276 -1073
rect 2080 -1133 2276 -1125
rect 1831 -1173 2027 -1163
rect 1831 -1225 1838 -1173
rect 1890 -1225 1902 -1173
rect 1954 -1225 1966 -1173
rect 2018 -1225 2027 -1173
rect 1831 -1233 2027 -1225
rect 1648 -1386 1654 -1352
rect 1688 -1386 1694 -1352
rect 1648 -1424 1694 -1386
rect 1648 -1458 1654 -1424
rect 1688 -1458 1694 -1424
rect 1648 -1505 1694 -1458
rect 1906 -1352 1952 -1233
rect 1906 -1386 1912 -1352
rect 1946 -1386 1952 -1352
rect 1906 -1424 1952 -1386
rect 1906 -1458 1912 -1424
rect 1946 -1458 1952 -1424
rect 1906 -1505 1952 -1458
rect 2153 -1352 2199 -1133
rect 2153 -1386 2159 -1352
rect 2193 -1386 2199 -1352
rect 2153 -1424 2199 -1386
rect 2153 -1458 2159 -1424
rect 2193 -1458 2199 -1424
rect 2153 -1505 2199 -1458
rect 2411 -1352 2457 -869
rect 2669 -1063 2715 -734
rect 2917 -592 3295 -558
rect 3329 -592 3707 -558
rect 6456 -558 6893 -543
rect 2917 -628 3707 -592
rect 2917 -662 2923 -628
rect 2957 -662 3181 -628
rect 3215 -630 3409 -628
rect 3215 -662 3295 -630
rect 2917 -664 3295 -662
rect 3329 -662 3409 -630
rect 3443 -662 3667 -628
rect 3701 -662 3707 -628
rect 3329 -664 3707 -662
rect 2917 -700 3707 -664
rect 2917 -734 2923 -700
rect 2957 -734 3181 -700
rect 3215 -702 3409 -700
rect 3215 -734 3295 -702
rect 2917 -736 3295 -734
rect 3329 -734 3409 -702
rect 3443 -734 3667 -700
rect 3701 -734 3707 -700
rect 3329 -736 3707 -734
rect 2917 -774 3707 -736
rect 2917 -808 3295 -774
rect 3329 -808 3707 -774
rect 2917 -846 3707 -808
rect 2917 -880 3295 -846
rect 3329 -880 3707 -846
rect 2917 -918 3707 -880
rect 2917 -952 3295 -918
rect 3329 -952 3707 -918
rect 2917 -990 3707 -952
rect 2917 -1024 3295 -990
rect 3329 -1024 3707 -990
rect 2917 -1062 3707 -1024
rect 2597 -1073 2793 -1063
rect 2597 -1125 2604 -1073
rect 2656 -1125 2668 -1073
rect 2720 -1125 2732 -1073
rect 2784 -1125 2793 -1073
rect 2597 -1133 2793 -1125
rect 2917 -1096 3295 -1062
rect 3329 -1096 3707 -1062
rect 3909 -628 3955 -581
rect 3909 -662 3915 -628
rect 3949 -662 3955 -628
rect 3909 -700 3955 -662
rect 3909 -734 3915 -700
rect 3949 -734 3955 -700
rect 3909 -1063 3955 -734
rect 4167 -628 4213 -581
rect 4167 -662 4173 -628
rect 4207 -662 4213 -628
rect 4167 -700 4213 -662
rect 4167 -734 4173 -700
rect 4207 -734 4213 -700
rect 4167 -799 4213 -734
rect 4425 -628 4471 -581
rect 4425 -662 4431 -628
rect 4465 -662 4471 -628
rect 4425 -700 4471 -662
rect 4425 -734 4431 -700
rect 4465 -734 4471 -700
rect 4091 -809 4287 -799
rect 4091 -861 4100 -809
rect 4152 -861 4164 -809
rect 4216 -861 4228 -809
rect 4280 -861 4287 -809
rect 4091 -869 4287 -861
rect 2411 -1386 2417 -1352
rect 2451 -1386 2457 -1352
rect 2411 -1424 2457 -1386
rect 2411 -1458 2417 -1424
rect 2451 -1458 2457 -1424
rect 2411 -1505 2457 -1458
rect 2669 -1352 2715 -1133
rect 2669 -1386 2675 -1352
rect 2709 -1386 2715 -1352
rect 2669 -1424 2715 -1386
rect 2669 -1458 2675 -1424
rect 2709 -1458 2715 -1424
rect 2669 -1505 2715 -1458
rect 2917 -1134 3707 -1096
rect 3831 -1073 4027 -1063
rect 3831 -1125 3840 -1073
rect 3892 -1125 3904 -1073
rect 3956 -1125 3968 -1073
rect 4020 -1125 4027 -1073
rect 3831 -1133 4027 -1125
rect 2917 -1168 3295 -1134
rect 3329 -1168 3707 -1134
rect 2917 -1206 3707 -1168
rect 2917 -1240 3295 -1206
rect 3329 -1240 3707 -1206
rect 2917 -1278 3707 -1240
rect 2917 -1312 3295 -1278
rect 3329 -1312 3707 -1278
rect 2917 -1350 3707 -1312
rect 2917 -1352 3295 -1350
rect 2917 -1386 2923 -1352
rect 2957 -1386 3181 -1352
rect 3215 -1384 3295 -1352
rect 3329 -1352 3707 -1350
rect 3329 -1384 3409 -1352
rect 3215 -1386 3409 -1384
rect 3443 -1386 3667 -1352
rect 3701 -1386 3707 -1352
rect 2917 -1422 3707 -1386
rect 2917 -1424 3295 -1422
rect 2917 -1458 2923 -1424
rect 2957 -1458 3181 -1424
rect 3215 -1456 3295 -1424
rect 3329 -1424 3707 -1422
rect 3329 -1456 3409 -1424
rect 3215 -1458 3409 -1456
rect 3443 -1458 3667 -1424
rect 3701 -1458 3707 -1424
rect 2917 -1494 3707 -1458
rect -269 -1543 168 -1528
rect 2917 -1528 3295 -1494
rect 3329 -1528 3707 -1494
rect 3909 -1352 3955 -1133
rect 3909 -1386 3915 -1352
rect 3949 -1386 3955 -1352
rect 3909 -1424 3955 -1386
rect 3909 -1458 3915 -1424
rect 3949 -1458 3955 -1424
rect 3909 -1505 3955 -1458
rect 4167 -1352 4213 -869
rect 4425 -1063 4471 -734
rect 4672 -628 4718 -581
rect 4672 -662 4678 -628
rect 4712 -662 4718 -628
rect 4672 -700 4718 -662
rect 4672 -734 4678 -700
rect 4712 -734 4718 -700
rect 4348 -1073 4544 -1063
rect 4348 -1125 4357 -1073
rect 4409 -1125 4421 -1073
rect 4473 -1125 4485 -1073
rect 4537 -1125 4544 -1073
rect 4348 -1133 4544 -1125
rect 4167 -1386 4173 -1352
rect 4207 -1386 4213 -1352
rect 4167 -1424 4213 -1386
rect 4167 -1458 4173 -1424
rect 4207 -1458 4213 -1424
rect 4167 -1505 4213 -1458
rect 4425 -1352 4471 -1133
rect 4672 -1163 4718 -734
rect 4930 -628 4976 -581
rect 4930 -662 4936 -628
rect 4970 -662 4976 -628
rect 4930 -700 4976 -662
rect 4930 -734 4936 -700
rect 4970 -734 4976 -700
rect 4930 -952 4976 -734
rect 5188 -628 5234 -581
rect 5188 -662 5194 -628
rect 5228 -662 5234 -628
rect 5188 -700 5234 -662
rect 5188 -734 5194 -700
rect 5228 -734 5234 -700
rect 4854 -962 5050 -952
rect 4854 -1014 4863 -962
rect 4915 -1014 4927 -962
rect 4979 -1014 4991 -962
rect 5043 -1014 5050 -962
rect 4854 -1022 5050 -1014
rect 4597 -1173 4793 -1163
rect 4597 -1225 4606 -1173
rect 4658 -1225 4670 -1173
rect 4722 -1225 4734 -1173
rect 4786 -1225 4793 -1173
rect 4597 -1233 4793 -1225
rect 4425 -1386 4431 -1352
rect 4465 -1386 4471 -1352
rect 4425 -1424 4471 -1386
rect 4425 -1458 4431 -1424
rect 4465 -1458 4471 -1424
rect 4425 -1505 4471 -1458
rect 4672 -1352 4718 -1233
rect 4672 -1386 4678 -1352
rect 4712 -1386 4718 -1352
rect 4672 -1424 4718 -1386
rect 4672 -1458 4678 -1424
rect 4712 -1458 4718 -1424
rect 4672 -1505 4718 -1458
rect 4930 -1352 4976 -1022
rect 5188 -1163 5234 -734
rect 5446 -628 5492 -581
rect 5446 -662 5452 -628
rect 5486 -662 5492 -628
rect 5446 -700 5492 -662
rect 5446 -734 5452 -700
rect 5486 -734 5492 -700
rect 5446 -952 5492 -734
rect 5693 -628 5739 -581
rect 5693 -662 5699 -628
rect 5733 -662 5739 -628
rect 5693 -700 5739 -662
rect 5693 -734 5699 -700
rect 5733 -734 5739 -700
rect 5371 -962 5567 -952
rect 5371 -1014 5380 -962
rect 5432 -1014 5444 -962
rect 5496 -1014 5508 -962
rect 5560 -1014 5567 -962
rect 5371 -1022 5567 -1014
rect 5114 -1173 5310 -1163
rect 5114 -1225 5123 -1173
rect 5175 -1225 5187 -1173
rect 5239 -1225 5251 -1173
rect 5303 -1225 5310 -1173
rect 5114 -1233 5310 -1225
rect 4930 -1386 4936 -1352
rect 4970 -1386 4976 -1352
rect 4930 -1424 4976 -1386
rect 4930 -1458 4936 -1424
rect 4970 -1458 4976 -1424
rect 4930 -1505 4976 -1458
rect 5188 -1352 5234 -1233
rect 5188 -1386 5194 -1352
rect 5228 -1386 5234 -1352
rect 5188 -1424 5234 -1386
rect 5188 -1458 5194 -1424
rect 5228 -1458 5234 -1424
rect 5188 -1505 5234 -1458
rect 5446 -1352 5492 -1022
rect 5693 -1063 5739 -734
rect 5951 -628 5997 -581
rect 5951 -662 5957 -628
rect 5991 -662 5997 -628
rect 5951 -700 5997 -662
rect 5951 -734 5957 -700
rect 5991 -734 5997 -700
rect 5951 -799 5997 -734
rect 6209 -628 6255 -581
rect 6209 -662 6215 -628
rect 6249 -662 6255 -628
rect 6209 -700 6255 -662
rect 6209 -734 6215 -700
rect 6249 -734 6255 -700
rect 5875 -809 6071 -799
rect 5875 -861 5884 -809
rect 5936 -861 5948 -809
rect 6000 -861 6012 -809
rect 6064 -861 6071 -809
rect 5875 -869 6071 -861
rect 5615 -1073 5811 -1063
rect 5615 -1125 5624 -1073
rect 5676 -1125 5688 -1073
rect 5740 -1125 5752 -1073
rect 5804 -1125 5811 -1073
rect 5615 -1133 5811 -1125
rect 5446 -1386 5452 -1352
rect 5486 -1386 5492 -1352
rect 5446 -1424 5492 -1386
rect 5446 -1458 5452 -1424
rect 5486 -1458 5492 -1424
rect 5446 -1505 5492 -1458
rect 5693 -1352 5739 -1133
rect 5693 -1386 5699 -1352
rect 5733 -1386 5739 -1352
rect 5693 -1424 5739 -1386
rect 5693 -1458 5699 -1424
rect 5733 -1458 5739 -1424
rect 5693 -1505 5739 -1458
rect 5951 -1352 5997 -869
rect 6209 -1063 6255 -734
rect 6456 -592 6834 -558
rect 6868 -592 6893 -558
rect 6456 -628 6893 -592
rect 6456 -662 6462 -628
rect 6496 -662 6720 -628
rect 6754 -630 6893 -628
rect 6754 -662 6834 -630
rect 6456 -664 6834 -662
rect 6868 -664 6893 -630
rect 6456 -700 6893 -664
rect 6456 -734 6462 -700
rect 6496 -734 6720 -700
rect 6754 -702 6893 -700
rect 6754 -734 6834 -702
rect 6456 -736 6834 -734
rect 6868 -736 6893 -702
rect 6456 -774 6893 -736
rect 6456 -808 6834 -774
rect 6868 -808 6893 -774
rect 6456 -846 6893 -808
rect 6456 -880 6834 -846
rect 6868 -880 6893 -846
rect 6456 -918 6893 -880
rect 6456 -952 6834 -918
rect 6868 -952 6893 -918
rect 6456 -990 6893 -952
rect 6456 -1024 6834 -990
rect 6868 -1024 6893 -990
rect 6456 -1062 6893 -1024
rect 6134 -1073 6330 -1063
rect 6134 -1125 6143 -1073
rect 6195 -1125 6207 -1073
rect 6259 -1125 6271 -1073
rect 6323 -1125 6330 -1073
rect 6134 -1133 6330 -1125
rect 6456 -1096 6834 -1062
rect 6868 -1096 6893 -1062
rect 5951 -1386 5957 -1352
rect 5991 -1386 5997 -1352
rect 5951 -1424 5997 -1386
rect 5951 -1458 5957 -1424
rect 5991 -1458 5997 -1424
rect 5951 -1505 5997 -1458
rect 6209 -1352 6255 -1133
rect 6209 -1386 6215 -1352
rect 6249 -1386 6255 -1352
rect 6209 -1424 6255 -1386
rect 6209 -1458 6215 -1424
rect 6249 -1458 6255 -1424
rect 6209 -1505 6255 -1458
rect 6456 -1134 6893 -1096
rect 6456 -1168 6834 -1134
rect 6868 -1168 6893 -1134
rect 6456 -1206 6893 -1168
rect 6456 -1240 6834 -1206
rect 6868 -1240 6893 -1206
rect 6456 -1278 6893 -1240
rect 6456 -1312 6834 -1278
rect 6868 -1312 6893 -1278
rect 6456 -1350 6893 -1312
rect 6456 -1352 6834 -1350
rect 6456 -1386 6462 -1352
rect 6496 -1386 6720 -1352
rect 6754 -1384 6834 -1352
rect 6868 -1384 6893 -1350
rect 6754 -1386 6893 -1384
rect 6456 -1422 6893 -1386
rect 6456 -1424 6834 -1422
rect 6456 -1458 6462 -1424
rect 6496 -1458 6720 -1424
rect 6754 -1456 6834 -1424
rect 6868 -1456 6893 -1422
rect 6754 -1458 6893 -1456
rect 6456 -1494 6893 -1458
rect -269 -1566 -37 -1543
rect -269 -1600 -244 -1566
rect -210 -1577 -37 -1566
rect -3 -1577 35 -1543
rect 69 -1577 168 -1543
rect -210 -1600 168 -1577
rect -269 -1638 168 -1600
rect 425 -1543 1099 -1537
rect 425 -1577 468 -1543
rect 502 -1577 540 -1543
rect 574 -1561 726 -1543
rect 425 -1613 551 -1577
rect 603 -1613 615 -1561
rect 667 -1613 679 -1561
rect 760 -1577 798 -1543
rect 832 -1577 1099 -1543
rect 731 -1613 1099 -1577
rect 425 -1633 1099 -1613
rect -269 -1672 -244 -1638
rect -210 -1672 168 -1638
rect -269 -1710 168 -1672
rect -269 -1744 -244 -1710
rect -210 -1744 168 -1710
rect -269 -1782 168 -1744
rect -269 -1816 -244 -1782
rect -210 -1816 168 -1782
rect -269 -1854 168 -1816
rect -269 -1888 -244 -1854
rect -210 -1888 168 -1854
rect -269 -1906 168 -1888
rect -269 -1926 -37 -1906
rect -269 -1960 -244 -1926
rect -210 -1940 -37 -1926
rect -3 -1940 35 -1906
rect 69 -1940 168 -1906
rect -210 -1960 168 -1940
rect 425 -1718 875 -1706
rect 425 -1770 551 -1718
rect 603 -1770 615 -1718
rect 667 -1770 679 -1718
rect 731 -1770 875 -1718
rect 425 -1870 875 -1770
rect 425 -1906 551 -1870
rect 425 -1940 468 -1906
rect 502 -1940 540 -1906
rect 603 -1922 615 -1870
rect 667 -1922 679 -1870
rect 731 -1906 875 -1870
rect 574 -1940 726 -1922
rect 760 -1940 798 -1906
rect 832 -1940 875 -1906
rect 425 -1946 875 -1940
rect 964 -1850 1099 -1633
rect 1188 -1543 1896 -1537
rect 1188 -1577 1231 -1543
rect 1265 -1577 1303 -1543
rect 1337 -1577 1489 -1543
rect 1523 -1577 1561 -1543
rect 1595 -1577 1747 -1543
rect 1781 -1577 1819 -1543
rect 1853 -1577 1896 -1543
rect 1188 -1718 1896 -1577
rect 1188 -1770 1217 -1718
rect 1269 -1770 1281 -1718
rect 1333 -1770 1345 -1718
rect 1397 -1770 1446 -1718
rect 1498 -1770 1510 -1718
rect 1562 -1770 1574 -1718
rect 1626 -1770 1684 -1718
rect 1736 -1770 1748 -1718
rect 1800 -1770 1812 -1718
rect 1864 -1770 1896 -1718
rect 1188 -1787 1896 -1770
rect 1988 -1543 2659 -1537
rect 1988 -1577 2252 -1543
rect 2286 -1577 2324 -1543
rect 2358 -1561 2510 -1543
rect 1988 -1613 2335 -1577
rect 2387 -1613 2399 -1561
rect 2451 -1613 2463 -1561
rect 2544 -1577 2582 -1543
rect 2616 -1577 2659 -1543
rect 2515 -1613 2659 -1577
rect 1988 -1633 2659 -1613
rect 2917 -1543 3707 -1528
rect 6456 -1528 6834 -1494
rect 6868 -1528 6893 -1494
rect 2917 -1577 3016 -1543
rect 3050 -1577 3088 -1543
rect 3122 -1566 3502 -1543
rect 3122 -1577 3295 -1566
rect 2917 -1600 3295 -1577
rect 3329 -1577 3502 -1566
rect 3536 -1577 3574 -1543
rect 3608 -1577 3707 -1543
rect 3329 -1600 3707 -1577
rect 1988 -1850 2121 -1633
rect 2917 -1638 3707 -1600
rect 3965 -1543 4636 -1537
rect 3965 -1577 4008 -1543
rect 4042 -1577 4080 -1543
rect 4114 -1561 4266 -1543
rect 3965 -1613 4109 -1577
rect 4161 -1613 4173 -1561
rect 4225 -1613 4237 -1561
rect 4300 -1577 4338 -1543
rect 4372 -1577 4636 -1543
rect 4289 -1613 4636 -1577
rect 3965 -1633 4636 -1613
rect 2917 -1672 3295 -1638
rect 3329 -1672 3707 -1638
rect 964 -1906 2121 -1850
rect 964 -1940 1231 -1906
rect 1265 -1940 1303 -1906
rect 1337 -1940 1489 -1906
rect 1523 -1940 1561 -1906
rect 1595 -1940 1747 -1906
rect 1781 -1940 1819 -1906
rect 1853 -1940 2121 -1906
rect 964 -1946 2121 -1940
rect 2209 -1718 2659 -1706
rect 2209 -1770 2335 -1718
rect 2387 -1770 2399 -1718
rect 2451 -1770 2463 -1718
rect 2515 -1770 2659 -1718
rect 2209 -1870 2659 -1770
rect 2209 -1906 2335 -1870
rect 2209 -1940 2252 -1906
rect 2286 -1940 2324 -1906
rect 2387 -1922 2399 -1870
rect 2451 -1922 2463 -1870
rect 2515 -1906 2659 -1870
rect 2358 -1940 2510 -1922
rect 2544 -1940 2582 -1906
rect 2616 -1940 2659 -1906
rect 2209 -1946 2659 -1940
rect 2917 -1710 3707 -1672
rect 2917 -1744 3295 -1710
rect 3329 -1744 3707 -1710
rect 2917 -1782 3707 -1744
rect 2917 -1816 3295 -1782
rect 3329 -1816 3707 -1782
rect 2917 -1854 3707 -1816
rect 2917 -1888 3295 -1854
rect 3329 -1888 3707 -1854
rect 2917 -1906 3707 -1888
rect 2917 -1940 3016 -1906
rect 3050 -1940 3088 -1906
rect 3122 -1926 3502 -1906
rect 3122 -1940 3295 -1926
rect -269 -1998 168 -1960
rect 2917 -1960 3295 -1940
rect 3329 -1940 3502 -1926
rect 3536 -1940 3574 -1906
rect 3608 -1940 3707 -1906
rect 3329 -1960 3707 -1940
rect 3965 -1718 4415 -1706
rect 3965 -1770 4109 -1718
rect 4161 -1770 4173 -1718
rect 4225 -1770 4237 -1718
rect 4289 -1770 4415 -1718
rect 3965 -1870 4415 -1770
rect 3965 -1906 4109 -1870
rect 3965 -1940 4008 -1906
rect 4042 -1940 4080 -1906
rect 4161 -1922 4173 -1870
rect 4225 -1922 4237 -1870
rect 4289 -1906 4415 -1870
rect 4114 -1940 4266 -1922
rect 4300 -1940 4338 -1906
rect 4372 -1940 4415 -1906
rect 3965 -1946 4415 -1940
rect 4503 -1850 4636 -1633
rect 4728 -1543 5436 -1537
rect 4728 -1577 4771 -1543
rect 4805 -1577 4843 -1543
rect 4877 -1577 5029 -1543
rect 5063 -1577 5101 -1543
rect 5135 -1577 5287 -1543
rect 5321 -1577 5359 -1543
rect 5393 -1577 5436 -1543
rect 4728 -1718 5436 -1577
rect 4728 -1770 4760 -1718
rect 4812 -1770 4824 -1718
rect 4876 -1770 4888 -1718
rect 4940 -1770 4998 -1718
rect 5050 -1770 5062 -1718
rect 5114 -1770 5126 -1718
rect 5178 -1770 5227 -1718
rect 5279 -1770 5291 -1718
rect 5343 -1770 5355 -1718
rect 5407 -1770 5436 -1718
rect 4728 -1787 5436 -1770
rect 5525 -1543 6199 -1537
rect 5525 -1577 5792 -1543
rect 5826 -1577 5864 -1543
rect 5898 -1561 6050 -1543
rect 5525 -1613 5893 -1577
rect 5945 -1613 5957 -1561
rect 6009 -1613 6021 -1561
rect 6084 -1577 6122 -1543
rect 6156 -1577 6199 -1543
rect 6073 -1613 6199 -1577
rect 5525 -1633 6199 -1613
rect 6456 -1543 6893 -1528
rect 6456 -1577 6555 -1543
rect 6589 -1577 6627 -1543
rect 6661 -1566 6893 -1543
rect 6661 -1577 6834 -1566
rect 6456 -1600 6834 -1577
rect 6868 -1600 6893 -1566
rect 5525 -1850 5660 -1633
rect 6456 -1638 6893 -1600
rect 6456 -1672 6834 -1638
rect 6868 -1672 6893 -1638
rect 4503 -1906 5660 -1850
rect 4503 -1940 4771 -1906
rect 4805 -1940 4843 -1906
rect 4877 -1940 5029 -1906
rect 5063 -1940 5101 -1906
rect 5135 -1940 5287 -1906
rect 5321 -1940 5359 -1906
rect 5393 -1940 5660 -1906
rect 4503 -1946 5660 -1940
rect 5749 -1718 6199 -1706
rect 5749 -1770 5893 -1718
rect 5945 -1770 5957 -1718
rect 6009 -1770 6021 -1718
rect 6073 -1770 6199 -1718
rect 5749 -1870 6199 -1770
rect 5749 -1906 5893 -1870
rect 5749 -1940 5792 -1906
rect 5826 -1940 5864 -1906
rect 5945 -1922 5957 -1870
rect 6009 -1922 6021 -1870
rect 6073 -1906 6199 -1870
rect 5898 -1940 6050 -1922
rect 6084 -1940 6122 -1906
rect 6156 -1940 6199 -1906
rect 5749 -1946 6199 -1940
rect 6456 -1710 6893 -1672
rect 6456 -1744 6834 -1710
rect 6868 -1744 6893 -1710
rect 6456 -1782 6893 -1744
rect 6456 -1816 6834 -1782
rect 6868 -1816 6893 -1782
rect 6456 -1854 6893 -1816
rect 6456 -1888 6834 -1854
rect 6868 -1888 6893 -1854
rect 6456 -1906 6893 -1888
rect 6456 -1940 6555 -1906
rect 6589 -1940 6627 -1906
rect 6661 -1926 6893 -1906
rect 6661 -1940 6834 -1926
rect -269 -2032 -244 -1998
rect -210 -2025 168 -1998
rect -210 -2032 -130 -2025
rect -269 -2059 -130 -2032
rect -96 -2059 128 -2025
rect 162 -2059 168 -2025
rect -269 -2070 168 -2059
rect -269 -2104 -244 -2070
rect -210 -2097 168 -2070
rect -210 -2104 -130 -2097
rect -269 -2131 -130 -2104
rect -96 -2131 128 -2097
rect 162 -2131 168 -2097
rect -269 -2142 168 -2131
rect -269 -2176 -244 -2142
rect -210 -2176 168 -2142
rect -269 -2214 168 -2176
rect -269 -2248 -244 -2214
rect -210 -2248 168 -2214
rect -269 -2286 168 -2248
rect -269 -2320 -244 -2286
rect -210 -2320 168 -2286
rect -269 -2358 168 -2320
rect -269 -2392 -244 -2358
rect -210 -2392 168 -2358
rect -269 -2430 168 -2392
rect -269 -2464 -244 -2430
rect -210 -2464 168 -2430
rect -269 -2502 168 -2464
rect -269 -2536 -244 -2502
rect -210 -2536 168 -2502
rect 369 -2025 415 -1978
rect 369 -2059 375 -2025
rect 409 -2059 415 -2025
rect 369 -2097 415 -2059
rect 369 -2131 375 -2097
rect 409 -2131 415 -2097
rect 369 -2446 415 -2131
rect 627 -2025 673 -1978
rect 627 -2059 633 -2025
rect 667 -2059 673 -2025
rect 627 -2097 673 -2059
rect 627 -2131 633 -2097
rect 667 -2131 673 -2097
rect 627 -2235 673 -2131
rect 885 -2025 931 -1978
rect 885 -2059 891 -2025
rect 925 -2059 931 -2025
rect 885 -2097 931 -2059
rect 885 -2131 891 -2097
rect 925 -2131 931 -2097
rect 553 -2245 749 -2235
rect 553 -2297 560 -2245
rect 612 -2297 624 -2245
rect 676 -2297 688 -2245
rect 740 -2297 749 -2245
rect 553 -2305 749 -2297
rect 885 -2446 931 -2131
rect 1132 -2025 1178 -1978
rect 1132 -2059 1138 -2025
rect 1172 -2059 1178 -2025
rect 1132 -2097 1178 -2059
rect 1132 -2131 1138 -2097
rect 1172 -2131 1178 -2097
rect 1132 -2334 1178 -2131
rect 1390 -2025 1436 -1978
rect 1390 -2059 1396 -2025
rect 1430 -2059 1436 -2025
rect 1390 -2097 1436 -2059
rect 1390 -2131 1396 -2097
rect 1430 -2131 1436 -2097
rect 1057 -2344 1253 -2334
rect 1057 -2396 1064 -2344
rect 1116 -2396 1128 -2344
rect 1180 -2396 1192 -2344
rect 1244 -2396 1253 -2344
rect 1057 -2404 1253 -2396
rect 369 -2456 931 -2446
rect 369 -2508 376 -2456
rect 428 -2508 440 -2456
rect 492 -2508 504 -2456
rect 556 -2508 742 -2456
rect 794 -2508 806 -2456
rect 858 -2508 870 -2456
rect 922 -2508 931 -2456
rect 369 -2516 931 -2508
rect -269 -2574 168 -2536
rect 1390 -2545 1436 -2131
rect 1648 -2025 1694 -1978
rect 1648 -2059 1654 -2025
rect 1688 -2059 1694 -2025
rect 1648 -2097 1694 -2059
rect 1648 -2131 1654 -2097
rect 1688 -2131 1694 -2097
rect 1648 -2334 1694 -2131
rect 1906 -2025 1952 -1978
rect 1906 -2059 1912 -2025
rect 1946 -2059 1952 -2025
rect 1906 -2097 1952 -2059
rect 1906 -2131 1912 -2097
rect 1946 -2131 1952 -2097
rect 1574 -2344 1770 -2334
rect 1574 -2396 1581 -2344
rect 1633 -2396 1645 -2344
rect 1697 -2396 1709 -2344
rect 1761 -2396 1770 -2344
rect 1574 -2404 1770 -2396
rect 1906 -2545 1952 -2131
rect 2153 -2025 2199 -1978
rect 2153 -2059 2159 -2025
rect 2193 -2059 2199 -2025
rect 2153 -2097 2199 -2059
rect 2153 -2131 2159 -2097
rect 2193 -2131 2199 -2097
rect 2153 -2446 2199 -2131
rect 2411 -2025 2457 -1978
rect 2411 -2059 2417 -2025
rect 2451 -2059 2457 -2025
rect 2411 -2097 2457 -2059
rect 2411 -2131 2417 -2097
rect 2451 -2131 2457 -2097
rect 2411 -2235 2457 -2131
rect 2669 -2025 2715 -1978
rect 2669 -2059 2675 -2025
rect 2709 -2059 2715 -2025
rect 2669 -2097 2715 -2059
rect 2669 -2131 2675 -2097
rect 2709 -2131 2715 -2097
rect 2337 -2245 2533 -2235
rect 2337 -2297 2344 -2245
rect 2396 -2297 2408 -2245
rect 2460 -2297 2472 -2245
rect 2524 -2297 2533 -2245
rect 2337 -2305 2533 -2297
rect 2669 -2446 2715 -2131
rect 2153 -2456 2715 -2446
rect 2153 -2508 2160 -2456
rect 2212 -2508 2224 -2456
rect 2276 -2508 2288 -2456
rect 2340 -2508 2526 -2456
rect 2578 -2508 2590 -2456
rect 2642 -2508 2654 -2456
rect 2706 -2508 2715 -2456
rect 2153 -2516 2715 -2508
rect 2917 -1998 3707 -1960
rect 6456 -1960 6834 -1940
rect 6868 -1960 6893 -1926
rect 2917 -2025 3295 -1998
rect 2917 -2059 2923 -2025
rect 2957 -2059 3181 -2025
rect 3215 -2032 3295 -2025
rect 3329 -2025 3707 -1998
rect 3329 -2032 3409 -2025
rect 3215 -2059 3409 -2032
rect 3443 -2059 3667 -2025
rect 3701 -2059 3707 -2025
rect 2917 -2070 3707 -2059
rect 2917 -2097 3295 -2070
rect 2917 -2131 2923 -2097
rect 2957 -2131 3181 -2097
rect 3215 -2104 3295 -2097
rect 3329 -2097 3707 -2070
rect 3329 -2104 3409 -2097
rect 3215 -2131 3409 -2104
rect 3443 -2131 3667 -2097
rect 3701 -2131 3707 -2097
rect 2917 -2142 3707 -2131
rect 2917 -2176 3295 -2142
rect 3329 -2176 3707 -2142
rect 2917 -2214 3707 -2176
rect 2917 -2248 3295 -2214
rect 3329 -2248 3707 -2214
rect 2917 -2286 3707 -2248
rect 2917 -2320 3295 -2286
rect 3329 -2320 3707 -2286
rect 2917 -2358 3707 -2320
rect 2917 -2392 3295 -2358
rect 3329 -2392 3707 -2358
rect 2917 -2430 3707 -2392
rect 2917 -2464 3295 -2430
rect 3329 -2464 3707 -2430
rect 2917 -2502 3707 -2464
rect 2917 -2536 3295 -2502
rect 3329 -2536 3707 -2502
rect 3909 -2025 3955 -1978
rect 3909 -2059 3915 -2025
rect 3949 -2059 3955 -2025
rect 3909 -2097 3955 -2059
rect 3909 -2131 3915 -2097
rect 3949 -2131 3955 -2097
rect 3909 -2446 3955 -2131
rect 4167 -2025 4213 -1978
rect 4167 -2059 4173 -2025
rect 4207 -2059 4213 -2025
rect 4167 -2097 4213 -2059
rect 4167 -2131 4173 -2097
rect 4207 -2131 4213 -2097
rect 4167 -2235 4213 -2131
rect 4425 -2025 4471 -1978
rect 4425 -2059 4431 -2025
rect 4465 -2059 4471 -2025
rect 4425 -2097 4471 -2059
rect 4425 -2131 4431 -2097
rect 4465 -2131 4471 -2097
rect 4091 -2245 4287 -2235
rect 4091 -2297 4100 -2245
rect 4152 -2297 4164 -2245
rect 4216 -2297 4228 -2245
rect 4280 -2297 4287 -2245
rect 4091 -2305 4287 -2297
rect 4425 -2446 4471 -2131
rect 3909 -2456 4471 -2446
rect 3909 -2508 3918 -2456
rect 3970 -2508 3982 -2456
rect 4034 -2508 4046 -2456
rect 4098 -2508 4284 -2456
rect 4336 -2508 4348 -2456
rect 4400 -2508 4412 -2456
rect 4464 -2508 4471 -2456
rect 3909 -2516 4471 -2508
rect 4672 -2025 4718 -1978
rect 4672 -2059 4678 -2025
rect 4712 -2059 4718 -2025
rect 4672 -2097 4718 -2059
rect 4672 -2131 4678 -2097
rect 4712 -2131 4718 -2097
rect -269 -2608 -244 -2574
rect -210 -2608 168 -2574
rect -269 -2646 168 -2608
rect 1314 -2555 1510 -2545
rect 1314 -2607 1321 -2555
rect 1373 -2607 1385 -2555
rect 1437 -2607 1449 -2555
rect 1501 -2607 1510 -2555
rect 1314 -2615 1510 -2607
rect 1831 -2555 2027 -2545
rect 1831 -2607 1838 -2555
rect 1890 -2607 1902 -2555
rect 1954 -2607 1966 -2555
rect 2018 -2607 2027 -2555
rect 1831 -2615 2027 -2607
rect 2917 -2574 3707 -2536
rect 4672 -2545 4718 -2131
rect 4930 -2025 4976 -1978
rect 4930 -2059 4936 -2025
rect 4970 -2059 4976 -2025
rect 4930 -2097 4976 -2059
rect 4930 -2131 4936 -2097
rect 4970 -2131 4976 -2097
rect 4930 -2334 4976 -2131
rect 5188 -2025 5234 -1978
rect 5188 -2059 5194 -2025
rect 5228 -2059 5234 -2025
rect 5188 -2097 5234 -2059
rect 5188 -2131 5194 -2097
rect 5228 -2131 5234 -2097
rect 4854 -2344 5050 -2334
rect 4854 -2396 4863 -2344
rect 4915 -2396 4927 -2344
rect 4979 -2396 4991 -2344
rect 5043 -2396 5050 -2344
rect 4854 -2404 5050 -2396
rect 5188 -2545 5234 -2131
rect 5446 -2025 5492 -1978
rect 5446 -2059 5452 -2025
rect 5486 -2059 5492 -2025
rect 5446 -2097 5492 -2059
rect 5446 -2131 5452 -2097
rect 5486 -2131 5492 -2097
rect 5446 -2334 5492 -2131
rect 5693 -2025 5739 -1978
rect 5693 -2059 5699 -2025
rect 5733 -2059 5739 -2025
rect 5693 -2097 5739 -2059
rect 5693 -2131 5699 -2097
rect 5733 -2131 5739 -2097
rect 5371 -2344 5567 -2334
rect 5371 -2396 5380 -2344
rect 5432 -2396 5444 -2344
rect 5496 -2396 5508 -2344
rect 5560 -2396 5567 -2344
rect 5371 -2404 5567 -2396
rect 5693 -2446 5739 -2131
rect 5951 -2025 5997 -1978
rect 5951 -2059 5957 -2025
rect 5991 -2059 5997 -2025
rect 5951 -2097 5997 -2059
rect 5951 -2131 5957 -2097
rect 5991 -2131 5997 -2097
rect 5951 -2235 5997 -2131
rect 6209 -2025 6255 -1978
rect 6209 -2059 6215 -2025
rect 6249 -2059 6255 -2025
rect 6209 -2097 6255 -2059
rect 6209 -2131 6215 -2097
rect 6249 -2131 6255 -2097
rect 5875 -2245 6071 -2235
rect 5875 -2297 5884 -2245
rect 5936 -2297 5948 -2245
rect 6000 -2297 6012 -2245
rect 6064 -2297 6071 -2245
rect 5875 -2305 6071 -2297
rect 6209 -2446 6255 -2131
rect 5693 -2456 6255 -2446
rect 5693 -2508 5702 -2456
rect 5754 -2508 5766 -2456
rect 5818 -2508 5830 -2456
rect 5882 -2508 6068 -2456
rect 6120 -2508 6132 -2456
rect 6184 -2508 6196 -2456
rect 6248 -2508 6255 -2456
rect 5693 -2516 6255 -2508
rect 6456 -1998 6893 -1960
rect 6456 -2025 6834 -1998
rect 6456 -2059 6462 -2025
rect 6496 -2059 6720 -2025
rect 6754 -2032 6834 -2025
rect 6868 -2032 6893 -1998
rect 6754 -2059 6893 -2032
rect 6456 -2070 6893 -2059
rect 6456 -2097 6834 -2070
rect 6456 -2131 6462 -2097
rect 6496 -2131 6720 -2097
rect 6754 -2104 6834 -2097
rect 6868 -2104 6893 -2070
rect 6754 -2131 6893 -2104
rect 6456 -2142 6893 -2131
rect 6456 -2176 6834 -2142
rect 6868 -2176 6893 -2142
rect 6456 -2214 6893 -2176
rect 6456 -2248 6834 -2214
rect 6868 -2248 6893 -2214
rect 6456 -2286 6893 -2248
rect 6456 -2320 6834 -2286
rect 6868 -2320 6893 -2286
rect 6456 -2358 6893 -2320
rect 6456 -2392 6834 -2358
rect 6868 -2392 6893 -2358
rect 6456 -2430 6893 -2392
rect 6456 -2464 6834 -2430
rect 6868 -2464 6893 -2430
rect 6456 -2502 6893 -2464
rect 6456 -2536 6834 -2502
rect 6868 -2536 6893 -2502
rect 2917 -2608 3295 -2574
rect 3329 -2608 3707 -2574
rect -269 -2680 -244 -2646
rect -210 -2680 168 -2646
rect -269 -2718 168 -2680
rect 2917 -2646 3707 -2608
rect 4597 -2555 4793 -2545
rect 4597 -2607 4606 -2555
rect 4658 -2607 4670 -2555
rect 4722 -2607 4734 -2555
rect 4786 -2607 4793 -2555
rect 4597 -2615 4793 -2607
rect 5114 -2555 5310 -2545
rect 5114 -2607 5123 -2555
rect 5175 -2607 5187 -2555
rect 5239 -2607 5251 -2555
rect 5303 -2607 5310 -2555
rect 5114 -2615 5310 -2607
rect 6456 -2574 6893 -2536
rect 6456 -2608 6834 -2574
rect 6868 -2608 6893 -2574
rect 2917 -2680 3295 -2646
rect 3329 -2680 3707 -2646
rect -269 -2752 -244 -2718
rect -210 -2751 168 -2718
rect -210 -2752 -130 -2751
rect -269 -2785 -130 -2752
rect -96 -2785 128 -2751
rect 162 -2785 168 -2751
rect -269 -2790 168 -2785
rect -269 -2824 -244 -2790
rect -210 -2823 168 -2790
rect -210 -2824 -130 -2823
rect -269 -2857 -130 -2824
rect -96 -2857 128 -2823
rect 162 -2857 168 -2823
rect -269 -2862 168 -2857
rect -269 -2896 -244 -2862
rect -210 -2896 168 -2862
rect -269 -2934 168 -2896
rect -269 -2968 -244 -2934
rect -210 -2936 168 -2934
rect 369 -2751 415 -2704
rect 369 -2785 375 -2751
rect 409 -2785 415 -2751
rect 369 -2823 415 -2785
rect 369 -2857 375 -2823
rect 409 -2857 415 -2823
rect 369 -2936 415 -2857
rect 627 -2751 673 -2704
rect 627 -2785 633 -2751
rect 667 -2785 673 -2751
rect 627 -2823 673 -2785
rect 627 -2857 633 -2823
rect 667 -2857 673 -2823
rect 627 -2936 673 -2857
rect 885 -2751 931 -2704
rect 885 -2785 891 -2751
rect 925 -2785 931 -2751
rect 885 -2823 931 -2785
rect 885 -2857 891 -2823
rect 925 -2857 931 -2823
rect 885 -2936 931 -2857
rect 1132 -2751 1178 -2704
rect 1132 -2785 1138 -2751
rect 1172 -2785 1178 -2751
rect 1132 -2823 1178 -2785
rect 1132 -2857 1138 -2823
rect 1172 -2857 1178 -2823
rect 1132 -2936 1178 -2857
rect 1390 -2751 1436 -2704
rect 1390 -2785 1396 -2751
rect 1430 -2785 1436 -2751
rect 1390 -2823 1436 -2785
rect 1390 -2857 1396 -2823
rect 1430 -2857 1436 -2823
rect 1390 -2936 1436 -2857
rect 1648 -2751 1694 -2704
rect 1648 -2785 1654 -2751
rect 1688 -2785 1694 -2751
rect 1648 -2823 1694 -2785
rect 1648 -2857 1654 -2823
rect 1688 -2857 1694 -2823
rect 1648 -2936 1694 -2857
rect 1906 -2751 1952 -2704
rect 1906 -2785 1912 -2751
rect 1946 -2785 1952 -2751
rect 1906 -2823 1952 -2785
rect 1906 -2857 1912 -2823
rect 1946 -2857 1952 -2823
rect 1906 -2936 1952 -2857
rect 2153 -2751 2199 -2704
rect 2153 -2785 2159 -2751
rect 2193 -2785 2199 -2751
rect 2153 -2823 2199 -2785
rect 2153 -2857 2159 -2823
rect 2193 -2857 2199 -2823
rect 2153 -2936 2199 -2857
rect 2411 -2751 2457 -2704
rect 2411 -2785 2417 -2751
rect 2451 -2785 2457 -2751
rect 2411 -2823 2457 -2785
rect 2411 -2857 2417 -2823
rect 2451 -2857 2457 -2823
rect 2411 -2936 2457 -2857
rect 2669 -2751 2715 -2704
rect 2669 -2785 2675 -2751
rect 2709 -2785 2715 -2751
rect 2669 -2823 2715 -2785
rect 2669 -2857 2675 -2823
rect 2709 -2857 2715 -2823
rect 2669 -2936 2715 -2857
rect 2917 -2718 3707 -2680
rect 6456 -2646 6893 -2608
rect 6456 -2680 6834 -2646
rect 6868 -2680 6893 -2646
rect 2917 -2751 3295 -2718
rect 2917 -2785 2923 -2751
rect 2957 -2785 3181 -2751
rect 3215 -2752 3295 -2751
rect 3329 -2751 3707 -2718
rect 3329 -2752 3409 -2751
rect 3215 -2785 3409 -2752
rect 3443 -2785 3667 -2751
rect 3701 -2785 3707 -2751
rect 2917 -2790 3707 -2785
rect 2917 -2823 3295 -2790
rect 2917 -2857 2923 -2823
rect 2957 -2857 3181 -2823
rect 3215 -2824 3295 -2823
rect 3329 -2823 3707 -2790
rect 3329 -2824 3409 -2823
rect 3215 -2857 3409 -2824
rect 3443 -2857 3667 -2823
rect 3701 -2857 3707 -2823
rect 2917 -2862 3707 -2857
rect 2917 -2896 3295 -2862
rect 3329 -2896 3707 -2862
rect 2917 -2934 3707 -2896
rect 2917 -2936 3295 -2934
rect -210 -2942 3295 -2936
rect -210 -2968 -37 -2942
rect -269 -2976 -37 -2968
rect -3 -2976 35 -2942
rect 69 -2976 468 -2942
rect 502 -2976 540 -2942
rect 574 -2976 726 -2942
rect 760 -2976 798 -2942
rect 832 -2976 1231 -2942
rect 1265 -2976 1303 -2942
rect 1337 -2976 1489 -2942
rect 1523 -2976 1561 -2942
rect 1595 -2976 1747 -2942
rect 1781 -2976 1819 -2942
rect 1853 -2976 2252 -2942
rect 2286 -2976 2324 -2942
rect 2358 -2976 2510 -2942
rect 2544 -2976 2582 -2942
rect 2616 -2976 3016 -2942
rect 3050 -2976 3088 -2942
rect 3122 -2968 3295 -2942
rect 3329 -2936 3707 -2934
rect 3909 -2751 3955 -2704
rect 3909 -2785 3915 -2751
rect 3949 -2785 3955 -2751
rect 3909 -2823 3955 -2785
rect 3909 -2857 3915 -2823
rect 3949 -2857 3955 -2823
rect 3909 -2936 3955 -2857
rect 4167 -2751 4213 -2704
rect 4167 -2785 4173 -2751
rect 4207 -2785 4213 -2751
rect 4167 -2823 4213 -2785
rect 4167 -2857 4173 -2823
rect 4207 -2857 4213 -2823
rect 4167 -2936 4213 -2857
rect 4425 -2751 4471 -2704
rect 4425 -2785 4431 -2751
rect 4465 -2785 4471 -2751
rect 4425 -2823 4471 -2785
rect 4425 -2857 4431 -2823
rect 4465 -2857 4471 -2823
rect 4425 -2936 4471 -2857
rect 4672 -2751 4718 -2704
rect 4672 -2785 4678 -2751
rect 4712 -2785 4718 -2751
rect 4672 -2823 4718 -2785
rect 4672 -2857 4678 -2823
rect 4712 -2857 4718 -2823
rect 4672 -2936 4718 -2857
rect 4930 -2751 4976 -2704
rect 4930 -2785 4936 -2751
rect 4970 -2785 4976 -2751
rect 4930 -2823 4976 -2785
rect 4930 -2857 4936 -2823
rect 4970 -2857 4976 -2823
rect 4930 -2936 4976 -2857
rect 5188 -2751 5234 -2704
rect 5188 -2785 5194 -2751
rect 5228 -2785 5234 -2751
rect 5188 -2823 5234 -2785
rect 5188 -2857 5194 -2823
rect 5228 -2857 5234 -2823
rect 5188 -2936 5234 -2857
rect 5446 -2751 5492 -2704
rect 5446 -2785 5452 -2751
rect 5486 -2785 5492 -2751
rect 5446 -2823 5492 -2785
rect 5446 -2857 5452 -2823
rect 5486 -2857 5492 -2823
rect 5446 -2936 5492 -2857
rect 5693 -2751 5739 -2704
rect 5693 -2785 5699 -2751
rect 5733 -2785 5739 -2751
rect 5693 -2823 5739 -2785
rect 5693 -2857 5699 -2823
rect 5733 -2857 5739 -2823
rect 5693 -2936 5739 -2857
rect 5951 -2751 5997 -2704
rect 5951 -2785 5957 -2751
rect 5991 -2785 5997 -2751
rect 5951 -2823 5997 -2785
rect 5951 -2857 5957 -2823
rect 5991 -2857 5997 -2823
rect 5951 -2936 5997 -2857
rect 6209 -2751 6255 -2704
rect 6209 -2785 6215 -2751
rect 6249 -2785 6255 -2751
rect 6209 -2823 6255 -2785
rect 6209 -2857 6215 -2823
rect 6249 -2857 6255 -2823
rect 6209 -2936 6255 -2857
rect 6456 -2718 6893 -2680
rect 6456 -2751 6834 -2718
rect 6456 -2785 6462 -2751
rect 6496 -2785 6720 -2751
rect 6754 -2752 6834 -2751
rect 6868 -2752 6893 -2718
rect 6754 -2785 6893 -2752
rect 6456 -2790 6893 -2785
rect 6456 -2823 6834 -2790
rect 6456 -2857 6462 -2823
rect 6496 -2857 6720 -2823
rect 6754 -2824 6834 -2823
rect 6868 -2824 6893 -2790
rect 6754 -2857 6893 -2824
rect 6456 -2862 6893 -2857
rect 6456 -2896 6834 -2862
rect 6868 -2896 6893 -2862
rect 6456 -2934 6893 -2896
rect 6456 -2936 6834 -2934
rect 3329 -2942 6834 -2936
rect 3329 -2968 3502 -2942
rect 3122 -2976 3502 -2968
rect 3536 -2976 3574 -2942
rect 3608 -2976 4008 -2942
rect 4042 -2976 4080 -2942
rect 4114 -2976 4266 -2942
rect 4300 -2976 4338 -2942
rect 4372 -2976 4771 -2942
rect 4805 -2976 4843 -2942
rect 4877 -2976 5029 -2942
rect 5063 -2976 5101 -2942
rect 5135 -2976 5287 -2942
rect 5321 -2976 5359 -2942
rect 5393 -2976 5792 -2942
rect 5826 -2976 5864 -2942
rect 5898 -2976 6050 -2942
rect 6084 -2976 6122 -2942
rect 6156 -2976 6555 -2942
rect 6589 -2976 6627 -2942
rect 6661 -2968 6834 -2942
rect 6868 -2968 6893 -2934
rect 6661 -2976 6893 -2968
rect -269 -3041 6893 -2976
rect -269 -3075 -80 -3041
rect -46 -3075 -8 -3041
rect 26 -3075 64 -3041
rect 98 -3075 136 -3041
rect 170 -3075 208 -3041
rect 242 -3075 280 -3041
rect 314 -3075 352 -3041
rect 386 -3075 424 -3041
rect 458 -3075 496 -3041
rect 530 -3075 568 -3041
rect 602 -3075 640 -3041
rect 674 -3075 712 -3041
rect 746 -3075 784 -3041
rect 818 -3075 856 -3041
rect 890 -3075 928 -3041
rect 962 -3075 1000 -3041
rect 1034 -3075 1072 -3041
rect 1106 -3075 1144 -3041
rect 1178 -3075 1216 -3041
rect 1250 -3075 1288 -3041
rect 1322 -3075 1360 -3041
rect 1394 -3075 1432 -3041
rect 1466 -3075 1504 -3041
rect 1538 -3075 1576 -3041
rect 1610 -3075 1648 -3041
rect 1682 -3075 1720 -3041
rect 1754 -3075 1792 -3041
rect 1826 -3075 1864 -3041
rect 1898 -3075 1936 -3041
rect 1970 -3075 2008 -3041
rect 2042 -3075 2080 -3041
rect 2114 -3075 2152 -3041
rect 2186 -3075 2224 -3041
rect 2258 -3075 2296 -3041
rect 2330 -3075 2368 -3041
rect 2402 -3075 2440 -3041
rect 2474 -3075 2512 -3041
rect 2546 -3075 2584 -3041
rect 2618 -3075 2656 -3041
rect 2690 -3075 2728 -3041
rect 2762 -3075 2800 -3041
rect 2834 -3075 2872 -3041
rect 2906 -3075 2944 -3041
rect 2978 -3075 3016 -3041
rect 3050 -3075 3088 -3041
rect 3122 -3075 3160 -3041
rect 3194 -3075 3430 -3041
rect 3464 -3075 3502 -3041
rect 3536 -3075 3574 -3041
rect 3608 -3075 3646 -3041
rect 3680 -3075 3718 -3041
rect 3752 -3075 3790 -3041
rect 3824 -3075 3862 -3041
rect 3896 -3075 3934 -3041
rect 3968 -3075 4006 -3041
rect 4040 -3075 4078 -3041
rect 4112 -3075 4150 -3041
rect 4184 -3075 4222 -3041
rect 4256 -3075 4294 -3041
rect 4328 -3075 4366 -3041
rect 4400 -3075 4438 -3041
rect 4472 -3075 4510 -3041
rect 4544 -3075 4582 -3041
rect 4616 -3075 4654 -3041
rect 4688 -3075 4726 -3041
rect 4760 -3075 4798 -3041
rect 4832 -3075 4870 -3041
rect 4904 -3075 4942 -3041
rect 4976 -3075 5014 -3041
rect 5048 -3075 5086 -3041
rect 5120 -3075 5158 -3041
rect 5192 -3075 5230 -3041
rect 5264 -3075 5302 -3041
rect 5336 -3075 5374 -3041
rect 5408 -3075 5446 -3041
rect 5480 -3075 5518 -3041
rect 5552 -3075 5590 -3041
rect 5624 -3075 5662 -3041
rect 5696 -3075 5734 -3041
rect 5768 -3075 5806 -3041
rect 5840 -3075 5878 -3041
rect 5912 -3075 5950 -3041
rect 5984 -3075 6022 -3041
rect 6056 -3075 6094 -3041
rect 6128 -3075 6166 -3041
rect 6200 -3075 6238 -3041
rect 6272 -3075 6310 -3041
rect 6344 -3075 6382 -3041
rect 6416 -3075 6454 -3041
rect 6488 -3075 6526 -3041
rect 6560 -3075 6598 -3041
rect 6632 -3075 6670 -3041
rect 6704 -3075 6893 -3041
rect -269 -3100 6893 -3075
<< via1 >>
rect 1067 500 1119 552
rect 1131 500 1183 552
rect 1195 500 1247 552
rect 1584 500 1636 552
rect 1648 500 1700 552
rect 1712 500 1764 552
rect 378 384 430 436
rect 442 384 494 436
rect 506 384 558 436
rect 744 384 796 436
rect 808 384 860 436
rect 872 384 924 436
rect 560 159 612 211
rect 624 159 676 211
rect 688 159 740 211
rect 1324 258 1376 310
rect 1388 258 1440 310
rect 1452 258 1504 310
rect 4860 500 4912 552
rect 4924 500 4976 552
rect 4988 500 5040 552
rect 5377 500 5429 552
rect 5441 500 5493 552
rect 5505 500 5557 552
rect 2162 384 2214 436
rect 2226 384 2278 436
rect 2290 384 2342 436
rect 2528 384 2580 436
rect 2592 384 2644 436
rect 2656 384 2708 436
rect 1841 258 1893 310
rect 1905 258 1957 310
rect 1969 258 2021 310
rect 2345 159 2397 211
rect 2409 159 2461 211
rect 2473 159 2525 211
rect 3916 384 3968 436
rect 3980 384 4032 436
rect 4044 384 4096 436
rect 4282 384 4334 436
rect 4346 384 4398 436
rect 4410 384 4462 436
rect 4099 159 4151 211
rect 4163 159 4215 211
rect 4227 159 4279 211
rect 4603 258 4655 310
rect 4667 258 4719 310
rect 4731 258 4783 310
rect 5120 258 5172 310
rect 5184 258 5236 310
rect 5248 258 5300 310
rect 5700 384 5752 436
rect 5764 384 5816 436
rect 5828 384 5880 436
rect 6066 384 6118 436
rect 6130 384 6182 436
rect 6194 384 6246 436
rect 5884 159 5936 211
rect 5948 159 6000 211
rect 6012 159 6064 211
rect 551 -180 574 -164
rect 574 -180 603 -164
rect 551 -216 603 -180
rect 615 -216 667 -164
rect 679 -180 726 -164
rect 726 -180 731 -164
rect 679 -216 731 -180
rect 551 -367 603 -315
rect 615 -367 667 -315
rect 679 -367 731 -315
rect 551 -509 603 -473
rect 551 -525 574 -509
rect 574 -525 603 -509
rect 615 -525 667 -473
rect 679 -509 731 -473
rect 679 -525 726 -509
rect 726 -525 731 -509
rect 1217 -367 1269 -315
rect 1281 -367 1333 -315
rect 1345 -367 1397 -315
rect 1446 -367 1498 -315
rect 1510 -367 1562 -315
rect 1574 -367 1626 -315
rect 1684 -367 1736 -315
rect 1748 -367 1800 -315
rect 1812 -367 1864 -315
rect 2335 -180 2358 -164
rect 2358 -180 2387 -164
rect 2335 -216 2387 -180
rect 2399 -216 2451 -164
rect 2463 -180 2510 -164
rect 2510 -180 2515 -164
rect 2463 -216 2515 -180
rect 2335 -367 2387 -315
rect 2399 -367 2451 -315
rect 2463 -367 2515 -315
rect 4109 -180 4114 -164
rect 4114 -180 4161 -164
rect 4109 -216 4161 -180
rect 4173 -216 4225 -164
rect 4237 -180 4266 -164
rect 4266 -180 4289 -164
rect 4237 -216 4289 -180
rect 4109 -367 4161 -315
rect 4173 -367 4225 -315
rect 4237 -367 4289 -315
rect 2335 -509 2387 -473
rect 2335 -525 2358 -509
rect 2358 -525 2387 -509
rect 2399 -525 2451 -473
rect 2463 -509 2515 -473
rect 2463 -525 2510 -509
rect 2510 -525 2515 -509
rect 4109 -509 4161 -473
rect 4109 -525 4114 -509
rect 4114 -525 4161 -509
rect 4173 -525 4225 -473
rect 4237 -509 4289 -473
rect 4237 -525 4266 -509
rect 4266 -525 4289 -509
rect 4760 -367 4812 -315
rect 4824 -367 4876 -315
rect 4888 -367 4940 -315
rect 4998 -367 5050 -315
rect 5062 -367 5114 -315
rect 5126 -367 5178 -315
rect 5227 -367 5279 -315
rect 5291 -367 5343 -315
rect 5355 -367 5407 -315
rect 5893 -180 5898 -164
rect 5898 -180 5945 -164
rect 5893 -216 5945 -180
rect 5957 -216 6009 -164
rect 6021 -180 6050 -164
rect 6050 -180 6073 -164
rect 6021 -216 6073 -180
rect 5893 -367 5945 -315
rect 5957 -367 6009 -315
rect 6021 -367 6073 -315
rect 5893 -509 5945 -473
rect 5893 -525 5898 -509
rect 5898 -525 5945 -509
rect 5957 -525 6009 -473
rect 6021 -509 6073 -473
rect 6021 -525 6050 -509
rect 6050 -525 6073 -509
rect 560 -861 612 -809
rect 624 -861 676 -809
rect 688 -861 740 -809
rect 301 -1125 353 -1073
rect 365 -1125 417 -1073
rect 429 -1125 481 -1073
rect 1064 -1014 1116 -962
rect 1128 -1014 1180 -962
rect 1192 -1014 1244 -962
rect 820 -1125 872 -1073
rect 884 -1125 936 -1073
rect 948 -1125 1000 -1073
rect 1581 -1014 1633 -962
rect 1645 -1014 1697 -962
rect 1709 -1014 1761 -962
rect 1321 -1225 1373 -1173
rect 1385 -1225 1437 -1173
rect 1449 -1225 1501 -1173
rect 2344 -861 2396 -809
rect 2408 -861 2460 -809
rect 2472 -861 2524 -809
rect 2087 -1125 2139 -1073
rect 2151 -1125 2203 -1073
rect 2215 -1125 2267 -1073
rect 1838 -1225 1890 -1173
rect 1902 -1225 1954 -1173
rect 1966 -1225 2018 -1173
rect 2604 -1125 2656 -1073
rect 2668 -1125 2720 -1073
rect 2732 -1125 2784 -1073
rect 4100 -861 4152 -809
rect 4164 -861 4216 -809
rect 4228 -861 4280 -809
rect 3840 -1125 3892 -1073
rect 3904 -1125 3956 -1073
rect 3968 -1125 4020 -1073
rect 4357 -1125 4409 -1073
rect 4421 -1125 4473 -1073
rect 4485 -1125 4537 -1073
rect 4863 -1014 4915 -962
rect 4927 -1014 4979 -962
rect 4991 -1014 5043 -962
rect 4606 -1225 4658 -1173
rect 4670 -1225 4722 -1173
rect 4734 -1225 4786 -1173
rect 5380 -1014 5432 -962
rect 5444 -1014 5496 -962
rect 5508 -1014 5560 -962
rect 5123 -1225 5175 -1173
rect 5187 -1225 5239 -1173
rect 5251 -1225 5303 -1173
rect 5884 -861 5936 -809
rect 5948 -861 6000 -809
rect 6012 -861 6064 -809
rect 5624 -1125 5676 -1073
rect 5688 -1125 5740 -1073
rect 5752 -1125 5804 -1073
rect 6143 -1125 6195 -1073
rect 6207 -1125 6259 -1073
rect 6271 -1125 6323 -1073
rect 551 -1577 574 -1561
rect 574 -1577 603 -1561
rect 551 -1613 603 -1577
rect 615 -1613 667 -1561
rect 679 -1577 726 -1561
rect 726 -1577 731 -1561
rect 679 -1613 731 -1577
rect 551 -1770 603 -1718
rect 615 -1770 667 -1718
rect 679 -1770 731 -1718
rect 551 -1906 603 -1870
rect 551 -1922 574 -1906
rect 574 -1922 603 -1906
rect 615 -1922 667 -1870
rect 679 -1906 731 -1870
rect 679 -1922 726 -1906
rect 726 -1922 731 -1906
rect 1217 -1770 1269 -1718
rect 1281 -1770 1333 -1718
rect 1345 -1770 1397 -1718
rect 1446 -1770 1498 -1718
rect 1510 -1770 1562 -1718
rect 1574 -1770 1626 -1718
rect 1684 -1770 1736 -1718
rect 1748 -1770 1800 -1718
rect 1812 -1770 1864 -1718
rect 2335 -1577 2358 -1561
rect 2358 -1577 2387 -1561
rect 2335 -1613 2387 -1577
rect 2399 -1613 2451 -1561
rect 2463 -1577 2510 -1561
rect 2510 -1577 2515 -1561
rect 2463 -1613 2515 -1577
rect 4109 -1577 4114 -1561
rect 4114 -1577 4161 -1561
rect 4109 -1613 4161 -1577
rect 4173 -1613 4225 -1561
rect 4237 -1577 4266 -1561
rect 4266 -1577 4289 -1561
rect 4237 -1613 4289 -1577
rect 2335 -1770 2387 -1718
rect 2399 -1770 2451 -1718
rect 2463 -1770 2515 -1718
rect 2335 -1906 2387 -1870
rect 2335 -1922 2358 -1906
rect 2358 -1922 2387 -1906
rect 2399 -1922 2451 -1870
rect 2463 -1906 2515 -1870
rect 2463 -1922 2510 -1906
rect 2510 -1922 2515 -1906
rect 4109 -1770 4161 -1718
rect 4173 -1770 4225 -1718
rect 4237 -1770 4289 -1718
rect 4109 -1906 4161 -1870
rect 4109 -1922 4114 -1906
rect 4114 -1922 4161 -1906
rect 4173 -1922 4225 -1870
rect 4237 -1906 4289 -1870
rect 4237 -1922 4266 -1906
rect 4266 -1922 4289 -1906
rect 4760 -1770 4812 -1718
rect 4824 -1770 4876 -1718
rect 4888 -1770 4940 -1718
rect 4998 -1770 5050 -1718
rect 5062 -1770 5114 -1718
rect 5126 -1770 5178 -1718
rect 5227 -1770 5279 -1718
rect 5291 -1770 5343 -1718
rect 5355 -1770 5407 -1718
rect 5893 -1577 5898 -1561
rect 5898 -1577 5945 -1561
rect 5893 -1613 5945 -1577
rect 5957 -1613 6009 -1561
rect 6021 -1577 6050 -1561
rect 6050 -1577 6073 -1561
rect 6021 -1613 6073 -1577
rect 5893 -1770 5945 -1718
rect 5957 -1770 6009 -1718
rect 6021 -1770 6073 -1718
rect 5893 -1906 5945 -1870
rect 5893 -1922 5898 -1906
rect 5898 -1922 5945 -1906
rect 5957 -1922 6009 -1870
rect 6021 -1906 6073 -1870
rect 6021 -1922 6050 -1906
rect 6050 -1922 6073 -1906
rect 560 -2297 612 -2245
rect 624 -2297 676 -2245
rect 688 -2297 740 -2245
rect 1064 -2396 1116 -2344
rect 1128 -2396 1180 -2344
rect 1192 -2396 1244 -2344
rect 376 -2508 428 -2456
rect 440 -2508 492 -2456
rect 504 -2508 556 -2456
rect 742 -2508 794 -2456
rect 806 -2508 858 -2456
rect 870 -2508 922 -2456
rect 1581 -2396 1633 -2344
rect 1645 -2396 1697 -2344
rect 1709 -2396 1761 -2344
rect 2344 -2297 2396 -2245
rect 2408 -2297 2460 -2245
rect 2472 -2297 2524 -2245
rect 2160 -2508 2212 -2456
rect 2224 -2508 2276 -2456
rect 2288 -2508 2340 -2456
rect 2526 -2508 2578 -2456
rect 2590 -2508 2642 -2456
rect 2654 -2508 2706 -2456
rect 4100 -2297 4152 -2245
rect 4164 -2297 4216 -2245
rect 4228 -2297 4280 -2245
rect 3918 -2508 3970 -2456
rect 3982 -2508 4034 -2456
rect 4046 -2508 4098 -2456
rect 4284 -2508 4336 -2456
rect 4348 -2508 4400 -2456
rect 4412 -2508 4464 -2456
rect 1321 -2607 1373 -2555
rect 1385 -2607 1437 -2555
rect 1449 -2607 1501 -2555
rect 1838 -2607 1890 -2555
rect 1902 -2607 1954 -2555
rect 1966 -2607 2018 -2555
rect 4863 -2396 4915 -2344
rect 4927 -2396 4979 -2344
rect 4991 -2396 5043 -2344
rect 5380 -2396 5432 -2344
rect 5444 -2396 5496 -2344
rect 5508 -2396 5560 -2344
rect 5884 -2297 5936 -2245
rect 5948 -2297 6000 -2245
rect 6012 -2297 6064 -2245
rect 5702 -2508 5754 -2456
rect 5766 -2508 5818 -2456
rect 5830 -2508 5882 -2456
rect 6068 -2508 6120 -2456
rect 6132 -2508 6184 -2456
rect 6196 -2508 6248 -2456
rect 4606 -2607 4658 -2555
rect 4670 -2607 4722 -2555
rect 4734 -2607 4786 -2555
rect 5123 -2607 5175 -2555
rect 5187 -2607 5239 -2555
rect 5251 -2607 5303 -2555
<< metal2 >>
rect -269 552 6893 560
rect -269 538 1067 552
rect -269 482 -229 538
rect -173 482 -149 538
rect -93 482 -69 538
rect -13 500 1067 538
rect 1119 500 1131 552
rect 1183 500 1195 552
rect 1247 500 1584 552
rect 1636 500 1648 552
rect 1700 500 1712 552
rect 1764 500 4860 552
rect 4912 500 4924 552
rect 4976 500 4988 552
rect 5040 500 5377 552
rect 5429 500 5441 552
rect 5493 500 5505 552
rect 5557 538 6893 552
rect 5557 500 6637 538
rect -13 490 6637 500
rect -13 482 31 490
rect -269 460 31 482
rect 6593 482 6637 490
rect 6693 482 6717 538
rect 6773 482 6797 538
rect 6853 482 6893 538
rect 6593 460 6893 482
rect 3054 444 3570 453
rect 369 436 6255 444
rect 369 384 378 436
rect 430 384 442 436
rect 494 384 506 436
rect 558 384 744 436
rect 796 384 808 436
rect 860 384 872 436
rect 924 384 2162 436
rect 2214 384 2226 436
rect 2278 384 2290 436
rect 2342 384 2528 436
rect 2580 384 2592 436
rect 2644 384 2656 436
rect 2708 431 3916 436
rect 2708 384 3094 431
rect 369 375 3094 384
rect 3150 375 3174 431
rect 3230 375 3254 431
rect 3310 375 3394 431
rect 3450 375 3474 431
rect 3530 384 3916 431
rect 3968 384 3980 436
rect 4032 384 4044 436
rect 4096 384 4282 436
rect 4334 384 4346 436
rect 4398 384 4410 436
rect 4462 384 5700 436
rect 5752 384 5764 436
rect 5816 384 5828 436
rect 5880 384 6066 436
rect 6118 384 6130 436
rect 6182 384 6194 436
rect 6246 384 6255 436
rect 3530 375 6255 384
rect 369 374 6255 375
rect 3054 353 3570 374
rect 163 310 6461 318
rect 163 296 1324 310
rect 163 240 203 296
rect 259 240 283 296
rect 339 240 363 296
rect 419 258 1324 296
rect 1376 258 1388 310
rect 1440 258 1452 310
rect 1504 258 1841 310
rect 1893 258 1905 310
rect 1957 258 1969 310
rect 2021 258 4603 310
rect 4655 258 4667 310
rect 4719 258 4731 310
rect 4783 258 5120 310
rect 5172 258 5184 310
rect 5236 258 5248 310
rect 5300 296 6461 310
rect 5300 258 6205 296
rect 419 248 6205 258
rect 419 240 463 248
rect 163 218 463 240
rect 6161 240 6205 248
rect 6261 240 6285 296
rect 6341 240 6365 296
rect 6421 240 6461 296
rect 551 211 6073 219
rect 6161 218 6461 240
rect 551 159 560 211
rect 612 159 624 211
rect 676 159 688 211
rect 740 159 2345 211
rect 2397 159 2409 211
rect 2461 159 2473 211
rect 2525 197 4099 211
rect 2525 159 2662 197
rect 551 149 2662 159
rect 2622 141 2662 149
rect 2718 141 2742 197
rect 2798 141 2822 197
rect 2878 149 3746 197
rect 2878 141 2922 149
rect 2622 119 2922 141
rect 3702 141 3746 149
rect 3802 141 3826 197
rect 3882 141 3906 197
rect 3962 159 4099 197
rect 4151 159 4163 211
rect 4215 159 4227 211
rect 4279 159 5884 211
rect 5936 159 5948 211
rect 6000 159 6012 211
rect 6064 159 6073 211
rect 3962 149 6073 159
rect 3962 141 4002 149
rect 3702 119 4002 141
rect 1906 -140 2206 -136
rect 4418 -140 4718 -136
rect 425 -158 6199 -140
rect 425 -164 1946 -158
rect 425 -216 551 -164
rect 603 -216 615 -164
rect 667 -216 679 -164
rect 731 -214 1946 -164
rect 2002 -214 2026 -158
rect 2082 -214 2106 -158
rect 2162 -164 4462 -158
rect 2162 -214 2335 -164
rect 731 -216 2335 -214
rect 2387 -216 2399 -164
rect 2451 -216 2463 -164
rect 2515 -216 4109 -164
rect 4161 -216 4173 -164
rect 4225 -216 4237 -164
rect 4289 -214 4462 -164
rect 4518 -214 4542 -158
rect 4598 -214 4622 -158
rect 4678 -164 6199 -158
rect 4678 -214 5893 -164
rect 4289 -216 5893 -214
rect 5945 -216 5957 -164
rect 6009 -216 6021 -164
rect 6073 -216 6199 -164
rect 425 -236 6199 -216
rect 425 -315 6199 -299
rect 425 -367 551 -315
rect 603 -367 615 -315
rect 667 -367 679 -315
rect 731 -367 1217 -315
rect 1269 -367 1281 -315
rect 1333 -367 1345 -315
rect 1397 -367 1446 -315
rect 1498 -367 1510 -315
rect 1562 -367 1574 -315
rect 1626 -367 1684 -315
rect 1736 -367 1748 -315
rect 1800 -367 1812 -315
rect 1864 -321 2335 -315
rect 1864 -367 1946 -321
rect 425 -377 1946 -367
rect 2002 -377 2026 -321
rect 2082 -377 2106 -321
rect 2162 -367 2335 -321
rect 2387 -367 2399 -315
rect 2451 -367 2463 -315
rect 2515 -367 4109 -315
rect 4161 -367 4173 -315
rect 4225 -367 4237 -315
rect 4289 -321 4760 -315
rect 4289 -367 4462 -321
rect 2162 -377 4462 -367
rect 4518 -377 4542 -321
rect 4598 -377 4622 -321
rect 4678 -367 4760 -321
rect 4812 -367 4824 -315
rect 4876 -367 4888 -315
rect 4940 -367 4998 -315
rect 5050 -367 5062 -315
rect 5114 -367 5126 -315
rect 5178 -367 5227 -315
rect 5279 -367 5291 -315
rect 5343 -367 5355 -315
rect 5407 -367 5893 -315
rect 5945 -367 5957 -315
rect 6009 -367 6021 -315
rect 6073 -367 6199 -315
rect 4678 -377 6199 -367
rect 425 -380 6199 -377
rect 1906 -399 2206 -380
rect 4418 -399 4718 -380
rect 425 -473 6199 -453
rect 425 -525 551 -473
rect 603 -525 615 -473
rect 667 -525 679 -473
rect 731 -475 2335 -473
rect 731 -525 919 -475
rect 425 -531 919 -525
rect 975 -531 999 -475
rect 1055 -531 1079 -475
rect 1135 -525 2335 -475
rect 2387 -525 2399 -473
rect 2451 -525 2463 -473
rect 2515 -525 4109 -473
rect 4161 -525 4173 -473
rect 4225 -525 4237 -473
rect 4289 -475 5893 -473
rect 4289 -525 5489 -475
rect 1135 -531 5489 -525
rect 5545 -531 5569 -475
rect 5625 -531 5649 -475
rect 5705 -525 5893 -475
rect 5945 -525 5957 -473
rect 6009 -525 6021 -473
rect 6073 -525 6199 -473
rect 5705 -531 6199 -525
rect 425 -549 6199 -531
rect 879 -553 1179 -549
rect 5445 -553 5745 -549
rect 163 -791 463 -769
rect 163 -847 203 -791
rect 259 -847 283 -791
rect 339 -847 363 -791
rect 419 -799 463 -791
rect 6161 -791 6461 -769
rect 6161 -799 6205 -791
rect 419 -809 6205 -799
rect 419 -847 560 -809
rect 163 -861 560 -847
rect 612 -861 624 -809
rect 676 -861 688 -809
rect 740 -861 2344 -809
rect 2396 -861 2408 -809
rect 2460 -861 2472 -809
rect 2524 -861 4100 -809
rect 4152 -861 4164 -809
rect 4216 -861 4228 -809
rect 4280 -861 5884 -809
rect 5936 -861 5948 -809
rect 6000 -861 6012 -809
rect 6064 -847 6205 -809
rect 6261 -847 6285 -791
rect 6341 -847 6365 -791
rect 6421 -847 6461 -791
rect 6064 -861 6461 -847
rect 163 -869 6461 -861
rect 2622 -944 2922 -922
rect 2622 -952 2662 -944
rect 1057 -962 2662 -952
rect 1057 -1014 1064 -962
rect 1116 -1014 1128 -962
rect 1180 -1014 1192 -962
rect 1244 -1014 1581 -962
rect 1633 -1014 1645 -962
rect 1697 -1014 1709 -962
rect 1761 -1000 2662 -962
rect 2718 -1000 2742 -944
rect 2798 -1000 2822 -944
rect 2878 -952 2922 -944
rect 3702 -944 4002 -922
rect 3702 -952 3746 -944
rect 2878 -1000 3746 -952
rect 3802 -1000 3826 -944
rect 3882 -1000 3906 -944
rect 3962 -952 4002 -944
rect 3962 -962 5567 -952
rect 3962 -1000 4863 -962
rect 1761 -1014 4863 -1000
rect 4915 -1014 4927 -962
rect 4979 -1014 4991 -962
rect 5043 -1014 5380 -962
rect 5432 -1014 5444 -962
rect 5496 -1014 5508 -962
rect 5560 -1014 5567 -962
rect 1057 -1022 5567 -1014
rect -269 -1055 31 -1033
rect -269 -1111 -229 -1055
rect -173 -1111 -149 -1055
rect -93 -1111 -69 -1055
rect -13 -1063 31 -1055
rect 6593 -1055 6893 -1033
rect 6593 -1063 6637 -1055
rect -13 -1073 6637 -1063
rect -13 -1111 301 -1073
rect -269 -1125 301 -1111
rect 353 -1125 365 -1073
rect 417 -1125 429 -1073
rect 481 -1125 820 -1073
rect 872 -1125 884 -1073
rect 936 -1125 948 -1073
rect 1000 -1125 2087 -1073
rect 2139 -1125 2151 -1073
rect 2203 -1125 2215 -1073
rect 2267 -1125 2604 -1073
rect 2656 -1125 2668 -1073
rect 2720 -1125 2732 -1073
rect 2784 -1125 3840 -1073
rect 3892 -1125 3904 -1073
rect 3956 -1125 3968 -1073
rect 4020 -1125 4357 -1073
rect 4409 -1125 4421 -1073
rect 4473 -1125 4485 -1073
rect 4537 -1125 5624 -1073
rect 5676 -1125 5688 -1073
rect 5740 -1125 5752 -1073
rect 5804 -1125 6143 -1073
rect 6195 -1125 6207 -1073
rect 6259 -1125 6271 -1073
rect 6323 -1111 6637 -1073
rect 6693 -1111 6717 -1055
rect 6773 -1111 6797 -1055
rect 6853 -1111 6893 -1055
rect 6323 -1125 6893 -1111
rect -269 -1133 6893 -1125
rect 1314 -1173 5310 -1163
rect 1314 -1225 1321 -1173
rect 1373 -1225 1385 -1173
rect 1437 -1225 1449 -1173
rect 1501 -1225 1838 -1173
rect 1890 -1225 1902 -1173
rect 1954 -1225 1966 -1173
rect 2018 -1185 4606 -1173
rect 2018 -1225 3094 -1185
rect 1314 -1233 3094 -1225
rect 3054 -1241 3094 -1233
rect 3150 -1241 3174 -1185
rect 3230 -1241 3314 -1185
rect 3370 -1241 3394 -1185
rect 3450 -1241 3474 -1185
rect 3530 -1225 4606 -1185
rect 4658 -1225 4670 -1173
rect 4722 -1225 4734 -1173
rect 4786 -1225 5123 -1173
rect 5175 -1225 5187 -1173
rect 5239 -1225 5251 -1173
rect 5303 -1225 5310 -1173
rect 3530 -1233 5310 -1225
rect 3530 -1241 3570 -1233
rect 3054 -1263 3570 -1241
rect 879 -1537 1179 -1533
rect 5445 -1537 5745 -1533
rect 425 -1555 6199 -1537
rect 425 -1561 919 -1555
rect 425 -1613 551 -1561
rect 603 -1613 615 -1561
rect 667 -1613 679 -1561
rect 731 -1611 919 -1561
rect 975 -1611 999 -1555
rect 1055 -1611 1079 -1555
rect 1135 -1561 5489 -1555
rect 1135 -1611 2335 -1561
rect 731 -1613 2335 -1611
rect 2387 -1613 2399 -1561
rect 2451 -1613 2463 -1561
rect 2515 -1613 4109 -1561
rect 4161 -1613 4173 -1561
rect 4225 -1613 4237 -1561
rect 4289 -1611 5489 -1561
rect 5545 -1611 5569 -1555
rect 5625 -1611 5649 -1555
rect 5705 -1561 6199 -1555
rect 5705 -1611 5893 -1561
rect 4289 -1613 5893 -1611
rect 5945 -1613 5957 -1561
rect 6009 -1613 6021 -1561
rect 6073 -1613 6199 -1561
rect 425 -1633 6199 -1613
rect 1906 -1706 2206 -1687
rect 4418 -1706 4718 -1687
rect 425 -1709 6199 -1706
rect 425 -1718 1946 -1709
rect 425 -1770 551 -1718
rect 603 -1770 615 -1718
rect 667 -1770 679 -1718
rect 731 -1770 1217 -1718
rect 1269 -1770 1281 -1718
rect 1333 -1770 1345 -1718
rect 1397 -1770 1446 -1718
rect 1498 -1770 1510 -1718
rect 1562 -1770 1574 -1718
rect 1626 -1770 1684 -1718
rect 1736 -1770 1748 -1718
rect 1800 -1770 1812 -1718
rect 1864 -1765 1946 -1718
rect 2002 -1765 2026 -1709
rect 2082 -1765 2106 -1709
rect 2162 -1718 4462 -1709
rect 2162 -1765 2335 -1718
rect 1864 -1770 2335 -1765
rect 2387 -1770 2399 -1718
rect 2451 -1770 2463 -1718
rect 2515 -1770 4109 -1718
rect 4161 -1770 4173 -1718
rect 4225 -1770 4237 -1718
rect 4289 -1765 4462 -1718
rect 4518 -1765 4542 -1709
rect 4598 -1765 4622 -1709
rect 4678 -1718 6199 -1709
rect 4678 -1765 4760 -1718
rect 4289 -1770 4760 -1765
rect 4812 -1770 4824 -1718
rect 4876 -1770 4888 -1718
rect 4940 -1770 4998 -1718
rect 5050 -1770 5062 -1718
rect 5114 -1770 5126 -1718
rect 5178 -1770 5227 -1718
rect 5279 -1770 5291 -1718
rect 5343 -1770 5355 -1718
rect 5407 -1770 5893 -1718
rect 5945 -1770 5957 -1718
rect 6009 -1770 6021 -1718
rect 6073 -1770 6199 -1718
rect 425 -1787 6199 -1770
rect 425 -1870 6199 -1850
rect 425 -1922 551 -1870
rect 603 -1922 615 -1870
rect 667 -1922 679 -1870
rect 731 -1872 2335 -1870
rect 731 -1922 1946 -1872
rect 425 -1928 1946 -1922
rect 2002 -1928 2026 -1872
rect 2082 -1928 2106 -1872
rect 2162 -1922 2335 -1872
rect 2387 -1922 2399 -1870
rect 2451 -1922 2463 -1870
rect 2515 -1922 4109 -1870
rect 4161 -1922 4173 -1870
rect 4225 -1922 4237 -1870
rect 4289 -1872 5893 -1870
rect 4289 -1922 4462 -1872
rect 2162 -1928 4462 -1922
rect 4518 -1928 4542 -1872
rect 4598 -1928 4622 -1872
rect 4678 -1922 5893 -1872
rect 5945 -1922 5957 -1870
rect 6009 -1922 6021 -1870
rect 6073 -1922 6199 -1870
rect 4678 -1928 6199 -1922
rect 425 -1946 6199 -1928
rect 1906 -1950 2206 -1946
rect 4418 -1950 4718 -1946
rect 2622 -2227 2922 -2205
rect 2622 -2235 2662 -2227
rect 550 -2245 2662 -2235
rect 550 -2297 560 -2245
rect 612 -2297 624 -2245
rect 676 -2297 688 -2245
rect 740 -2297 2344 -2245
rect 2396 -2297 2408 -2245
rect 2460 -2297 2472 -2245
rect 2524 -2283 2662 -2245
rect 2718 -2283 2742 -2227
rect 2798 -2283 2822 -2227
rect 2878 -2235 2922 -2227
rect 3702 -2227 4002 -2205
rect 3702 -2235 3746 -2227
rect 2878 -2283 3746 -2235
rect 3802 -2283 3826 -2227
rect 3882 -2283 3906 -2227
rect 3962 -2235 4002 -2227
rect 3962 -2245 6074 -2235
rect 3962 -2283 4100 -2245
rect 2524 -2297 4100 -2283
rect 4152 -2297 4164 -2245
rect 4216 -2297 4228 -2245
rect 4280 -2297 5884 -2245
rect 5936 -2297 5948 -2245
rect 6000 -2297 6012 -2245
rect 6064 -2297 6074 -2245
rect 550 -2305 6074 -2297
rect 163 -2327 463 -2305
rect 163 -2383 203 -2327
rect 259 -2383 283 -2327
rect 339 -2383 363 -2327
rect 419 -2334 463 -2327
rect 6161 -2327 6461 -2305
rect 6161 -2334 6205 -2327
rect 419 -2344 1770 -2334
rect 419 -2383 1064 -2344
rect 163 -2396 1064 -2383
rect 1116 -2396 1128 -2344
rect 1180 -2396 1192 -2344
rect 1244 -2396 1581 -2344
rect 1633 -2396 1645 -2344
rect 1697 -2396 1709 -2344
rect 1761 -2396 1770 -2344
rect 163 -2405 1770 -2396
rect 4854 -2344 6205 -2334
rect 4854 -2396 4863 -2344
rect 4915 -2396 4927 -2344
rect 4979 -2396 4991 -2344
rect 5043 -2396 5380 -2344
rect 5432 -2396 5444 -2344
rect 5496 -2396 5508 -2344
rect 5560 -2383 6205 -2344
rect 6261 -2383 6285 -2327
rect 6341 -2383 6365 -2327
rect 6421 -2383 6461 -2327
rect 5560 -2396 6461 -2383
rect 4854 -2405 6461 -2396
rect 3054 -2438 3570 -2416
rect 3054 -2446 3094 -2438
rect 369 -2456 3094 -2446
rect 369 -2508 376 -2456
rect 428 -2508 440 -2456
rect 492 -2508 504 -2456
rect 556 -2508 742 -2456
rect 794 -2508 806 -2456
rect 858 -2508 870 -2456
rect 922 -2508 2160 -2456
rect 2212 -2508 2224 -2456
rect 2276 -2508 2288 -2456
rect 2340 -2508 2526 -2456
rect 2578 -2508 2590 -2456
rect 2642 -2508 2654 -2456
rect 2706 -2494 3094 -2456
rect 3150 -2494 3174 -2438
rect 3230 -2494 3254 -2438
rect 3310 -2494 3394 -2438
rect 3450 -2494 3474 -2438
rect 3530 -2446 3570 -2438
rect 3530 -2456 6255 -2446
rect 3530 -2494 3918 -2456
rect 2706 -2508 3918 -2494
rect 3970 -2508 3982 -2456
rect 4034 -2508 4046 -2456
rect 4098 -2508 4284 -2456
rect 4336 -2508 4348 -2456
rect 4400 -2508 4412 -2456
rect 4464 -2508 5702 -2456
rect 5754 -2508 5766 -2456
rect 5818 -2508 5830 -2456
rect 5882 -2508 6068 -2456
rect 6120 -2508 6132 -2456
rect 6184 -2508 6196 -2456
rect 6248 -2508 6255 -2456
rect -269 -2537 31 -2515
rect 369 -2516 6255 -2508
rect -269 -2593 -229 -2537
rect -173 -2593 -149 -2537
rect -93 -2593 -69 -2537
rect -13 -2545 31 -2537
rect 6593 -2537 6893 -2515
rect 6593 -2545 6637 -2537
rect -13 -2555 6637 -2545
rect -13 -2593 1321 -2555
rect -269 -2607 1321 -2593
rect 1373 -2607 1385 -2555
rect 1437 -2607 1449 -2555
rect 1501 -2607 1838 -2555
rect 1890 -2607 1902 -2555
rect 1954 -2607 1966 -2555
rect 2018 -2607 4606 -2555
rect 4658 -2607 4670 -2555
rect 4722 -2607 4734 -2555
rect 4786 -2607 5123 -2555
rect 5175 -2607 5187 -2555
rect 5239 -2607 5251 -2555
rect 5303 -2593 6637 -2555
rect 6693 -2593 6717 -2537
rect 6773 -2593 6797 -2537
rect 6853 -2593 6893 -2537
rect 5303 -2607 6893 -2593
rect -269 -2615 6893 -2607
<< via2 >>
rect -229 482 -173 538
rect -149 482 -93 538
rect -69 482 -13 538
rect 6637 482 6693 538
rect 6717 482 6773 538
rect 6797 482 6853 538
rect 3094 375 3150 431
rect 3174 375 3230 431
rect 3254 375 3310 431
rect 3394 375 3450 431
rect 3474 375 3530 431
rect 203 240 259 296
rect 283 240 339 296
rect 363 240 419 296
rect 6205 240 6261 296
rect 6285 240 6341 296
rect 6365 240 6421 296
rect 2662 141 2718 197
rect 2742 141 2798 197
rect 2822 141 2878 197
rect 3746 141 3802 197
rect 3826 141 3882 197
rect 3906 141 3962 197
rect 1946 -214 2002 -158
rect 2026 -214 2082 -158
rect 2106 -214 2162 -158
rect 4462 -214 4518 -158
rect 4542 -214 4598 -158
rect 4622 -214 4678 -158
rect 1946 -377 2002 -321
rect 2026 -377 2082 -321
rect 2106 -377 2162 -321
rect 4462 -377 4518 -321
rect 4542 -377 4598 -321
rect 4622 -377 4678 -321
rect 919 -531 975 -475
rect 999 -531 1055 -475
rect 1079 -531 1135 -475
rect 5489 -531 5545 -475
rect 5569 -531 5625 -475
rect 5649 -531 5705 -475
rect 203 -847 259 -791
rect 283 -847 339 -791
rect 363 -847 419 -791
rect 6205 -847 6261 -791
rect 6285 -847 6341 -791
rect 6365 -847 6421 -791
rect 2662 -1000 2718 -944
rect 2742 -1000 2798 -944
rect 2822 -1000 2878 -944
rect 3746 -1000 3802 -944
rect 3826 -1000 3882 -944
rect 3906 -1000 3962 -944
rect -229 -1111 -173 -1055
rect -149 -1111 -93 -1055
rect -69 -1111 -13 -1055
rect 6637 -1111 6693 -1055
rect 6717 -1111 6773 -1055
rect 6797 -1111 6853 -1055
rect 3094 -1241 3150 -1185
rect 3174 -1241 3230 -1185
rect 3314 -1241 3370 -1185
rect 3394 -1241 3450 -1185
rect 3474 -1241 3530 -1185
rect 919 -1611 975 -1555
rect 999 -1611 1055 -1555
rect 1079 -1611 1135 -1555
rect 5489 -1611 5545 -1555
rect 5569 -1611 5625 -1555
rect 5649 -1611 5705 -1555
rect 1946 -1765 2002 -1709
rect 2026 -1765 2082 -1709
rect 2106 -1765 2162 -1709
rect 4462 -1765 4518 -1709
rect 4542 -1765 4598 -1709
rect 4622 -1765 4678 -1709
rect 1946 -1928 2002 -1872
rect 2026 -1928 2082 -1872
rect 2106 -1928 2162 -1872
rect 4462 -1928 4518 -1872
rect 4542 -1928 4598 -1872
rect 4622 -1928 4678 -1872
rect 2662 -2283 2718 -2227
rect 2742 -2283 2798 -2227
rect 2822 -2283 2878 -2227
rect 3746 -2283 3802 -2227
rect 3826 -2283 3882 -2227
rect 3906 -2283 3962 -2227
rect 203 -2383 259 -2327
rect 283 -2383 339 -2327
rect 363 -2383 419 -2327
rect 6205 -2383 6261 -2327
rect 6285 -2383 6341 -2327
rect 6365 -2383 6421 -2327
rect 3094 -2494 3150 -2438
rect 3174 -2494 3230 -2438
rect 3254 -2494 3310 -2438
rect 3394 -2494 3450 -2438
rect 3474 -2494 3530 -2438
rect -229 -2593 -173 -2537
rect -149 -2593 -93 -2537
rect -69 -2593 -13 -2537
rect 6637 -2593 6693 -2537
rect 6717 -2593 6773 -2537
rect 6797 -2593 6853 -2537
<< metal3 >>
rect -269 538 31 560
rect -269 482 -229 538
rect -173 482 -149 538
rect -93 482 -69 538
rect -13 482 31 538
rect -269 -1055 31 482
rect 6593 538 6893 560
rect 6593 482 6637 538
rect 6693 482 6717 538
rect 6773 482 6797 538
rect 6853 482 6893 538
rect 3054 431 3570 453
rect 3054 375 3094 431
rect 3150 375 3174 431
rect 3230 375 3254 431
rect 3310 375 3394 431
rect 3450 375 3474 431
rect 3530 375 3570 431
rect -269 -1111 -229 -1055
rect -173 -1111 -149 -1055
rect -93 -1111 -69 -1055
rect -13 -1111 31 -1055
rect -269 -2537 31 -1111
rect 163 296 463 318
rect 163 240 203 296
rect 259 240 283 296
rect 339 240 363 296
rect 419 240 463 296
rect 163 -791 463 240
rect 2622 197 2922 219
rect 2622 141 2662 197
rect 2718 141 2742 197
rect 2798 141 2822 197
rect 2878 141 2922 197
rect 1906 -158 2206 -136
rect 1906 -214 1946 -158
rect 2002 -214 2026 -158
rect 2082 -214 2106 -158
rect 2162 -214 2206 -158
rect 1906 -321 2206 -214
rect 1906 -377 1946 -321
rect 2002 -377 2026 -321
rect 2082 -377 2106 -321
rect 2162 -377 2206 -321
rect 163 -847 203 -791
rect 259 -847 283 -791
rect 339 -847 363 -791
rect 419 -847 463 -791
rect 163 -2327 463 -847
rect 879 -475 1180 -453
rect 879 -531 919 -475
rect 975 -531 999 -475
rect 1055 -531 1079 -475
rect 1135 -531 1180 -475
rect 879 -1555 1180 -531
rect 879 -1611 919 -1555
rect 975 -1611 999 -1555
rect 1055 -1611 1079 -1555
rect 1135 -1611 1180 -1555
rect 879 -1633 1180 -1611
rect 1906 -1709 2206 -377
rect 1906 -1765 1946 -1709
rect 2002 -1765 2026 -1709
rect 2082 -1765 2106 -1709
rect 2162 -1765 2206 -1709
rect 1906 -1872 2206 -1765
rect 1906 -1928 1946 -1872
rect 2002 -1928 2026 -1872
rect 2082 -1928 2106 -1872
rect 2162 -1928 2206 -1872
rect 1906 -1950 2206 -1928
rect 2622 -944 2922 141
rect 2622 -1000 2662 -944
rect 2718 -1000 2742 -944
rect 2798 -1000 2822 -944
rect 2878 -1000 2922 -944
rect 2622 -2227 2922 -1000
rect 2622 -2283 2662 -2227
rect 2718 -2283 2742 -2227
rect 2798 -2283 2822 -2227
rect 2878 -2283 2922 -2227
rect 2622 -2305 2922 -2283
rect 3054 -1185 3570 375
rect 6161 296 6461 318
rect 6161 240 6205 296
rect 6261 240 6285 296
rect 6341 240 6365 296
rect 6421 240 6461 296
rect 3054 -1241 3094 -1185
rect 3150 -1241 3174 -1185
rect 3230 -1241 3314 -1185
rect 3370 -1241 3394 -1185
rect 3450 -1241 3474 -1185
rect 3530 -1241 3570 -1185
rect 163 -2383 203 -2327
rect 259 -2383 283 -2327
rect 339 -2383 363 -2327
rect 419 -2383 463 -2327
rect 163 -2405 463 -2383
rect 3054 -2438 3570 -1241
rect 3702 197 4002 219
rect 3702 141 3746 197
rect 3802 141 3826 197
rect 3882 141 3906 197
rect 3962 141 4002 197
rect 3702 -944 4002 141
rect 3702 -1000 3746 -944
rect 3802 -1000 3826 -944
rect 3882 -1000 3906 -944
rect 3962 -1000 4002 -944
rect 3702 -2227 4002 -1000
rect 4418 -158 4718 -136
rect 4418 -214 4462 -158
rect 4518 -214 4542 -158
rect 4598 -214 4622 -158
rect 4678 -214 4718 -158
rect 4418 -321 4718 -214
rect 4418 -377 4462 -321
rect 4518 -377 4542 -321
rect 4598 -377 4622 -321
rect 4678 -377 4718 -321
rect 4418 -1709 4718 -377
rect 5444 -475 5745 -453
rect 5444 -531 5489 -475
rect 5545 -531 5569 -475
rect 5625 -531 5649 -475
rect 5705 -531 5745 -475
rect 5444 -1555 5745 -531
rect 5444 -1611 5489 -1555
rect 5545 -1611 5569 -1555
rect 5625 -1611 5649 -1555
rect 5705 -1611 5745 -1555
rect 5444 -1633 5745 -1611
rect 6161 -791 6461 240
rect 6161 -847 6205 -791
rect 6261 -847 6285 -791
rect 6341 -847 6365 -791
rect 6421 -847 6461 -791
rect 4418 -1765 4462 -1709
rect 4518 -1765 4542 -1709
rect 4598 -1765 4622 -1709
rect 4678 -1765 4718 -1709
rect 4418 -1872 4718 -1765
rect 4418 -1928 4462 -1872
rect 4518 -1928 4542 -1872
rect 4598 -1928 4622 -1872
rect 4678 -1928 4718 -1872
rect 4418 -1950 4718 -1928
rect 3702 -2283 3746 -2227
rect 3802 -2283 3826 -2227
rect 3882 -2283 3906 -2227
rect 3962 -2283 4002 -2227
rect 3702 -2305 4002 -2283
rect 6161 -2327 6461 -847
rect 6161 -2383 6205 -2327
rect 6261 -2383 6285 -2327
rect 6341 -2383 6365 -2327
rect 6421 -2383 6461 -2327
rect 6161 -2405 6461 -2383
rect 6593 -1055 6893 482
rect 6593 -1111 6637 -1055
rect 6693 -1111 6717 -1055
rect 6773 -1111 6797 -1055
rect 6853 -1111 6893 -1055
rect 3054 -2494 3094 -2438
rect 3150 -2494 3174 -2438
rect 3230 -2494 3254 -2438
rect 3310 -2494 3394 -2438
rect 3450 -2494 3474 -2438
rect 3530 -2494 3570 -2438
rect 3054 -2516 3570 -2494
rect -269 -2593 -229 -2537
rect -173 -2593 -149 -2537
rect -93 -2593 -69 -2537
rect -13 -2593 31 -2537
rect -269 -2615 31 -2593
rect 6593 -2537 6893 -1111
rect 6593 -2593 6637 -2537
rect 6693 -2593 6717 -2537
rect 6773 -2593 6797 -2537
rect 6853 -2593 6893 -2537
rect 6593 -2615 6893 -2593
<< end >>
