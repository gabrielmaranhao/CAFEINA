magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< pwell >>
rect 1048 -158 3305 562
rect 1048 -358 1134 -158
rect 3219 -358 3305 -158
rect 1048 -754 3305 -358
<< nmos >>
rect 1238 165 1438 365
rect 1689 165 1889 365
rect 1947 165 2147 365
rect 2205 165 2405 365
rect 2463 165 2663 365
rect 2915 165 3115 365
rect 1238 -132 1438 68
rect 1689 -132 1889 68
rect 1947 -132 2147 68
rect 2205 -132 2405 68
rect 2463 -132 2663 68
rect 2915 -132 3115 68
rect 1238 -584 1438 -384
rect 1689 -584 1889 -384
rect 1947 -584 2147 -384
rect 2205 -584 2405 -384
rect 2463 -584 2663 -384
rect 2915 -584 3115 -384
<< ndiff >>
rect 1180 350 1238 365
rect 1180 316 1192 350
rect 1226 316 1238 350
rect 1180 282 1238 316
rect 1180 248 1192 282
rect 1226 248 1238 282
rect 1180 214 1238 248
rect 1180 180 1192 214
rect 1226 180 1238 214
rect 1180 165 1238 180
rect 1438 350 1496 365
rect 1438 316 1450 350
rect 1484 316 1496 350
rect 1438 282 1496 316
rect 1438 248 1450 282
rect 1484 248 1496 282
rect 1438 214 1496 248
rect 1438 180 1450 214
rect 1484 180 1496 214
rect 1438 165 1496 180
rect 1631 350 1689 365
rect 1631 316 1643 350
rect 1677 316 1689 350
rect 1631 282 1689 316
rect 1631 248 1643 282
rect 1677 248 1689 282
rect 1631 214 1689 248
rect 1631 180 1643 214
rect 1677 180 1689 214
rect 1631 165 1689 180
rect 1889 350 1947 365
rect 1889 316 1901 350
rect 1935 316 1947 350
rect 1889 282 1947 316
rect 1889 248 1901 282
rect 1935 248 1947 282
rect 1889 214 1947 248
rect 1889 180 1901 214
rect 1935 180 1947 214
rect 1889 165 1947 180
rect 2147 350 2205 365
rect 2147 316 2159 350
rect 2193 316 2205 350
rect 2147 282 2205 316
rect 2147 248 2159 282
rect 2193 248 2205 282
rect 2147 214 2205 248
rect 2147 180 2159 214
rect 2193 180 2205 214
rect 2147 165 2205 180
rect 2405 350 2463 365
rect 2405 316 2417 350
rect 2451 316 2463 350
rect 2405 282 2463 316
rect 2405 248 2417 282
rect 2451 248 2463 282
rect 2405 214 2463 248
rect 2405 180 2417 214
rect 2451 180 2463 214
rect 2405 165 2463 180
rect 2663 350 2721 365
rect 2663 316 2675 350
rect 2709 316 2721 350
rect 2663 282 2721 316
rect 2663 248 2675 282
rect 2709 248 2721 282
rect 2663 214 2721 248
rect 2663 180 2675 214
rect 2709 180 2721 214
rect 2663 165 2721 180
rect 2857 350 2915 365
rect 2857 316 2869 350
rect 2903 316 2915 350
rect 2857 282 2915 316
rect 2857 248 2869 282
rect 2903 248 2915 282
rect 2857 214 2915 248
rect 2857 180 2869 214
rect 2903 180 2915 214
rect 2857 165 2915 180
rect 3115 350 3173 365
rect 3115 316 3127 350
rect 3161 316 3173 350
rect 3115 282 3173 316
rect 3115 248 3127 282
rect 3161 248 3173 282
rect 3115 214 3173 248
rect 3115 180 3127 214
rect 3161 180 3173 214
rect 3115 165 3173 180
rect 1180 53 1238 68
rect 1180 19 1192 53
rect 1226 19 1238 53
rect 1180 -15 1238 19
rect 1180 -49 1192 -15
rect 1226 -49 1238 -15
rect 1180 -83 1238 -49
rect 1180 -117 1192 -83
rect 1226 -117 1238 -83
rect 1180 -132 1238 -117
rect 1438 53 1496 68
rect 1438 19 1450 53
rect 1484 19 1496 53
rect 1438 -15 1496 19
rect 1438 -49 1450 -15
rect 1484 -49 1496 -15
rect 1438 -83 1496 -49
rect 1438 -117 1450 -83
rect 1484 -117 1496 -83
rect 1438 -132 1496 -117
rect 1631 53 1689 68
rect 1631 19 1643 53
rect 1677 19 1689 53
rect 1631 -15 1689 19
rect 1631 -49 1643 -15
rect 1677 -49 1689 -15
rect 1631 -83 1689 -49
rect 1631 -117 1643 -83
rect 1677 -117 1689 -83
rect 1631 -132 1689 -117
rect 1889 53 1947 68
rect 1889 19 1901 53
rect 1935 19 1947 53
rect 1889 -15 1947 19
rect 1889 -49 1901 -15
rect 1935 -49 1947 -15
rect 1889 -83 1947 -49
rect 1889 -117 1901 -83
rect 1935 -117 1947 -83
rect 1889 -132 1947 -117
rect 2147 53 2205 68
rect 2147 19 2159 53
rect 2193 19 2205 53
rect 2147 -15 2205 19
rect 2147 -49 2159 -15
rect 2193 -49 2205 -15
rect 2147 -83 2205 -49
rect 2147 -117 2159 -83
rect 2193 -117 2205 -83
rect 2147 -132 2205 -117
rect 2405 53 2463 68
rect 2405 19 2417 53
rect 2451 19 2463 53
rect 2405 -15 2463 19
rect 2405 -49 2417 -15
rect 2451 -49 2463 -15
rect 2405 -83 2463 -49
rect 2405 -117 2417 -83
rect 2451 -117 2463 -83
rect 2405 -132 2463 -117
rect 2663 53 2721 68
rect 2663 19 2675 53
rect 2709 19 2721 53
rect 2663 -15 2721 19
rect 2663 -49 2675 -15
rect 2709 -49 2721 -15
rect 2663 -83 2721 -49
rect 2663 -117 2675 -83
rect 2709 -117 2721 -83
rect 2663 -132 2721 -117
rect 2857 53 2915 68
rect 2857 19 2869 53
rect 2903 19 2915 53
rect 2857 -15 2915 19
rect 2857 -49 2869 -15
rect 2903 -49 2915 -15
rect 2857 -83 2915 -49
rect 2857 -117 2869 -83
rect 2903 -117 2915 -83
rect 2857 -132 2915 -117
rect 3115 53 3173 68
rect 3115 19 3127 53
rect 3161 19 3173 53
rect 3115 -15 3173 19
rect 3115 -49 3127 -15
rect 3161 -49 3173 -15
rect 3115 -83 3173 -49
rect 3115 -117 3127 -83
rect 3161 -117 3173 -83
rect 3115 -132 3173 -117
rect 1180 -399 1238 -384
rect 1180 -433 1192 -399
rect 1226 -433 1238 -399
rect 1180 -467 1238 -433
rect 1180 -501 1192 -467
rect 1226 -501 1238 -467
rect 1180 -535 1238 -501
rect 1180 -569 1192 -535
rect 1226 -569 1238 -535
rect 1180 -584 1238 -569
rect 1438 -399 1496 -384
rect 1438 -433 1450 -399
rect 1484 -433 1496 -399
rect 1438 -467 1496 -433
rect 1438 -501 1450 -467
rect 1484 -501 1496 -467
rect 1438 -535 1496 -501
rect 1438 -569 1450 -535
rect 1484 -569 1496 -535
rect 1438 -584 1496 -569
rect 1631 -399 1689 -384
rect 1631 -433 1643 -399
rect 1677 -433 1689 -399
rect 1631 -467 1689 -433
rect 1631 -501 1643 -467
rect 1677 -501 1689 -467
rect 1631 -535 1689 -501
rect 1631 -569 1643 -535
rect 1677 -569 1689 -535
rect 1631 -584 1689 -569
rect 1889 -399 1947 -384
rect 1889 -433 1901 -399
rect 1935 -433 1947 -399
rect 1889 -467 1947 -433
rect 1889 -501 1901 -467
rect 1935 -501 1947 -467
rect 1889 -535 1947 -501
rect 1889 -569 1901 -535
rect 1935 -569 1947 -535
rect 1889 -584 1947 -569
rect 2147 -399 2205 -384
rect 2147 -433 2159 -399
rect 2193 -433 2205 -399
rect 2147 -467 2205 -433
rect 2147 -501 2159 -467
rect 2193 -501 2205 -467
rect 2147 -535 2205 -501
rect 2147 -569 2159 -535
rect 2193 -569 2205 -535
rect 2147 -584 2205 -569
rect 2405 -399 2463 -384
rect 2405 -433 2417 -399
rect 2451 -433 2463 -399
rect 2405 -467 2463 -433
rect 2405 -501 2417 -467
rect 2451 -501 2463 -467
rect 2405 -535 2463 -501
rect 2405 -569 2417 -535
rect 2451 -569 2463 -535
rect 2405 -584 2463 -569
rect 2663 -399 2721 -384
rect 2663 -433 2675 -399
rect 2709 -433 2721 -399
rect 2663 -467 2721 -433
rect 2663 -501 2675 -467
rect 2709 -501 2721 -467
rect 2663 -535 2721 -501
rect 2663 -569 2675 -535
rect 2709 -569 2721 -535
rect 2663 -584 2721 -569
rect 2857 -399 2915 -384
rect 2857 -433 2869 -399
rect 2903 -433 2915 -399
rect 2857 -467 2915 -433
rect 2857 -501 2869 -467
rect 2903 -501 2915 -467
rect 2857 -535 2915 -501
rect 2857 -569 2869 -535
rect 2903 -569 2915 -535
rect 2857 -584 2915 -569
rect 3115 -399 3173 -384
rect 3115 -433 3127 -399
rect 3161 -433 3173 -399
rect 3115 -467 3173 -433
rect 3115 -501 3127 -467
rect 3161 -501 3173 -467
rect 3115 -535 3173 -501
rect 3115 -569 3127 -535
rect 3161 -569 3173 -535
rect 3115 -584 3173 -569
<< ndiffc >>
rect 1192 316 1226 350
rect 1192 248 1226 282
rect 1192 180 1226 214
rect 1450 316 1484 350
rect 1450 248 1484 282
rect 1450 180 1484 214
rect 1643 316 1677 350
rect 1643 248 1677 282
rect 1643 180 1677 214
rect 1901 316 1935 350
rect 1901 248 1935 282
rect 1901 180 1935 214
rect 2159 316 2193 350
rect 2159 248 2193 282
rect 2159 180 2193 214
rect 2417 316 2451 350
rect 2417 248 2451 282
rect 2417 180 2451 214
rect 2675 316 2709 350
rect 2675 248 2709 282
rect 2675 180 2709 214
rect 2869 316 2903 350
rect 2869 248 2903 282
rect 2869 180 2903 214
rect 3127 316 3161 350
rect 3127 248 3161 282
rect 3127 180 3161 214
rect 1192 19 1226 53
rect 1192 -49 1226 -15
rect 1192 -117 1226 -83
rect 1450 19 1484 53
rect 1450 -49 1484 -15
rect 1450 -117 1484 -83
rect 1643 19 1677 53
rect 1643 -49 1677 -15
rect 1643 -117 1677 -83
rect 1901 19 1935 53
rect 1901 -49 1935 -15
rect 1901 -117 1935 -83
rect 2159 19 2193 53
rect 2159 -49 2193 -15
rect 2159 -117 2193 -83
rect 2417 19 2451 53
rect 2417 -49 2451 -15
rect 2417 -117 2451 -83
rect 2675 19 2709 53
rect 2675 -49 2709 -15
rect 2675 -117 2709 -83
rect 2869 19 2903 53
rect 2869 -49 2903 -15
rect 2869 -117 2903 -83
rect 3127 19 3161 53
rect 3127 -49 3161 -15
rect 3127 -117 3161 -83
rect 1192 -433 1226 -399
rect 1192 -501 1226 -467
rect 1192 -569 1226 -535
rect 1450 -433 1484 -399
rect 1450 -501 1484 -467
rect 1450 -569 1484 -535
rect 1643 -433 1677 -399
rect 1643 -501 1677 -467
rect 1643 -569 1677 -535
rect 1901 -433 1935 -399
rect 1901 -501 1935 -467
rect 1901 -569 1935 -535
rect 2159 -433 2193 -399
rect 2159 -501 2193 -467
rect 2159 -569 2193 -535
rect 2417 -433 2451 -399
rect 2417 -501 2451 -467
rect 2417 -569 2451 -535
rect 2675 -433 2709 -399
rect 2675 -501 2709 -467
rect 2675 -569 2709 -535
rect 2869 -433 2903 -399
rect 2869 -501 2903 -467
rect 2869 -569 2903 -535
rect 3127 -433 3161 -399
rect 3127 -501 3161 -467
rect 3127 -569 3161 -535
<< psubdiff >>
rect 1074 502 1259 536
rect 1293 502 1327 536
rect 1361 502 1395 536
rect 1429 502 1463 536
rect 1497 502 1531 536
rect 1565 502 1599 536
rect 1633 502 1667 536
rect 1701 502 1735 536
rect 1769 502 1803 536
rect 1837 502 1871 536
rect 1905 502 1939 536
rect 1973 502 2007 536
rect 2041 502 2075 536
rect 2109 502 2143 536
rect 2177 502 2211 536
rect 2245 502 2279 536
rect 2313 502 2347 536
rect 2381 502 2415 536
rect 2449 502 2483 536
rect 2517 502 2551 536
rect 2585 502 2619 536
rect 2653 502 2687 536
rect 2721 502 2755 536
rect 2789 502 2823 536
rect 2857 502 2891 536
rect 2925 502 2959 536
rect 2993 502 3027 536
rect 3061 502 3095 536
rect 3129 502 3279 536
rect 1074 351 1108 502
rect 1074 283 1108 317
rect 1074 215 1108 249
rect 1074 147 1108 181
rect 3245 351 3279 502
rect 3245 283 3279 317
rect 3245 215 3279 249
rect 3245 147 3279 181
rect 1074 54 1108 113
rect 1074 -14 1108 20
rect 1074 -82 1108 -48
rect 1074 -150 1108 -116
rect 3245 54 3279 113
rect 3245 -14 3279 20
rect 3245 -82 3279 -48
rect 1074 -218 1108 -184
rect 3245 -150 3279 -116
rect 3245 -218 3279 -184
rect 1074 -286 1108 -252
rect 3245 -286 3279 -252
rect 1074 -354 1108 -320
rect 3245 -354 3279 -320
rect 1074 -422 1108 -388
rect 1074 -490 1108 -456
rect 1074 -558 1108 -524
rect 3245 -422 3279 -388
rect 3245 -490 3279 -456
rect 3245 -558 3279 -524
rect 1074 -694 1108 -592
rect 3245 -694 3279 -592
rect 1074 -728 1259 -694
rect 1293 -728 1327 -694
rect 1361 -728 1395 -694
rect 1429 -728 1463 -694
rect 1497 -728 1531 -694
rect 1565 -728 1599 -694
rect 1633 -728 1667 -694
rect 1701 -728 1735 -694
rect 1769 -728 1803 -694
rect 1837 -728 1871 -694
rect 1905 -728 1939 -694
rect 1973 -728 2007 -694
rect 2041 -728 2075 -694
rect 2109 -728 2143 -694
rect 2177 -728 2211 -694
rect 2245 -728 2279 -694
rect 2313 -728 2347 -694
rect 2381 -728 2415 -694
rect 2449 -728 2483 -694
rect 2517 -728 2551 -694
rect 2585 -728 2619 -694
rect 2653 -728 2687 -694
rect 2721 -728 2755 -694
rect 2789 -728 2823 -694
rect 2857 -728 2891 -694
rect 2925 -728 2959 -694
rect 2993 -728 3027 -694
rect 3061 -728 3095 -694
rect 3129 -728 3279 -694
<< psubdiffcont >>
rect 1259 502 1293 536
rect 1327 502 1361 536
rect 1395 502 1429 536
rect 1463 502 1497 536
rect 1531 502 1565 536
rect 1599 502 1633 536
rect 1667 502 1701 536
rect 1735 502 1769 536
rect 1803 502 1837 536
rect 1871 502 1905 536
rect 1939 502 1973 536
rect 2007 502 2041 536
rect 2075 502 2109 536
rect 2143 502 2177 536
rect 2211 502 2245 536
rect 2279 502 2313 536
rect 2347 502 2381 536
rect 2415 502 2449 536
rect 2483 502 2517 536
rect 2551 502 2585 536
rect 2619 502 2653 536
rect 2687 502 2721 536
rect 2755 502 2789 536
rect 2823 502 2857 536
rect 2891 502 2925 536
rect 2959 502 2993 536
rect 3027 502 3061 536
rect 3095 502 3129 536
rect 1074 317 1108 351
rect 1074 249 1108 283
rect 1074 181 1108 215
rect 3245 317 3279 351
rect 3245 249 3279 283
rect 3245 181 3279 215
rect 1074 113 1108 147
rect 3245 113 3279 147
rect 1074 20 1108 54
rect 1074 -48 1108 -14
rect 1074 -116 1108 -82
rect 3245 20 3279 54
rect 3245 -48 3279 -14
rect 3245 -116 3279 -82
rect 1074 -184 1108 -150
rect 1074 -252 1108 -218
rect 3245 -184 3279 -150
rect 1074 -320 1108 -286
rect 3245 -252 3279 -218
rect 1074 -388 1108 -354
rect 3245 -320 3279 -286
rect 1074 -456 1108 -422
rect 1074 -524 1108 -490
rect 1074 -592 1108 -558
rect 3245 -388 3279 -354
rect 3245 -456 3279 -422
rect 3245 -524 3279 -490
rect 3245 -592 3279 -558
rect 1259 -728 1293 -694
rect 1327 -728 1361 -694
rect 1395 -728 1429 -694
rect 1463 -728 1497 -694
rect 1531 -728 1565 -694
rect 1599 -728 1633 -694
rect 1667 -728 1701 -694
rect 1735 -728 1769 -694
rect 1803 -728 1837 -694
rect 1871 -728 1905 -694
rect 1939 -728 1973 -694
rect 2007 -728 2041 -694
rect 2075 -728 2109 -694
rect 2143 -728 2177 -694
rect 2211 -728 2245 -694
rect 2279 -728 2313 -694
rect 2347 -728 2381 -694
rect 2415 -728 2449 -694
rect 2483 -728 2517 -694
rect 2551 -728 2585 -694
rect 2619 -728 2653 -694
rect 2687 -728 2721 -694
rect 2755 -728 2789 -694
rect 2823 -728 2857 -694
rect 2891 -728 2925 -694
rect 2959 -728 2993 -694
rect 3027 -728 3061 -694
rect 3095 -728 3129 -694
<< poly >>
rect 1238 437 1438 453
rect 1238 403 1287 437
rect 1321 403 1355 437
rect 1389 403 1438 437
rect 1238 365 1438 403
rect 1689 437 1889 453
rect 1689 403 1738 437
rect 1772 403 1806 437
rect 1840 403 1889 437
rect 1689 365 1889 403
rect 1947 437 2147 453
rect 1947 403 1996 437
rect 2030 403 2064 437
rect 2098 403 2147 437
rect 1947 365 2147 403
rect 2205 437 2405 453
rect 2205 403 2254 437
rect 2288 403 2322 437
rect 2356 403 2405 437
rect 2205 365 2405 403
rect 2463 437 2663 453
rect 2463 403 2512 437
rect 2546 403 2580 437
rect 2614 403 2663 437
rect 2463 365 2663 403
rect 2915 437 3115 453
rect 2915 403 2964 437
rect 2998 403 3032 437
rect 3066 403 3115 437
rect 2915 365 3115 403
rect 1238 139 1438 165
rect 1689 139 1889 165
rect 1947 139 2147 165
rect 2205 139 2405 165
rect 2463 139 2663 165
rect 2915 139 3115 165
rect 1238 68 1438 94
rect 1689 68 1889 94
rect 1947 68 2147 94
rect 2205 68 2405 94
rect 2463 68 2663 94
rect 2915 68 3115 94
rect 1238 -170 1438 -132
rect 1238 -204 1287 -170
rect 1321 -204 1355 -170
rect 1389 -204 1438 -170
rect 1238 -220 1438 -204
rect 1689 -170 1889 -132
rect 1689 -204 1738 -170
rect 1772 -204 1806 -170
rect 1840 -204 1889 -170
rect 1689 -220 1889 -204
rect 1947 -170 2147 -132
rect 1947 -204 1996 -170
rect 2030 -204 2064 -170
rect 2098 -204 2147 -170
rect 1947 -220 2147 -204
rect 2205 -170 2405 -132
rect 2205 -204 2254 -170
rect 2288 -204 2322 -170
rect 2356 -204 2405 -170
rect 2205 -220 2405 -204
rect 2463 -170 2663 -132
rect 2463 -204 2512 -170
rect 2546 -204 2580 -170
rect 2614 -204 2663 -170
rect 2463 -220 2663 -204
rect 2915 -170 3115 -132
rect 2915 -204 2964 -170
rect 2998 -204 3032 -170
rect 3066 -204 3115 -170
rect 2915 -220 3115 -204
rect 1238 -312 1438 -296
rect 1238 -346 1287 -312
rect 1321 -346 1355 -312
rect 1389 -346 1438 -312
rect 1238 -384 1438 -346
rect 1689 -312 1889 -296
rect 1689 -346 1738 -312
rect 1772 -346 1806 -312
rect 1840 -346 1889 -312
rect 1689 -384 1889 -346
rect 1947 -312 2147 -296
rect 1947 -346 1996 -312
rect 2030 -346 2064 -312
rect 2098 -346 2147 -312
rect 1947 -384 2147 -346
rect 2205 -312 2405 -296
rect 2205 -346 2254 -312
rect 2288 -346 2322 -312
rect 2356 -346 2405 -312
rect 2205 -384 2405 -346
rect 2463 -312 2663 -296
rect 2463 -346 2512 -312
rect 2546 -346 2580 -312
rect 2614 -346 2663 -312
rect 2463 -384 2663 -346
rect 2915 -312 3115 -296
rect 2915 -346 2964 -312
rect 2998 -346 3032 -312
rect 3066 -346 3115 -312
rect 2915 -384 3115 -346
rect 1238 -610 1438 -584
rect 1689 -610 1889 -584
rect 1947 -610 2147 -584
rect 2205 -610 2405 -584
rect 2463 -610 2663 -584
rect 2915 -610 3115 -584
<< polycont >>
rect 1287 403 1321 437
rect 1355 403 1389 437
rect 1738 403 1772 437
rect 1806 403 1840 437
rect 1996 403 2030 437
rect 2064 403 2098 437
rect 2254 403 2288 437
rect 2322 403 2356 437
rect 2512 403 2546 437
rect 2580 403 2614 437
rect 2964 403 2998 437
rect 3032 403 3066 437
rect 1287 -204 1321 -170
rect 1355 -204 1389 -170
rect 1738 -204 1772 -170
rect 1806 -204 1840 -170
rect 1996 -204 2030 -170
rect 2064 -204 2098 -170
rect 2254 -204 2288 -170
rect 2322 -204 2356 -170
rect 2512 -204 2546 -170
rect 2580 -204 2614 -170
rect 2964 -204 2998 -170
rect 3032 -204 3066 -170
rect 1287 -346 1321 -312
rect 1355 -346 1389 -312
rect 1738 -346 1772 -312
rect 1806 -346 1840 -312
rect 1996 -346 2030 -312
rect 2064 -346 2098 -312
rect 2254 -346 2288 -312
rect 2322 -346 2356 -312
rect 2512 -346 2546 -312
rect 2580 -346 2614 -312
rect 2964 -346 2998 -312
rect 3032 -346 3066 -312
<< locali >>
rect 1074 502 1238 536
rect 1293 502 1310 536
rect 1361 502 1382 536
rect 1429 502 1454 536
rect 1497 502 1526 536
rect 1565 502 1598 536
rect 1633 502 1667 536
rect 1704 502 1735 536
rect 1776 502 1803 536
rect 1848 502 1871 536
rect 1920 502 1939 536
rect 1992 502 2007 536
rect 2064 502 2075 536
rect 2136 502 2143 536
rect 2208 502 2211 536
rect 2245 502 2246 536
rect 2313 502 2318 536
rect 2381 502 2390 536
rect 2449 502 2462 536
rect 2517 502 2534 536
rect 2585 502 2606 536
rect 2653 502 2678 536
rect 2721 502 2750 536
rect 2789 502 2822 536
rect 2857 502 2891 536
rect 2928 502 2959 536
rect 3000 502 3027 536
rect 3072 502 3095 536
rect 3144 502 3279 536
rect 1074 371 1108 502
rect 1238 403 1285 437
rect 1321 403 1355 437
rect 1391 403 1438 437
rect 1689 403 1736 437
rect 1772 403 1806 437
rect 1842 403 1889 437
rect 1947 403 1994 437
rect 2030 403 2064 437
rect 2100 403 2147 437
rect 2205 403 2252 437
rect 2288 403 2322 437
rect 2358 403 2405 437
rect 2463 403 2510 437
rect 2546 403 2580 437
rect 2616 403 2663 437
rect 2915 403 2962 437
rect 2998 403 3032 437
rect 3068 403 3115 437
rect 3245 371 3279 502
rect 1074 299 1108 317
rect 1074 227 1108 249
rect 1074 155 1108 181
rect 1192 350 1226 369
rect 1192 282 1226 284
rect 1192 246 1226 248
rect 1192 161 1226 180
rect 1450 350 1484 369
rect 1450 282 1484 284
rect 1450 246 1484 248
rect 1450 161 1484 180
rect 1643 350 1677 369
rect 1643 282 1677 284
rect 1643 246 1677 248
rect 1643 161 1677 180
rect 1901 350 1935 369
rect 1901 282 1935 284
rect 1901 246 1935 248
rect 1901 161 1935 180
rect 2159 350 2193 369
rect 2159 282 2193 284
rect 2159 246 2193 248
rect 2159 161 2193 180
rect 2417 350 2451 369
rect 2417 282 2451 284
rect 2417 246 2451 248
rect 2417 161 2451 180
rect 2675 350 2709 369
rect 2675 282 2709 284
rect 2675 246 2709 248
rect 2675 161 2709 180
rect 2869 350 2903 369
rect 2869 282 2903 284
rect 2869 246 2903 248
rect 2869 161 2903 180
rect 3127 350 3161 369
rect 3127 282 3161 284
rect 3127 246 3161 248
rect 3127 161 3161 180
rect 3245 299 3279 317
rect 3245 227 3279 249
rect 1074 59 1108 113
rect 3245 155 3279 181
rect 1074 -13 1108 20
rect 1074 -82 1108 -48
rect 1074 -150 1108 -119
rect 1192 53 1226 72
rect 1192 -15 1226 -13
rect 1192 -51 1226 -49
rect 1192 -136 1226 -117
rect 1450 53 1484 72
rect 1450 -15 1484 -13
rect 1450 -51 1484 -49
rect 1450 -136 1484 -117
rect 1643 53 1677 72
rect 1643 -15 1677 -13
rect 1643 -51 1677 -49
rect 1643 -136 1677 -117
rect 1901 53 1935 72
rect 1901 -15 1935 -13
rect 1901 -51 1935 -49
rect 1901 -136 1935 -117
rect 2159 53 2193 72
rect 2159 -15 2193 -13
rect 2159 -51 2193 -49
rect 2159 -136 2193 -117
rect 2417 53 2451 72
rect 2417 -15 2451 -13
rect 2417 -51 2451 -49
rect 2417 -136 2451 -117
rect 2675 53 2709 72
rect 2675 -15 2709 -13
rect 2675 -51 2709 -49
rect 2675 -136 2709 -117
rect 2869 53 2903 72
rect 2869 -15 2903 -13
rect 2869 -51 2903 -49
rect 2869 -136 2903 -117
rect 3127 53 3161 72
rect 3127 -15 3161 -13
rect 3127 -51 3161 -49
rect 3127 -136 3161 -117
rect 3245 59 3279 113
rect 3245 -13 3279 20
rect 3245 -82 3279 -48
rect 3245 -150 3279 -119
rect 1074 -218 1108 -191
rect 1238 -204 1285 -170
rect 1321 -204 1355 -170
rect 1391 -204 1438 -170
rect 1689 -204 1736 -170
rect 1772 -204 1806 -170
rect 1842 -204 1889 -170
rect 1947 -204 1994 -170
rect 2030 -204 2064 -170
rect 2100 -204 2147 -170
rect 2205 -204 2252 -170
rect 2288 -204 2322 -170
rect 2358 -204 2405 -170
rect 2463 -204 2510 -170
rect 2546 -204 2580 -170
rect 2616 -204 2663 -170
rect 2915 -204 2962 -170
rect 2998 -204 3032 -170
rect 3068 -204 3115 -170
rect 1074 -286 1108 -263
rect 3245 -218 3279 -191
rect 3245 -286 3279 -263
rect 1074 -354 1108 -335
rect 1238 -346 1285 -312
rect 1321 -346 1355 -312
rect 1391 -346 1438 -312
rect 1689 -346 1736 -312
rect 1772 -346 1806 -312
rect 1842 -346 1889 -312
rect 1947 -346 1994 -312
rect 2030 -346 2064 -312
rect 2100 -346 2147 -312
rect 2205 -346 2252 -312
rect 2288 -346 2322 -312
rect 2358 -346 2405 -312
rect 2463 -346 2510 -312
rect 2546 -346 2580 -312
rect 2616 -346 2663 -312
rect 2915 -346 2962 -312
rect 2998 -346 3032 -312
rect 3068 -346 3115 -312
rect 3245 -354 3279 -335
rect 1074 -422 1108 -407
rect 1074 -490 1108 -479
rect 1074 -558 1108 -551
rect 1192 -399 1226 -380
rect 1192 -467 1226 -465
rect 1192 -503 1226 -501
rect 1192 -588 1226 -569
rect 1450 -399 1484 -380
rect 1450 -467 1484 -465
rect 1450 -503 1484 -501
rect 1450 -588 1484 -569
rect 1643 -399 1677 -380
rect 1643 -467 1677 -465
rect 1643 -503 1677 -501
rect 1643 -588 1677 -569
rect 1901 -399 1935 -380
rect 1901 -467 1935 -465
rect 1901 -503 1935 -501
rect 1901 -588 1935 -569
rect 2159 -399 2193 -380
rect 2159 -467 2193 -465
rect 2159 -503 2193 -501
rect 2159 -588 2193 -569
rect 2417 -399 2451 -380
rect 2417 -467 2451 -465
rect 2417 -503 2451 -501
rect 2417 -588 2451 -569
rect 2675 -399 2709 -380
rect 2675 -467 2709 -465
rect 2675 -503 2709 -501
rect 2675 -588 2709 -569
rect 2869 -399 2903 -380
rect 2869 -467 2903 -465
rect 2869 -503 2903 -501
rect 2869 -588 2903 -569
rect 3127 -399 3161 -380
rect 3127 -467 3161 -465
rect 3127 -503 3161 -501
rect 3127 -588 3161 -569
rect 3245 -422 3279 -407
rect 3245 -490 3279 -479
rect 3245 -558 3279 -551
rect 1074 -694 1108 -592
rect 3245 -694 3279 -592
rect 1074 -728 1238 -694
rect 1293 -728 1310 -694
rect 1361 -728 1382 -694
rect 1429 -728 1454 -694
rect 1497 -728 1526 -694
rect 1565 -728 1598 -694
rect 1633 -728 1667 -694
rect 1704 -728 1735 -694
rect 1776 -728 1803 -694
rect 1848 -728 1871 -694
rect 1920 -728 1939 -694
rect 1992 -728 2007 -694
rect 2064 -728 2075 -694
rect 2136 -728 2143 -694
rect 2208 -728 2211 -694
rect 2245 -728 2246 -694
rect 2313 -728 2318 -694
rect 2381 -728 2390 -694
rect 2449 -728 2462 -694
rect 2517 -728 2534 -694
rect 2585 -728 2606 -694
rect 2653 -728 2678 -694
rect 2721 -728 2750 -694
rect 2789 -728 2822 -694
rect 2857 -728 2891 -694
rect 2928 -728 2959 -694
rect 3000 -728 3027 -694
rect 3072 -728 3095 -694
rect 3129 -728 3279 -694
<< viali >>
rect 1238 502 1259 536
rect 1259 502 1272 536
rect 1310 502 1327 536
rect 1327 502 1344 536
rect 1382 502 1395 536
rect 1395 502 1416 536
rect 1454 502 1463 536
rect 1463 502 1488 536
rect 1526 502 1531 536
rect 1531 502 1560 536
rect 1598 502 1599 536
rect 1599 502 1632 536
rect 1670 502 1701 536
rect 1701 502 1704 536
rect 1742 502 1769 536
rect 1769 502 1776 536
rect 1814 502 1837 536
rect 1837 502 1848 536
rect 1886 502 1905 536
rect 1905 502 1920 536
rect 1958 502 1973 536
rect 1973 502 1992 536
rect 2030 502 2041 536
rect 2041 502 2064 536
rect 2102 502 2109 536
rect 2109 502 2136 536
rect 2174 502 2177 536
rect 2177 502 2208 536
rect 2246 502 2279 536
rect 2279 502 2280 536
rect 2318 502 2347 536
rect 2347 502 2352 536
rect 2390 502 2415 536
rect 2415 502 2424 536
rect 2462 502 2483 536
rect 2483 502 2496 536
rect 2534 502 2551 536
rect 2551 502 2568 536
rect 2606 502 2619 536
rect 2619 502 2640 536
rect 2678 502 2687 536
rect 2687 502 2712 536
rect 2750 502 2755 536
rect 2755 502 2784 536
rect 2822 502 2823 536
rect 2823 502 2856 536
rect 2894 502 2925 536
rect 2925 502 2928 536
rect 2966 502 2993 536
rect 2993 502 3000 536
rect 3038 502 3061 536
rect 3061 502 3072 536
rect 3110 502 3129 536
rect 3129 502 3144 536
rect 1285 403 1287 437
rect 1287 403 1319 437
rect 1357 403 1389 437
rect 1389 403 1391 437
rect 1736 403 1738 437
rect 1738 403 1770 437
rect 1808 403 1840 437
rect 1840 403 1842 437
rect 1994 403 1996 437
rect 1996 403 2028 437
rect 2066 403 2098 437
rect 2098 403 2100 437
rect 2252 403 2254 437
rect 2254 403 2286 437
rect 2324 403 2356 437
rect 2356 403 2358 437
rect 2510 403 2512 437
rect 2512 403 2544 437
rect 2582 403 2614 437
rect 2614 403 2616 437
rect 2962 403 2964 437
rect 2964 403 2996 437
rect 3034 403 3066 437
rect 3066 403 3068 437
rect 1074 351 1108 371
rect 1074 337 1108 351
rect 1074 283 1108 299
rect 1074 265 1108 283
rect 1074 215 1108 227
rect 1074 193 1108 215
rect 1192 316 1226 318
rect 1192 284 1226 316
rect 1192 214 1226 246
rect 1192 212 1226 214
rect 1450 316 1484 318
rect 1450 284 1484 316
rect 1450 214 1484 246
rect 1450 212 1484 214
rect 1643 316 1677 318
rect 1643 284 1677 316
rect 1643 214 1677 246
rect 1643 212 1677 214
rect 1901 316 1935 318
rect 1901 284 1935 316
rect 1901 214 1935 246
rect 1901 212 1935 214
rect 2159 316 2193 318
rect 2159 284 2193 316
rect 2159 214 2193 246
rect 2159 212 2193 214
rect 2417 316 2451 318
rect 2417 284 2451 316
rect 2417 214 2451 246
rect 2417 212 2451 214
rect 2675 316 2709 318
rect 2675 284 2709 316
rect 2675 214 2709 246
rect 2675 212 2709 214
rect 2869 316 2903 318
rect 2869 284 2903 316
rect 2869 214 2903 246
rect 2869 212 2903 214
rect 3127 316 3161 318
rect 3127 284 3161 316
rect 3127 214 3161 246
rect 3127 212 3161 214
rect 3245 351 3279 371
rect 3245 337 3279 351
rect 3245 283 3279 299
rect 3245 265 3279 283
rect 3245 215 3279 227
rect 3245 193 3279 215
rect 1074 147 1108 155
rect 1074 121 1108 147
rect 3245 147 3279 155
rect 3245 121 3279 147
rect 1074 54 1108 59
rect 1074 25 1108 54
rect 1074 -14 1108 -13
rect 1074 -47 1108 -14
rect 1074 -116 1108 -85
rect 1074 -119 1108 -116
rect 1192 19 1226 21
rect 1192 -13 1226 19
rect 1192 -83 1226 -51
rect 1192 -85 1226 -83
rect 1450 19 1484 21
rect 1450 -13 1484 19
rect 1450 -83 1484 -51
rect 1450 -85 1484 -83
rect 1643 19 1677 21
rect 1643 -13 1677 19
rect 1643 -83 1677 -51
rect 1643 -85 1677 -83
rect 1901 19 1935 21
rect 1901 -13 1935 19
rect 1901 -83 1935 -51
rect 1901 -85 1935 -83
rect 2159 19 2193 21
rect 2159 -13 2193 19
rect 2159 -83 2193 -51
rect 2159 -85 2193 -83
rect 2417 19 2451 21
rect 2417 -13 2451 19
rect 2417 -83 2451 -51
rect 2417 -85 2451 -83
rect 2675 19 2709 21
rect 2675 -13 2709 19
rect 2675 -83 2709 -51
rect 2675 -85 2709 -83
rect 2869 19 2903 21
rect 2869 -13 2903 19
rect 2869 -83 2903 -51
rect 2869 -85 2903 -83
rect 3127 19 3161 21
rect 3127 -13 3161 19
rect 3127 -83 3161 -51
rect 3127 -85 3161 -83
rect 3245 54 3279 59
rect 3245 25 3279 54
rect 3245 -14 3279 -13
rect 3245 -47 3279 -14
rect 3245 -116 3279 -85
rect 3245 -119 3279 -116
rect 1074 -184 1108 -157
rect 1074 -191 1108 -184
rect 1285 -204 1287 -170
rect 1287 -204 1319 -170
rect 1357 -204 1389 -170
rect 1389 -204 1391 -170
rect 1736 -204 1738 -170
rect 1738 -204 1770 -170
rect 1808 -204 1840 -170
rect 1840 -204 1842 -170
rect 1994 -204 1996 -170
rect 1996 -204 2028 -170
rect 2066 -204 2098 -170
rect 2098 -204 2100 -170
rect 2252 -204 2254 -170
rect 2254 -204 2286 -170
rect 2324 -204 2356 -170
rect 2356 -204 2358 -170
rect 2510 -204 2512 -170
rect 2512 -204 2544 -170
rect 2582 -204 2614 -170
rect 2614 -204 2616 -170
rect 2962 -204 2964 -170
rect 2964 -204 2996 -170
rect 3034 -204 3066 -170
rect 3066 -204 3068 -170
rect 3245 -184 3279 -157
rect 3245 -191 3279 -184
rect 1074 -252 1108 -229
rect 1074 -263 1108 -252
rect 1074 -320 1108 -301
rect 3245 -252 3279 -229
rect 3245 -263 3279 -252
rect 1074 -335 1108 -320
rect 1285 -346 1287 -312
rect 1287 -346 1319 -312
rect 1357 -346 1389 -312
rect 1389 -346 1391 -312
rect 1736 -346 1738 -312
rect 1738 -346 1770 -312
rect 1808 -346 1840 -312
rect 1840 -346 1842 -312
rect 1994 -346 1996 -312
rect 1996 -346 2028 -312
rect 2066 -346 2098 -312
rect 2098 -346 2100 -312
rect 2252 -346 2254 -312
rect 2254 -346 2286 -312
rect 2324 -346 2356 -312
rect 2356 -346 2358 -312
rect 2510 -346 2512 -312
rect 2512 -346 2544 -312
rect 2582 -346 2614 -312
rect 2614 -346 2616 -312
rect 2962 -346 2964 -312
rect 2964 -346 2996 -312
rect 3034 -346 3066 -312
rect 3066 -346 3068 -312
rect 3245 -320 3279 -301
rect 3245 -335 3279 -320
rect 1074 -388 1108 -373
rect 1074 -407 1108 -388
rect 1074 -456 1108 -445
rect 1074 -479 1108 -456
rect 1074 -524 1108 -517
rect 1074 -551 1108 -524
rect 1192 -433 1226 -431
rect 1192 -465 1226 -433
rect 1192 -535 1226 -503
rect 1192 -537 1226 -535
rect 1450 -433 1484 -431
rect 1450 -465 1484 -433
rect 1450 -535 1484 -503
rect 1450 -537 1484 -535
rect 1643 -433 1677 -431
rect 1643 -465 1677 -433
rect 1643 -535 1677 -503
rect 1643 -537 1677 -535
rect 1901 -433 1935 -431
rect 1901 -465 1935 -433
rect 1901 -535 1935 -503
rect 1901 -537 1935 -535
rect 2159 -433 2193 -431
rect 2159 -465 2193 -433
rect 2159 -535 2193 -503
rect 2159 -537 2193 -535
rect 2417 -433 2451 -431
rect 2417 -465 2451 -433
rect 2417 -535 2451 -503
rect 2417 -537 2451 -535
rect 2675 -433 2709 -431
rect 2675 -465 2709 -433
rect 2675 -535 2709 -503
rect 2675 -537 2709 -535
rect 2869 -433 2903 -431
rect 2869 -465 2903 -433
rect 2869 -535 2903 -503
rect 2869 -537 2903 -535
rect 3127 -433 3161 -431
rect 3127 -465 3161 -433
rect 3127 -535 3161 -503
rect 3127 -537 3161 -535
rect 3245 -388 3279 -373
rect 3245 -407 3279 -388
rect 3245 -456 3279 -445
rect 3245 -479 3279 -456
rect 3245 -524 3279 -517
rect 3245 -551 3279 -524
rect 1238 -728 1259 -694
rect 1259 -728 1272 -694
rect 1310 -728 1327 -694
rect 1327 -728 1344 -694
rect 1382 -728 1395 -694
rect 1395 -728 1416 -694
rect 1454 -728 1463 -694
rect 1463 -728 1488 -694
rect 1526 -728 1531 -694
rect 1531 -728 1560 -694
rect 1598 -728 1599 -694
rect 1599 -728 1632 -694
rect 1670 -728 1701 -694
rect 1701 -728 1704 -694
rect 1742 -728 1769 -694
rect 1769 -728 1776 -694
rect 1814 -728 1837 -694
rect 1837 -728 1848 -694
rect 1886 -728 1905 -694
rect 1905 -728 1920 -694
rect 1958 -728 1973 -694
rect 1973 -728 1992 -694
rect 2030 -728 2041 -694
rect 2041 -728 2064 -694
rect 2102 -728 2109 -694
rect 2109 -728 2136 -694
rect 2174 -728 2177 -694
rect 2177 -728 2208 -694
rect 2246 -728 2279 -694
rect 2279 -728 2280 -694
rect 2318 -728 2347 -694
rect 2347 -728 2352 -694
rect 2390 -728 2415 -694
rect 2415 -728 2424 -694
rect 2462 -728 2483 -694
rect 2483 -728 2496 -694
rect 2534 -728 2551 -694
rect 2551 -728 2568 -694
rect 2606 -728 2619 -694
rect 2619 -728 2640 -694
rect 2678 -728 2687 -694
rect 2687 -728 2712 -694
rect 2750 -728 2755 -694
rect 2755 -728 2784 -694
rect 2822 -728 2823 -694
rect 2823 -728 2856 -694
rect 2894 -728 2925 -694
rect 2925 -728 2928 -694
rect 2966 -728 2993 -694
rect 2993 -728 3000 -694
rect 3038 -728 3061 -694
rect 3061 -728 3072 -694
<< metal1 >>
rect 1049 536 3304 561
rect 1049 502 1238 536
rect 1272 502 1310 536
rect 1344 502 1382 536
rect 1416 502 1454 536
rect 1488 502 1526 536
rect 1560 502 1598 536
rect 1632 502 1670 536
rect 1704 502 1742 536
rect 1776 502 1814 536
rect 1848 502 1886 536
rect 1920 502 1958 536
rect 1992 502 2030 536
rect 2064 502 2102 536
rect 2136 502 2174 536
rect 2208 502 2246 536
rect 2280 502 2318 536
rect 2352 502 2390 536
rect 2424 502 2462 536
rect 2496 502 2534 536
rect 2568 502 2606 536
rect 2640 502 2678 536
rect 2712 502 2750 536
rect 2784 502 2822 536
rect 2856 502 2894 536
rect 2928 502 2966 536
rect 3000 502 3038 536
rect 3072 502 3110 536
rect 3144 502 3304 536
rect 1049 437 3304 502
rect 1049 403 1285 437
rect 1319 403 1357 437
rect 1391 403 1736 437
rect 1770 403 1808 437
rect 1842 403 1994 437
rect 2028 403 2066 437
rect 2100 403 2252 437
rect 2286 403 2324 437
rect 2358 403 2510 437
rect 2544 403 2582 437
rect 2616 403 2962 437
rect 2996 403 3034 437
rect 3068 403 3304 437
rect 1049 371 3304 403
rect 1049 337 1074 371
rect 1108 337 3245 371
rect 3279 337 3304 371
rect 1049 318 3304 337
rect 1049 299 1192 318
rect 1049 265 1074 299
rect 1108 284 1192 299
rect 1226 284 1450 318
rect 1484 284 1643 318
rect 1677 284 1901 318
rect 1935 284 2159 318
rect 2193 284 2417 318
rect 2451 284 2675 318
rect 2709 284 2869 318
rect 2903 284 3127 318
rect 3161 299 3304 318
rect 3161 284 3245 299
rect 1108 265 3245 284
rect 3279 265 3304 299
rect 1049 246 3304 265
rect 1049 227 1192 246
rect 1049 193 1074 227
rect 1108 212 1192 227
rect 1226 212 1450 246
rect 1484 212 1643 246
rect 1677 212 1901 246
rect 1935 212 2159 246
rect 2193 212 2417 246
rect 2451 212 2675 246
rect 2709 212 2869 246
rect 2903 212 3127 246
rect 3161 227 3304 246
rect 3161 212 3245 227
rect 1108 193 3245 212
rect 3279 193 3304 227
rect 1049 165 3304 193
rect 1049 155 1563 165
rect 1049 121 1074 155
rect 1108 121 1563 155
rect 1049 68 1563 121
rect 2863 155 3304 165
rect 2863 121 3245 155
rect 3279 121 3304 155
rect 1049 59 1683 68
rect 1049 25 1074 59
rect 1108 25 1683 59
rect 1049 21 1683 25
rect 1049 -13 1192 21
rect 1226 -13 1450 21
rect 1484 -13 1643 21
rect 1677 -13 1683 21
rect 1049 -47 1074 -13
rect 1108 -47 1683 -13
rect 1049 -51 1683 -47
rect 1049 -85 1192 -51
rect 1226 -85 1450 -51
rect 1484 -85 1643 -51
rect 1677 -85 1683 -51
rect 1049 -119 1074 -85
rect 1108 -119 1683 -85
rect 1049 -132 1683 -119
rect 1895 21 1941 68
rect 1895 -13 1901 21
rect 1935 -13 1941 21
rect 1895 -51 1941 -13
rect 1895 -85 1901 -51
rect 1935 -85 1941 -51
rect 1895 -132 1941 -85
rect 2153 21 2199 68
rect 2153 -13 2159 21
rect 2193 -13 2199 21
rect 2153 -51 2199 -13
rect 2153 -85 2159 -51
rect 2193 -85 2199 -51
rect 2153 -132 2199 -85
rect 2411 21 2457 68
rect 2411 -13 2417 21
rect 2451 -13 2457 21
rect 2411 -51 2457 -13
rect 2411 -85 2417 -51
rect 2451 -85 2457 -51
rect 2411 -132 2457 -85
rect 2669 21 2790 68
rect 2669 -13 2675 21
rect 2709 -13 2790 21
rect 2669 -51 2790 -13
rect 2669 -85 2675 -51
rect 2709 -85 2790 -51
rect 1049 -157 1563 -132
rect 1049 -191 1074 -157
rect 1108 -170 1563 -157
rect 2669 -164 2790 -85
rect 1108 -191 1285 -170
rect 1049 -204 1285 -191
rect 1319 -204 1357 -170
rect 1391 -204 1563 -170
rect 1049 -229 1563 -204
rect 1049 -263 1074 -229
rect 1108 -263 1563 -229
rect 1693 -170 2790 -164
rect 1693 -172 1736 -170
rect 1770 -172 1808 -170
rect 1842 -172 1994 -170
rect 2028 -172 2066 -170
rect 2100 -172 2252 -170
rect 2286 -172 2324 -170
rect 2358 -172 2510 -170
rect 1693 -224 1722 -172
rect 1774 -224 1786 -172
rect 1842 -204 1850 -172
rect 1838 -224 1850 -204
rect 1902 -224 1956 -172
rect 2008 -224 2020 -204
rect 2072 -224 2084 -204
rect 2136 -224 2196 -172
rect 2248 -204 2252 -172
rect 2248 -224 2260 -204
rect 2312 -224 2324 -172
rect 2376 -204 2510 -172
rect 2544 -204 2582 -170
rect 2616 -204 2790 -170
rect 2376 -210 2790 -204
rect 2863 59 3304 121
rect 2863 25 3245 59
rect 3279 25 3304 59
rect 2863 21 3304 25
rect 2863 -13 2869 21
rect 2903 -13 3127 21
rect 3161 -13 3304 21
rect 2863 -47 3245 -13
rect 3279 -47 3304 -13
rect 2863 -51 3304 -47
rect 2863 -85 2869 -51
rect 2903 -85 3127 -51
rect 3161 -85 3304 -51
rect 2863 -119 3245 -85
rect 3279 -119 3304 -85
rect 2863 -157 3304 -119
rect 2863 -170 3245 -157
rect 2863 -204 2962 -170
rect 2996 -204 3034 -170
rect 3068 -191 3245 -170
rect 3279 -191 3304 -157
rect 3068 -204 3304 -191
rect 2376 -224 2532 -210
rect 1693 -234 2532 -224
rect 2863 -229 3304 -204
rect 1049 -301 1563 -263
rect 1049 -335 1074 -301
rect 1108 -306 1563 -301
rect 2863 -263 3245 -229
rect 3279 -263 3304 -229
rect 2863 -301 3304 -263
rect 2863 -306 3245 -301
rect 1108 -312 3245 -306
rect 1108 -335 1285 -312
rect 1049 -346 1285 -335
rect 1319 -346 1357 -312
rect 1391 -346 1736 -312
rect 1770 -346 1808 -312
rect 1842 -346 1994 -312
rect 2028 -346 2066 -312
rect 2100 -346 2252 -312
rect 2286 -346 2324 -312
rect 2358 -346 2510 -312
rect 2544 -346 2582 -312
rect 2616 -346 2962 -312
rect 2996 -346 3034 -312
rect 3068 -335 3245 -312
rect 3279 -335 3304 -301
rect 3068 -346 3304 -335
rect 1049 -373 3304 -346
rect 1049 -407 1074 -373
rect 1108 -407 3245 -373
rect 3279 -407 3304 -373
rect 1049 -431 3304 -407
rect 1049 -445 1192 -431
rect 1049 -479 1074 -445
rect 1108 -465 1192 -445
rect 1226 -465 1450 -431
rect 1484 -465 1643 -431
rect 1677 -465 1901 -431
rect 1935 -465 2159 -431
rect 2193 -465 2417 -431
rect 2451 -465 2675 -431
rect 2709 -465 2869 -431
rect 2903 -465 3127 -431
rect 3161 -445 3304 -431
rect 3161 -465 3245 -445
rect 1108 -479 3245 -465
rect 3279 -479 3304 -445
rect 1049 -503 3304 -479
rect 1049 -517 1192 -503
rect 1049 -551 1074 -517
rect 1108 -537 1192 -517
rect 1226 -537 1450 -503
rect 1484 -537 1643 -503
rect 1677 -537 1901 -503
rect 1935 -537 2159 -503
rect 2193 -537 2417 -503
rect 2451 -537 2675 -503
rect 2709 -537 2869 -503
rect 2903 -537 3127 -503
rect 3161 -517 3304 -503
rect 3161 -537 3245 -517
rect 1108 -551 3245 -537
rect 3279 -551 3304 -517
rect 1049 -694 3304 -551
rect 1049 -728 1238 -694
rect 1272 -728 1310 -694
rect 1344 -728 1382 -694
rect 1416 -728 1454 -694
rect 1488 -728 1526 -694
rect 1560 -728 1598 -694
rect 1632 -728 1670 -694
rect 1704 -728 1742 -694
rect 1776 -728 1814 -694
rect 1848 -728 1886 -694
rect 1920 -728 1958 -694
rect 1992 -728 2030 -694
rect 2064 -728 2102 -694
rect 2136 -728 2174 -694
rect 2208 -728 2246 -694
rect 2280 -728 2318 -694
rect 2352 -728 2390 -694
rect 2424 -728 2462 -694
rect 2496 -728 2534 -694
rect 2568 -728 2606 -694
rect 2640 -728 2678 -694
rect 2712 -728 2750 -694
rect 2784 -728 2822 -694
rect 2856 -728 2894 -694
rect 2928 -728 2966 -694
rect 3000 -728 3038 -694
rect 3072 -728 3304 -694
rect 1049 -753 3304 -728
<< via1 >>
rect 1722 -204 1736 -172
rect 1736 -204 1770 -172
rect 1770 -204 1774 -172
rect 1722 -224 1774 -204
rect 1786 -204 1808 -172
rect 1808 -204 1838 -172
rect 1786 -224 1838 -204
rect 1850 -224 1902 -172
rect 1956 -204 1994 -172
rect 1994 -204 2008 -172
rect 2020 -204 2028 -172
rect 2028 -204 2066 -172
rect 2066 -204 2072 -172
rect 2084 -204 2100 -172
rect 2100 -204 2136 -172
rect 1956 -224 2008 -204
rect 2020 -224 2072 -204
rect 2084 -224 2136 -204
rect 2196 -224 2248 -172
rect 2260 -204 2286 -172
rect 2286 -204 2312 -172
rect 2260 -224 2312 -204
rect 2324 -204 2358 -172
rect 2358 -204 2376 -172
rect 2324 -224 2376 -204
<< metal2 >>
rect 1713 -172 2702 -164
rect 1713 -224 1722 -172
rect 1774 -224 1786 -172
rect 1838 -224 1850 -172
rect 1902 -224 1956 -172
rect 2008 -224 2020 -172
rect 2072 -224 2084 -172
rect 2136 -224 2196 -172
rect 2248 -224 2260 -172
rect 2312 -224 2324 -172
rect 2376 -224 2702 -172
rect 1713 -265 2702 -224
<< labels >>
flabel metal1 s 1120 -651 1537 466 2 FreeSans 3126 0 0 0 AVSS
port 1 nsew
flabel metal2 s 1724 -250 2688 -180 2 FreeSans 3126 0 0 0 VB3
port 2 nsew
<< end >>
