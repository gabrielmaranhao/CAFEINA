magic
tech sky130A
magscale 1 2
timestamp 1698351692
<< nwell >>
rect 70 7344 6652 7795
rect 7401 6799 10893 7301
<< pwell >>
rect 7412 7361 10882 7481
<< mvpsubdiff >>
rect 7438 7387 10856 7455
<< mvnsubdiff >>
rect 7467 7201 10827 7235
<< locali >>
rect 41 8249 183 8288
rect 41 8215 60 8249
rect 94 8215 132 8249
rect 166 8215 183 8249
rect 41 7451 183 8215
rect 6891 8245 7134 8286
rect 6891 8139 6937 8245
rect 7115 8139 7134 8245
rect 6891 7455 7134 8139
rect 9224 8046 9270 8060
rect 9224 8012 9230 8046
rect 9264 8012 9270 8046
rect 9224 7974 9270 8012
rect 9224 7940 9230 7974
rect 9264 7940 9270 7974
rect 9224 7902 9270 7940
rect 9224 7868 9230 7902
rect 9264 7868 9270 7902
rect 9224 7854 9270 7868
rect 10785 7870 10819 7879
rect 7604 7794 7807 7801
rect 7604 7760 7616 7794
rect 7650 7760 7688 7794
rect 7722 7760 7760 7794
rect 7794 7760 7807 7794
rect 7604 7754 7807 7760
rect 9459 7794 9796 7801
rect 9459 7760 9466 7794
rect 9500 7760 9538 7794
rect 9572 7760 9610 7794
rect 9644 7760 9682 7794
rect 9716 7760 9754 7794
rect 9788 7760 9796 7794
rect 9459 7754 9796 7760
rect 10785 7798 10819 7836
rect 10785 7726 10819 7764
rect 10785 7683 10819 7692
rect 3043 7451 7134 7455
rect 41 7425 7134 7451
rect 41 7305 6929 7425
rect 35 6388 121 7179
rect 3043 7031 6929 7305
rect 7107 7322 7134 7425
rect 7107 7201 10829 7322
rect 7107 7031 7134 7201
rect 3043 7005 7134 7031
rect 8439 6870 8506 6878
rect 2907 6670 7134 6838
rect 8439 6836 8455 6870
rect 8489 6836 8506 6870
rect 7870 6821 8128 6834
rect 7870 6787 7874 6821
rect 7908 6787 7946 6821
rect 7980 6787 8018 6821
rect 8052 6787 8090 6821
rect 8124 6787 8128 6821
rect 7870 6775 8128 6787
rect 8439 6798 8506 6836
rect 8439 6764 8455 6798
rect 8489 6764 8506 6798
rect 10270 6868 10316 6896
rect 10270 6834 10276 6868
rect 10310 6834 10316 6868
rect 10270 6796 10316 6834
rect 8439 6726 8506 6764
rect 8439 6692 8455 6726
rect 8489 6692 8506 6726
rect 8650 6760 8853 6767
rect 8650 6726 8662 6760
rect 8696 6726 8734 6760
rect 8768 6726 8806 6760
rect 8840 6726 8853 6760
rect 10270 6762 10276 6796
rect 10310 6762 10316 6796
rect 10270 6735 10316 6762
rect 8650 6720 8853 6726
rect 8439 6684 8506 6692
rect 2907 6388 3247 6670
rect 35 6308 3247 6388
rect 35 6202 78 6308
rect 256 6202 523 6308
rect 2933 6276 3247 6308
rect 6089 6388 7134 6670
rect 6089 6276 10860 6388
rect 2933 6202 10860 6276
rect 35 6143 10860 6202
rect 35 5813 689 6143
rect 1006 5813 1393 6029
rect 1778 5813 2165 6029
rect 2550 6011 2937 6029
rect 2550 5833 2655 6011
rect 2833 5833 2937 6011
rect 2550 5813 2937 5833
rect 3322 5813 3709 6029
rect 4094 5813 4481 6029
rect 4866 5813 5253 6029
rect 5638 5813 6025 6029
rect 6410 5813 6797 6029
rect 7182 5813 7569 6029
rect 7954 5813 8341 6029
rect 8726 5813 9113 6029
rect 9498 5813 9885 6029
rect 10202 6011 10340 6030
rect 10202 5617 10218 6011
rect 10324 5617 10340 6011
rect 10656 5813 10837 6029
rect 10202 5598 10340 5617
rect 51 165 234 381
rect 619 165 1006 381
rect 1391 165 1778 381
rect 2163 165 2550 381
rect 2935 165 3322 381
rect 3707 165 4094 381
rect 4479 165 4866 381
rect 5251 165 5638 381
rect 6023 165 6410 381
rect 6795 165 7182 381
rect 7567 165 7954 381
rect 8339 165 8726 381
rect 9111 165 9498 381
rect 9883 165 10270 381
rect 10655 165 10835 381
<< viali >>
rect 60 8215 94 8249
rect 132 8215 166 8249
rect 6937 8139 7115 8245
rect 9230 8012 9264 8046
rect 9230 7940 9264 7974
rect 9230 7868 9264 7902
rect 10785 7836 10819 7870
rect 7616 7760 7650 7794
rect 7688 7760 7722 7794
rect 7760 7760 7794 7794
rect 9466 7760 9500 7794
rect 9538 7760 9572 7794
rect 9610 7760 9644 7794
rect 9682 7760 9716 7794
rect 9754 7760 9788 7794
rect 10785 7764 10819 7798
rect 10785 7692 10819 7726
rect 6929 7031 7107 7425
rect 8455 6836 8489 6870
rect 7874 6787 7908 6821
rect 7946 6787 7980 6821
rect 8018 6787 8052 6821
rect 8090 6787 8124 6821
rect 8455 6764 8489 6798
rect 10276 6834 10310 6868
rect 8455 6692 8489 6726
rect 8662 6726 8696 6760
rect 8734 6726 8768 6760
rect 8806 6726 8840 6760
rect 10276 6762 10310 6796
rect 78 6202 256 6308
rect 523 6202 2933 6308
rect 3247 6276 6089 6670
rect 2655 5833 2833 6011
rect 10218 5617 10324 6011
<< metal1 >>
rect 40 8261 7133 8286
rect 40 8209 60 8261
rect 112 8209 124 8261
rect 176 8209 188 8261
rect 240 8209 252 8261
rect 304 8209 316 8261
rect 368 8209 380 8261
rect 432 8209 444 8261
rect 496 8209 508 8261
rect 560 8209 572 8261
rect 624 8252 7133 8261
rect 624 8209 1057 8252
rect 40 8200 1057 8209
rect 1109 8200 1121 8252
rect 1173 8200 1185 8252
rect 1237 8200 1249 8252
rect 1301 8200 1313 8252
rect 1365 8200 1377 8252
rect 1429 8200 1441 8252
rect 1493 8200 1505 8252
rect 1557 8200 1569 8252
rect 1621 8200 1633 8252
rect 1685 8200 1697 8252
rect 1749 8200 1761 8252
rect 1813 8200 1825 8252
rect 1877 8200 1889 8252
rect 1941 8200 1953 8252
rect 2005 8200 2017 8252
rect 2069 8200 2081 8252
rect 2133 8200 2145 8252
rect 2197 8200 2209 8252
rect 2261 8200 2273 8252
rect 2325 8200 2337 8252
rect 2389 8200 2401 8252
rect 2453 8200 2465 8252
rect 2517 8200 2529 8252
rect 2581 8200 2593 8252
rect 2645 8200 2657 8252
rect 2709 8200 2721 8252
rect 2773 8200 2785 8252
rect 2837 8200 2849 8252
rect 2901 8200 2913 8252
rect 2965 8200 2977 8252
rect 3029 8200 3041 8252
rect 3093 8200 3105 8252
rect 3157 8200 3169 8252
rect 3221 8200 3233 8252
rect 3285 8200 3297 8252
rect 3349 8200 3361 8252
rect 3413 8200 3425 8252
rect 3477 8200 3489 8252
rect 3541 8200 3553 8252
rect 3605 8200 3617 8252
rect 3669 8200 3681 8252
rect 3733 8200 3745 8252
rect 3797 8200 3809 8252
rect 3861 8200 3873 8252
rect 3925 8200 3937 8252
rect 3989 8200 4001 8252
rect 4053 8200 4065 8252
rect 4117 8200 4129 8252
rect 4181 8200 4193 8252
rect 4245 8200 4257 8252
rect 4309 8200 4321 8252
rect 4373 8200 4385 8252
rect 4437 8200 4449 8252
rect 4501 8200 4513 8252
rect 4565 8200 4577 8252
rect 4629 8200 4641 8252
rect 4693 8200 4705 8252
rect 4757 8200 4769 8252
rect 4821 8200 4833 8252
rect 4885 8200 4897 8252
rect 4949 8200 4961 8252
rect 5013 8200 5025 8252
rect 5077 8200 5089 8252
rect 5141 8200 5153 8252
rect 5205 8200 5217 8252
rect 5269 8200 5281 8252
rect 5333 8200 5345 8252
rect 5397 8200 5409 8252
rect 5461 8200 5473 8252
rect 5525 8200 5537 8252
rect 5589 8200 5601 8252
rect 5653 8200 5665 8252
rect 5717 8200 5729 8252
rect 5781 8200 5793 8252
rect 5845 8200 5857 8252
rect 5909 8200 5921 8252
rect 5973 8200 5985 8252
rect 6037 8200 6049 8252
rect 6101 8200 6113 8252
rect 6165 8200 6177 8252
rect 6229 8200 6241 8252
rect 6293 8200 6305 8252
rect 6357 8200 6369 8252
rect 6421 8200 6433 8252
rect 6485 8200 6497 8252
rect 6549 8200 6561 8252
rect 6613 8200 6625 8252
rect 6677 8200 6689 8252
rect 6741 8200 6753 8252
rect 6805 8200 6817 8252
rect 6869 8200 6881 8252
rect 6933 8245 6945 8252
rect 6997 8245 7009 8252
rect 7061 8245 7133 8252
rect 6933 8200 6937 8245
rect 7115 8209 7133 8245
rect 7284 8228 10841 8278
rect 40 8179 6937 8200
rect 709 8139 818 8144
rect 218 8110 376 8127
rect 218 8038 436 8110
rect 709 8087 734 8139
rect 786 8129 818 8139
rect 6910 8139 6937 8179
rect 7115 8139 7134 8209
rect 786 8087 2498 8129
rect 709 8085 2498 8087
rect 2829 8085 2990 8129
rect 709 8082 818 8085
rect 218 8024 282 8038
rect 218 7641 313 8024
rect 375 7641 436 8038
rect 521 7788 567 8040
rect 627 7892 2821 8028
rect 502 7653 2537 7788
rect 218 7568 436 7641
rect 521 7597 567 7653
rect 709 7601 818 7606
rect 709 7597 734 7601
rect 218 7554 375 7568
rect 218 7501 282 7554
rect 521 7553 734 7597
rect 709 7549 734 7553
rect 786 7597 818 7601
rect 2866 7597 2944 8085
rect 2993 7658 3300 7804
rect 786 7556 2990 7597
rect 786 7553 2922 7556
rect 786 7549 818 7553
rect 709 7544 818 7549
rect 3360 7501 3433 8122
rect 3699 8082 3959 8128
rect 3486 7636 3556 8035
rect 218 7453 3433 7501
rect 218 7248 282 7453
rect 3497 7344 3556 7636
rect 185 7121 282 7248
rect 2382 7274 3556 7344
rect 3699 7642 3781 8082
rect 4283 8081 5747 8125
rect 6083 8081 6237 8125
rect 3988 7805 4025 8041
rect 4109 7872 6071 8033
rect 3966 7645 5802 7805
rect 3699 7600 3773 7642
rect 3699 7554 3958 7600
rect 3988 7597 4025 7645
rect 6126 7597 6188 8081
rect 6249 7884 6537 8029
rect 6249 7690 6262 7884
rect 3699 7501 3773 7554
rect 3988 7553 6239 7597
rect 6612 7501 6674 8112
rect 3699 7453 6674 7501
rect 185 6969 263 7121
rect 2382 7074 2452 7274
rect 3699 7165 3773 7453
rect 2265 7064 2452 7074
rect 2265 7047 2287 7064
rect 185 6573 282 6969
rect 25 6308 301 6326
rect 25 6202 78 6308
rect 256 6202 301 6308
rect 25 6185 301 6202
rect 25 5348 133 6185
rect 345 5944 399 7033
rect 781 7012 2287 7047
rect 2339 7047 2452 7064
rect 2767 7074 3773 7165
rect 2339 7012 2738 7047
rect 781 7003 2738 7012
rect 463 6745 634 6972
rect 2382 6952 2452 7003
rect 721 6815 2452 6952
rect 463 6579 2560 6745
rect 463 6569 634 6579
rect 505 6326 634 6569
rect 2629 6533 2693 7003
rect 2767 6949 2842 7074
rect 6752 7065 6823 8044
rect 6910 7425 7134 8139
rect 7284 8176 7338 8228
rect 7390 8176 7402 8228
rect 7454 8176 7466 8228
rect 7518 8176 7530 8228
rect 7582 8176 7594 8228
rect 7646 8176 7658 8228
rect 7710 8176 7722 8228
rect 7774 8176 7786 8228
rect 7838 8176 7850 8228
rect 7902 8176 7914 8228
rect 7966 8176 7978 8228
rect 8030 8176 8042 8228
rect 8094 8176 8106 8228
rect 8158 8176 8170 8228
rect 8222 8176 8234 8228
rect 8286 8176 8298 8228
rect 8350 8176 8362 8228
rect 8414 8176 8426 8228
rect 8478 8176 8490 8228
rect 8542 8176 8554 8228
rect 8606 8176 8618 8228
rect 8670 8176 8682 8228
rect 8734 8176 8746 8228
rect 8798 8176 8810 8228
rect 8862 8176 8874 8228
rect 8926 8176 8938 8228
rect 8990 8176 9002 8228
rect 9054 8176 9066 8228
rect 9118 8176 9130 8228
rect 9182 8176 9194 8228
rect 9246 8176 9258 8228
rect 9310 8176 9322 8228
rect 9374 8176 9386 8228
rect 9438 8176 9450 8228
rect 9502 8176 9514 8228
rect 9566 8176 9578 8228
rect 9630 8176 9642 8228
rect 9694 8176 9706 8228
rect 9758 8176 9770 8228
rect 9822 8176 9834 8228
rect 9886 8176 9898 8228
rect 9950 8176 9962 8228
rect 10014 8176 10026 8228
rect 10078 8176 10090 8228
rect 10142 8176 10154 8228
rect 10206 8176 10218 8228
rect 10270 8176 10282 8228
rect 10334 8176 10346 8228
rect 10398 8176 10410 8228
rect 10462 8176 10474 8228
rect 10526 8176 10538 8228
rect 10590 8176 10602 8228
rect 10654 8176 10666 8228
rect 10718 8176 10730 8228
rect 10782 8176 10841 8228
rect 7284 8125 10841 8176
rect 9218 8051 9276 8072
rect 10128 8052 10300 8053
rect 10128 8051 10156 8052
rect 9218 8046 10156 8051
rect 9218 8012 9230 8046
rect 9264 8012 10156 8046
rect 9218 8001 10156 8012
rect 9218 7974 9276 8001
rect 10128 8000 10156 8001
rect 10208 8000 10220 8052
rect 10272 8000 10300 8052
rect 10128 7999 10300 8000
rect 9218 7940 9230 7974
rect 9264 7940 9276 7974
rect 9218 7902 9276 7940
rect 9218 7868 9230 7902
rect 9264 7868 9276 7902
rect 9218 7842 9276 7868
rect 10779 7870 10825 7891
rect 10779 7836 10785 7870
rect 10819 7836 10825 7870
rect 7592 7803 9808 7807
rect 7592 7794 8339 7803
rect 7592 7760 7616 7794
rect 7650 7760 7688 7794
rect 7722 7760 7760 7794
rect 7794 7760 8339 7794
rect 7592 7751 8339 7760
rect 8391 7751 8403 7803
rect 8455 7751 8467 7803
rect 8519 7794 9808 7803
rect 8519 7760 9466 7794
rect 9500 7760 9538 7794
rect 9572 7760 9610 7794
rect 9644 7760 9682 7794
rect 9716 7760 9754 7794
rect 9788 7760 9808 7794
rect 8519 7751 9808 7760
rect 7592 7748 9808 7751
rect 10779 7798 10825 7836
rect 10779 7764 10785 7798
rect 10819 7764 10825 7798
rect 10779 7728 10825 7764
rect 10743 7727 10915 7728
rect 10743 7675 10771 7727
rect 10823 7675 10835 7727
rect 10887 7675 10915 7727
rect 10743 7674 10915 7675
rect 10779 7671 10825 7674
rect 2756 6573 2842 6949
rect 6407 7015 6825 7065
rect 3167 6794 6174 6842
rect 3167 6670 4362 6794
rect 5246 6670 6174 6794
rect 781 6522 2360 6533
rect 781 6489 2286 6522
rect 2265 6470 2286 6489
rect 2338 6470 2360 6522
rect 2585 6489 2739 6533
rect 2265 6460 2360 6470
rect 3167 6326 3247 6670
rect 493 6308 3247 6326
rect 493 6202 523 6308
rect 2933 6276 3247 6308
rect 6089 6531 6174 6670
rect 6407 6643 6463 7015
rect 6771 6840 6825 7015
rect 6910 7031 6929 7425
rect 7107 7324 7134 7425
rect 7279 7522 10836 7570
rect 7279 7470 7318 7522
rect 7370 7470 7382 7522
rect 7434 7470 7446 7522
rect 7498 7470 7510 7522
rect 7562 7470 7574 7522
rect 7626 7470 7638 7522
rect 7690 7470 7702 7522
rect 7754 7470 7766 7522
rect 7818 7470 7830 7522
rect 7882 7470 7894 7522
rect 7946 7470 7958 7522
rect 8010 7470 8022 7522
rect 8074 7470 8086 7522
rect 8138 7470 8150 7522
rect 8202 7470 8214 7522
rect 8266 7470 8278 7522
rect 8330 7470 8647 7522
rect 8699 7470 8711 7522
rect 8763 7470 8775 7522
rect 8827 7470 8839 7522
rect 8891 7470 8903 7522
rect 8955 7470 8967 7522
rect 9019 7470 9031 7522
rect 9083 7470 9095 7522
rect 9147 7470 9159 7522
rect 9211 7470 9223 7522
rect 9275 7470 9287 7522
rect 9339 7470 9351 7522
rect 9403 7470 9415 7522
rect 9467 7470 9479 7522
rect 9531 7470 9543 7522
rect 9595 7470 9607 7522
rect 9659 7470 9671 7522
rect 9723 7470 9735 7522
rect 9787 7470 9799 7522
rect 9851 7470 9863 7522
rect 9915 7470 9927 7522
rect 9979 7470 9991 7522
rect 10043 7470 10055 7522
rect 10107 7470 10119 7522
rect 10171 7470 10183 7522
rect 10235 7470 10247 7522
rect 10299 7470 10311 7522
rect 10363 7470 10375 7522
rect 10427 7470 10439 7522
rect 10491 7470 10503 7522
rect 10555 7470 10567 7522
rect 10619 7470 10836 7522
rect 7279 7417 10836 7470
rect 7107 7269 10832 7324
rect 7107 7153 7175 7269
rect 8315 7153 8626 7269
rect 10726 7153 10832 7269
rect 7107 7094 10832 7153
rect 7107 7031 7134 7094
rect 10516 7093 10832 7094
rect 6910 6994 7134 7031
rect 8433 6878 8512 6890
rect 8429 6871 8516 6878
rect 6771 6821 8140 6840
rect 6771 6787 7874 6821
rect 7908 6787 7946 6821
rect 7980 6787 8018 6821
rect 8052 6787 8090 6821
rect 8124 6787 8140 6821
rect 6771 6769 8140 6787
rect 8429 6819 8446 6871
rect 8498 6819 8516 6871
rect 8429 6807 8516 6819
rect 6771 6643 6825 6769
rect 8429 6755 8446 6807
rect 8498 6773 8516 6807
rect 10264 6868 10322 6908
rect 10264 6834 10276 6868
rect 10310 6834 10322 6868
rect 10264 6825 10682 6834
rect 10264 6796 10531 6825
rect 8498 6760 8865 6773
rect 8498 6755 8662 6760
rect 8429 6743 8662 6755
rect 8429 6691 8446 6743
rect 8498 6726 8662 6743
rect 8696 6726 8734 6760
rect 8768 6726 8806 6760
rect 8840 6726 8865 6760
rect 8498 6714 8865 6726
rect 10264 6762 10276 6796
rect 10310 6773 10531 6796
rect 10583 6773 10595 6825
rect 10647 6773 10682 6825
rect 10310 6765 10682 6773
rect 10310 6762 10322 6765
rect 10264 6723 10322 6762
rect 8498 6691 8516 6714
rect 8429 6684 8516 6691
rect 8433 6672 8512 6684
rect 6407 6600 6825 6643
rect 6089 6319 10827 6531
rect 6089 6276 6174 6319
rect 2933 6237 6174 6276
rect 10221 6249 10716 6270
rect 2933 6202 6175 6237
rect 493 6185 6175 6202
rect 10221 6197 10248 6249
rect 10300 6197 10312 6249
rect 10364 6197 10376 6249
rect 10428 6197 10440 6249
rect 10492 6197 10504 6249
rect 10556 6197 10568 6249
rect 10620 6197 10632 6249
rect 10684 6197 10716 6249
rect 10221 6176 10716 6197
rect 10221 6045 10315 6176
rect 2635 6011 2853 6026
rect 2635 5944 2655 6011
rect 345 5890 2655 5944
rect 2635 5833 2655 5890
rect 2833 5833 2853 6011
rect 2635 5816 2853 5833
rect 10187 6011 10353 6045
rect 10187 5617 10218 6011
rect 10324 5617 10353 6011
rect 10187 5582 10353 5617
rect 10805 5348 10867 6079
rect 25 4748 10867 5348
rect 25 4348 133 4748
rect 10805 4348 10867 4748
rect 25 3748 10867 4348
rect 25 3348 133 3748
rect 10805 3348 10867 3748
rect 25 2748 10867 3348
rect 25 2348 133 2748
rect 10805 2348 10867 2748
rect 25 1748 10867 2348
rect 25 1348 133 1748
rect 10805 1348 10867 1748
rect 25 748 10867 1348
rect 25 99 133 748
rect 10805 99 10867 748
rect 25 11 10867 99
<< via1 >>
rect 60 8249 112 8261
rect 60 8215 94 8249
rect 94 8215 112 8249
rect 60 8209 112 8215
rect 124 8249 176 8261
rect 124 8215 132 8249
rect 132 8215 166 8249
rect 166 8215 176 8249
rect 124 8209 176 8215
rect 188 8209 240 8261
rect 252 8209 304 8261
rect 316 8209 368 8261
rect 380 8209 432 8261
rect 444 8209 496 8261
rect 508 8209 560 8261
rect 572 8209 624 8261
rect 1057 8200 1109 8252
rect 1121 8200 1173 8252
rect 1185 8200 1237 8252
rect 1249 8200 1301 8252
rect 1313 8200 1365 8252
rect 1377 8200 1429 8252
rect 1441 8200 1493 8252
rect 1505 8200 1557 8252
rect 1569 8200 1621 8252
rect 1633 8200 1685 8252
rect 1697 8200 1749 8252
rect 1761 8200 1813 8252
rect 1825 8200 1877 8252
rect 1889 8200 1941 8252
rect 1953 8200 2005 8252
rect 2017 8200 2069 8252
rect 2081 8200 2133 8252
rect 2145 8200 2197 8252
rect 2209 8200 2261 8252
rect 2273 8200 2325 8252
rect 2337 8200 2389 8252
rect 2401 8200 2453 8252
rect 2465 8200 2517 8252
rect 2529 8200 2581 8252
rect 2593 8200 2645 8252
rect 2657 8200 2709 8252
rect 2721 8200 2773 8252
rect 2785 8200 2837 8252
rect 2849 8200 2901 8252
rect 2913 8200 2965 8252
rect 2977 8200 3029 8252
rect 3041 8200 3093 8252
rect 3105 8200 3157 8252
rect 3169 8200 3221 8252
rect 3233 8200 3285 8252
rect 3297 8200 3349 8252
rect 3361 8200 3413 8252
rect 3425 8200 3477 8252
rect 3489 8200 3541 8252
rect 3553 8200 3605 8252
rect 3617 8200 3669 8252
rect 3681 8200 3733 8252
rect 3745 8200 3797 8252
rect 3809 8200 3861 8252
rect 3873 8200 3925 8252
rect 3937 8200 3989 8252
rect 4001 8200 4053 8252
rect 4065 8200 4117 8252
rect 4129 8200 4181 8252
rect 4193 8200 4245 8252
rect 4257 8200 4309 8252
rect 4321 8200 4373 8252
rect 4385 8200 4437 8252
rect 4449 8200 4501 8252
rect 4513 8200 4565 8252
rect 4577 8200 4629 8252
rect 4641 8200 4693 8252
rect 4705 8200 4757 8252
rect 4769 8200 4821 8252
rect 4833 8200 4885 8252
rect 4897 8200 4949 8252
rect 4961 8200 5013 8252
rect 5025 8200 5077 8252
rect 5089 8200 5141 8252
rect 5153 8200 5205 8252
rect 5217 8200 5269 8252
rect 5281 8200 5333 8252
rect 5345 8200 5397 8252
rect 5409 8200 5461 8252
rect 5473 8200 5525 8252
rect 5537 8200 5589 8252
rect 5601 8200 5653 8252
rect 5665 8200 5717 8252
rect 5729 8200 5781 8252
rect 5793 8200 5845 8252
rect 5857 8200 5909 8252
rect 5921 8200 5973 8252
rect 5985 8200 6037 8252
rect 6049 8200 6101 8252
rect 6113 8200 6165 8252
rect 6177 8200 6229 8252
rect 6241 8200 6293 8252
rect 6305 8200 6357 8252
rect 6369 8200 6421 8252
rect 6433 8200 6485 8252
rect 6497 8200 6549 8252
rect 6561 8200 6613 8252
rect 6625 8200 6677 8252
rect 6689 8200 6741 8252
rect 6753 8200 6805 8252
rect 6817 8200 6869 8252
rect 6881 8200 6933 8252
rect 6945 8245 6997 8252
rect 7009 8245 7061 8252
rect 6945 8200 6997 8245
rect 7009 8200 7061 8245
rect 734 8087 786 8139
rect 734 7549 786 7601
rect 2287 7012 2339 7064
rect 7338 8176 7390 8228
rect 7402 8176 7454 8228
rect 7466 8176 7518 8228
rect 7530 8176 7582 8228
rect 7594 8176 7646 8228
rect 7658 8176 7710 8228
rect 7722 8176 7774 8228
rect 7786 8176 7838 8228
rect 7850 8176 7902 8228
rect 7914 8176 7966 8228
rect 7978 8176 8030 8228
rect 8042 8176 8094 8228
rect 8106 8176 8158 8228
rect 8170 8176 8222 8228
rect 8234 8176 8286 8228
rect 8298 8176 8350 8228
rect 8362 8176 8414 8228
rect 8426 8176 8478 8228
rect 8490 8176 8542 8228
rect 8554 8176 8606 8228
rect 8618 8176 8670 8228
rect 8682 8176 8734 8228
rect 8746 8176 8798 8228
rect 8810 8176 8862 8228
rect 8874 8176 8926 8228
rect 8938 8176 8990 8228
rect 9002 8176 9054 8228
rect 9066 8176 9118 8228
rect 9130 8176 9182 8228
rect 9194 8176 9246 8228
rect 9258 8176 9310 8228
rect 9322 8176 9374 8228
rect 9386 8176 9438 8228
rect 9450 8176 9502 8228
rect 9514 8176 9566 8228
rect 9578 8176 9630 8228
rect 9642 8176 9694 8228
rect 9706 8176 9758 8228
rect 9770 8176 9822 8228
rect 9834 8176 9886 8228
rect 9898 8176 9950 8228
rect 9962 8176 10014 8228
rect 10026 8176 10078 8228
rect 10090 8176 10142 8228
rect 10154 8176 10206 8228
rect 10218 8176 10270 8228
rect 10282 8176 10334 8228
rect 10346 8176 10398 8228
rect 10410 8176 10462 8228
rect 10474 8176 10526 8228
rect 10538 8176 10590 8228
rect 10602 8176 10654 8228
rect 10666 8176 10718 8228
rect 10730 8176 10782 8228
rect 10156 8000 10208 8052
rect 10220 8000 10272 8052
rect 8339 7751 8391 7803
rect 8403 7751 8455 7803
rect 8467 7751 8519 7803
rect 10771 7726 10823 7727
rect 10771 7692 10785 7726
rect 10785 7692 10819 7726
rect 10819 7692 10823 7726
rect 10771 7675 10823 7692
rect 10835 7675 10887 7727
rect 4362 6670 5246 6794
rect 2286 6470 2338 6522
rect 4362 6294 5246 6670
rect 6463 6643 6771 7015
rect 7318 7470 7370 7522
rect 7382 7470 7434 7522
rect 7446 7470 7498 7522
rect 7510 7470 7562 7522
rect 7574 7470 7626 7522
rect 7638 7470 7690 7522
rect 7702 7470 7754 7522
rect 7766 7470 7818 7522
rect 7830 7470 7882 7522
rect 7894 7470 7946 7522
rect 7958 7470 8010 7522
rect 8022 7470 8074 7522
rect 8086 7470 8138 7522
rect 8150 7470 8202 7522
rect 8214 7470 8266 7522
rect 8278 7470 8330 7522
rect 8647 7470 8699 7522
rect 8711 7470 8763 7522
rect 8775 7470 8827 7522
rect 8839 7470 8891 7522
rect 8903 7470 8955 7522
rect 8967 7470 9019 7522
rect 9031 7470 9083 7522
rect 9095 7470 9147 7522
rect 9159 7470 9211 7522
rect 9223 7470 9275 7522
rect 9287 7470 9339 7522
rect 9351 7470 9403 7522
rect 9415 7470 9467 7522
rect 9479 7470 9531 7522
rect 9543 7470 9595 7522
rect 9607 7470 9659 7522
rect 9671 7470 9723 7522
rect 9735 7470 9787 7522
rect 9799 7470 9851 7522
rect 9863 7470 9915 7522
rect 9927 7470 9979 7522
rect 9991 7470 10043 7522
rect 10055 7470 10107 7522
rect 10119 7470 10171 7522
rect 10183 7470 10235 7522
rect 10247 7470 10299 7522
rect 10311 7470 10363 7522
rect 10375 7470 10427 7522
rect 10439 7470 10491 7522
rect 10503 7470 10555 7522
rect 10567 7470 10619 7522
rect 7175 7153 8315 7269
rect 8626 7153 10726 7269
rect 8446 6870 8498 6871
rect 8446 6836 8455 6870
rect 8455 6836 8489 6870
rect 8489 6836 8498 6870
rect 8446 6819 8498 6836
rect 8446 6798 8498 6807
rect 8446 6764 8455 6798
rect 8455 6764 8489 6798
rect 8489 6764 8498 6798
rect 8446 6755 8498 6764
rect 8446 6726 8498 6743
rect 8446 6692 8455 6726
rect 8455 6692 8489 6726
rect 8489 6692 8498 6726
rect 10531 6773 10583 6825
rect 10595 6773 10647 6825
rect 8446 6691 8498 6692
rect 10248 6197 10300 6249
rect 10312 6197 10364 6249
rect 10376 6197 10428 6249
rect 10440 6197 10492 6249
rect 10504 6197 10556 6249
rect 10568 6197 10620 6249
rect 10632 6197 10684 6249
<< metal2 >>
rect 985 8286 7132 8287
rect 38 8261 7132 8286
rect 38 8209 60 8261
rect 112 8250 124 8261
rect 176 8250 188 8261
rect 240 8250 252 8261
rect 304 8250 316 8261
rect 368 8250 380 8261
rect 432 8250 444 8261
rect 496 8250 508 8261
rect 560 8250 572 8261
rect 624 8252 7132 8261
rect 624 8250 1057 8252
rect 1109 8250 1121 8252
rect 1173 8250 1185 8252
rect 1237 8250 1249 8252
rect 1301 8250 1313 8252
rect 1365 8250 1377 8252
rect 1429 8250 1441 8252
rect 1493 8250 1505 8252
rect 1557 8250 1569 8252
rect 1621 8250 1633 8252
rect 1685 8250 1697 8252
rect 1749 8250 1761 8252
rect 1813 8250 1825 8252
rect 1877 8250 1889 8252
rect 1941 8250 1953 8252
rect 2005 8250 2017 8252
rect 2069 8250 2081 8252
rect 2133 8250 2145 8252
rect 2197 8250 2209 8252
rect 2261 8250 2273 8252
rect 2325 8250 2337 8252
rect 2389 8250 2401 8252
rect 2453 8250 2465 8252
rect 2517 8250 2529 8252
rect 2581 8250 2593 8252
rect 2645 8250 2657 8252
rect 2709 8250 2721 8252
rect 2773 8250 2785 8252
rect 2837 8250 2849 8252
rect 2901 8250 2913 8252
rect 2965 8250 2977 8252
rect 3029 8250 3041 8252
rect 3093 8250 3105 8252
rect 3157 8250 3169 8252
rect 3221 8250 3233 8252
rect 3285 8250 3297 8252
rect 3349 8250 3361 8252
rect 3413 8250 3425 8252
rect 3477 8250 3489 8252
rect 3541 8250 3553 8252
rect 3605 8250 3617 8252
rect 3669 8250 3681 8252
rect 3733 8250 3745 8252
rect 3797 8250 3809 8252
rect 3861 8250 3873 8252
rect 3925 8250 3937 8252
rect 3989 8250 4001 8252
rect 4053 8250 4065 8252
rect 4117 8250 4129 8252
rect 4181 8250 4193 8252
rect 4245 8250 4257 8252
rect 4309 8250 4321 8252
rect 4373 8250 4385 8252
rect 4437 8250 4449 8252
rect 4501 8250 4513 8252
rect 4565 8250 4577 8252
rect 4629 8250 4641 8252
rect 4693 8250 4705 8252
rect 4757 8250 4769 8252
rect 4821 8250 4833 8252
rect 4885 8250 4897 8252
rect 4949 8250 4961 8252
rect 5013 8250 5025 8252
rect 5077 8250 5089 8252
rect 5141 8250 5153 8252
rect 5205 8250 5217 8252
rect 5269 8250 5281 8252
rect 5333 8250 5345 8252
rect 5397 8250 5409 8252
rect 5461 8250 5473 8252
rect 5525 8250 5537 8252
rect 5589 8250 5601 8252
rect 5653 8250 5665 8252
rect 5717 8250 5729 8252
rect 5781 8250 5793 8252
rect 5845 8250 5857 8252
rect 5909 8250 5921 8252
rect 5973 8250 5985 8252
rect 6037 8250 6049 8252
rect 6101 8250 6113 8252
rect 6165 8250 6177 8252
rect 6229 8250 6241 8252
rect 6293 8250 6305 8252
rect 6357 8250 6369 8252
rect 6421 8250 6433 8252
rect 6485 8250 6497 8252
rect 6549 8250 6561 8252
rect 6613 8250 6625 8252
rect 6677 8250 6689 8252
rect 6741 8250 6753 8252
rect 6805 8250 6817 8252
rect 6869 8250 6881 8252
rect 6933 8250 6945 8252
rect 6997 8250 7009 8252
rect 624 8209 920 8250
rect 38 8114 87 8209
rect 623 8187 920 8209
rect 7061 8200 7132 8252
rect 623 8114 654 8187
rect 38 8061 654 8114
rect 719 8139 801 8154
rect 719 8087 734 8139
rect 786 8087 801 8139
rect 719 8072 801 8087
rect 866 8114 920 8187
rect 7056 8114 7132 8200
rect 7284 8230 10841 8278
rect 7284 8228 7352 8230
rect 7408 8228 7432 8230
rect 7488 8228 7512 8230
rect 7568 8228 7592 8230
rect 7648 8228 7672 8230
rect 7728 8228 7752 8230
rect 7808 8228 7832 8230
rect 7888 8228 7912 8230
rect 7968 8228 7992 8230
rect 8048 8228 8072 8230
rect 8128 8228 8152 8230
rect 8208 8228 8232 8230
rect 8288 8228 8312 8230
rect 8368 8228 8392 8230
rect 8448 8228 8472 8230
rect 8528 8228 8552 8230
rect 8608 8228 8632 8230
rect 8688 8228 8712 8230
rect 8768 8228 8792 8230
rect 8848 8228 8872 8230
rect 8928 8228 8952 8230
rect 9008 8228 9032 8230
rect 9088 8228 9112 8230
rect 9168 8228 9192 8230
rect 9248 8228 9272 8230
rect 9328 8228 9352 8230
rect 9408 8228 9432 8230
rect 9488 8228 9512 8230
rect 9568 8228 9592 8230
rect 9648 8228 9672 8230
rect 9728 8228 9752 8230
rect 9808 8228 9832 8230
rect 9888 8228 9912 8230
rect 9968 8228 9992 8230
rect 10048 8228 10072 8230
rect 10128 8228 10152 8230
rect 10208 8228 10232 8230
rect 10288 8228 10312 8230
rect 10368 8228 10392 8230
rect 10448 8228 10472 8230
rect 10528 8228 10552 8230
rect 10608 8228 10632 8230
rect 10688 8228 10712 8230
rect 10768 8228 10841 8230
rect 7284 8176 7338 8228
rect 7582 8176 7592 8228
rect 7648 8176 7658 8228
rect 7902 8176 7912 8228
rect 7968 8176 7978 8228
rect 8222 8176 8232 8228
rect 8288 8176 8298 8228
rect 8542 8176 8552 8228
rect 8608 8176 8618 8228
rect 8862 8176 8872 8228
rect 8928 8176 8938 8228
rect 9182 8176 9192 8228
rect 9248 8176 9258 8228
rect 9502 8176 9512 8228
rect 9568 8176 9578 8228
rect 9822 8176 9832 8228
rect 9888 8176 9898 8228
rect 10142 8176 10152 8228
rect 10208 8176 10218 8228
rect 10462 8176 10472 8228
rect 10528 8176 10538 8228
rect 10782 8176 10841 8228
rect 7284 8174 7352 8176
rect 7408 8174 7432 8176
rect 7488 8174 7512 8176
rect 7568 8174 7592 8176
rect 7648 8174 7672 8176
rect 7728 8174 7752 8176
rect 7808 8174 7832 8176
rect 7888 8174 7912 8176
rect 7968 8174 7992 8176
rect 8048 8174 8072 8176
rect 8128 8174 8152 8176
rect 8208 8174 8232 8176
rect 8288 8174 8312 8176
rect 8368 8174 8392 8176
rect 8448 8174 8472 8176
rect 8528 8174 8552 8176
rect 8608 8174 8632 8176
rect 8688 8174 8712 8176
rect 8768 8174 8792 8176
rect 8848 8174 8872 8176
rect 8928 8174 8952 8176
rect 9008 8174 9032 8176
rect 9088 8174 9112 8176
rect 9168 8174 9192 8176
rect 9248 8174 9272 8176
rect 9328 8174 9352 8176
rect 9408 8174 9432 8176
rect 9488 8174 9512 8176
rect 9568 8174 9592 8176
rect 9648 8174 9672 8176
rect 9728 8174 9752 8176
rect 9808 8174 9832 8176
rect 9888 8174 9912 8176
rect 9968 8174 9992 8176
rect 10048 8174 10072 8176
rect 10128 8174 10152 8176
rect 10208 8174 10232 8176
rect 10288 8174 10312 8176
rect 10368 8174 10392 8176
rect 10448 8174 10472 8176
rect 10528 8174 10552 8176
rect 10608 8174 10632 8176
rect 10688 8174 10712 8176
rect 10768 8174 10841 8176
rect 7284 8125 10841 8174
rect 729 7616 785 8072
rect 866 8060 7132 8114
rect 10138 8054 10290 8066
rect 10138 7998 10146 8054
rect 10202 8052 10226 8054
rect 10208 8000 10220 8052
rect 10202 7998 10226 8000
rect 10282 7998 10290 8054
rect 10138 7986 10290 7998
rect 8339 7803 8519 7817
rect 8391 7751 8403 7803
rect 8455 7751 8467 7803
rect 8339 7738 8519 7751
rect 719 7601 801 7616
rect 719 7549 734 7601
rect 786 7549 801 7601
rect 719 7534 801 7549
rect 7279 7524 8374 7570
rect 7279 7468 7316 7524
rect 7372 7522 7396 7524
rect 7452 7522 7476 7524
rect 7532 7522 7556 7524
rect 7612 7522 7636 7524
rect 7692 7522 7716 7524
rect 7772 7522 7796 7524
rect 7852 7522 7876 7524
rect 7932 7522 7956 7524
rect 8012 7522 8036 7524
rect 8092 7522 8116 7524
rect 8172 7522 8196 7524
rect 8252 7522 8276 7524
rect 7372 7470 7382 7522
rect 7626 7470 7636 7522
rect 7692 7470 7702 7522
rect 7946 7470 7956 7522
rect 8012 7470 8022 7522
rect 8266 7470 8276 7522
rect 7372 7468 7396 7470
rect 7452 7468 7476 7470
rect 7532 7468 7556 7470
rect 7612 7468 7636 7470
rect 7692 7468 7716 7470
rect 7772 7468 7796 7470
rect 7852 7468 7876 7470
rect 7932 7468 7956 7470
rect 8012 7468 8036 7470
rect 8092 7468 8116 7470
rect 8172 7468 8196 7470
rect 8252 7468 8276 7470
rect 8332 7468 8374 7524
rect 7279 7417 8374 7468
rect 7141 7269 8355 7324
rect 7141 7153 7175 7269
rect 8315 7153 8355 7269
rect 7141 7094 8355 7153
rect 2275 7064 2351 7084
rect 2275 7012 2287 7064
rect 2339 7012 2351 7064
rect 2275 6993 2351 7012
rect 6407 7017 6825 7065
rect 6407 7015 6469 7017
rect 6765 7015 6825 7017
rect 2288 6543 2340 6993
rect 4308 6833 5298 6868
rect 2275 6522 2350 6543
rect 2275 6470 2286 6522
rect 2338 6470 2350 6522
rect 2275 6450 2350 6470
rect 4308 6537 4336 6833
rect 5272 6537 5298 6833
rect 6407 6643 6463 7015
rect 6771 6643 6825 7015
rect 8443 6888 8500 7738
rect 10753 7729 10905 7741
rect 10753 7673 10761 7729
rect 10817 7727 10841 7729
rect 10823 7675 10835 7727
rect 10817 7673 10841 7675
rect 10897 7673 10905 7729
rect 10753 7661 10905 7673
rect 8588 7543 10667 7570
rect 8587 7524 10667 7543
rect 8587 7468 8645 7524
rect 8701 7522 8725 7524
rect 8781 7522 8805 7524
rect 8861 7522 8885 7524
rect 8941 7522 8965 7524
rect 9021 7522 9045 7524
rect 9101 7522 9125 7524
rect 9181 7522 9205 7524
rect 9261 7522 9285 7524
rect 9341 7522 9365 7524
rect 9421 7522 9445 7524
rect 9501 7522 9525 7524
rect 9581 7522 9605 7524
rect 9661 7522 9685 7524
rect 9741 7522 9765 7524
rect 9821 7522 9845 7524
rect 9901 7522 9925 7524
rect 9981 7522 10005 7524
rect 10061 7522 10085 7524
rect 10141 7522 10165 7524
rect 10221 7522 10245 7524
rect 10301 7522 10325 7524
rect 10381 7522 10405 7524
rect 10461 7522 10485 7524
rect 10541 7522 10565 7524
rect 8701 7470 8711 7522
rect 8955 7470 8965 7522
rect 9021 7470 9031 7522
rect 9275 7470 9285 7522
rect 9341 7470 9351 7522
rect 9595 7470 9605 7522
rect 9661 7470 9671 7522
rect 9915 7470 9925 7522
rect 9981 7470 9991 7522
rect 10235 7470 10245 7522
rect 10301 7470 10311 7522
rect 10555 7470 10565 7522
rect 8701 7468 8725 7470
rect 8781 7468 8805 7470
rect 8861 7468 8885 7470
rect 8941 7468 8965 7470
rect 9021 7468 9045 7470
rect 9101 7468 9125 7470
rect 9181 7468 9205 7470
rect 9261 7468 9285 7470
rect 9341 7468 9365 7470
rect 9421 7468 9445 7470
rect 9501 7468 9525 7470
rect 9581 7468 9605 7470
rect 9661 7468 9685 7470
rect 9741 7468 9765 7470
rect 9821 7468 9845 7470
rect 9901 7468 9925 7470
rect 9981 7468 10005 7470
rect 10061 7468 10085 7470
rect 10141 7468 10165 7470
rect 10221 7468 10245 7470
rect 10301 7468 10325 7470
rect 10381 7468 10405 7470
rect 10461 7468 10485 7470
rect 10541 7468 10565 7470
rect 10621 7468 10667 7524
rect 8587 7449 10667 7468
rect 8588 7417 10667 7449
rect 8567 7269 10798 7324
rect 8567 7153 8626 7269
rect 10726 7153 10798 7269
rect 8567 7094 10798 7153
rect 8439 6871 8506 6888
rect 8439 6819 8446 6871
rect 8498 6819 8506 6871
rect 8439 6807 8506 6819
rect 8439 6755 8446 6807
rect 8498 6755 8506 6807
rect 8439 6743 8506 6755
rect 8439 6691 8446 6743
rect 8498 6691 8506 6743
rect 8439 6674 8506 6691
rect 6407 6641 6469 6643
rect 6765 6641 6825 6643
rect 6407 6600 6825 6641
rect 4308 6294 4362 6537
rect 5246 6294 5298 6537
rect 4308 6249 5298 6294
rect 10221 6270 10431 7094
rect 10498 6827 10918 6834
rect 10498 6825 10765 6827
rect 10498 6773 10531 6825
rect 10583 6773 10595 6825
rect 10647 6773 10765 6825
rect 10498 6771 10765 6773
rect 10821 6771 10845 6827
rect 10901 6771 10918 6827
rect 10498 6765 10918 6771
rect 10221 6249 10716 6270
rect 10221 6197 10248 6249
rect 10300 6197 10312 6249
rect 10364 6197 10376 6249
rect 10428 6197 10440 6249
rect 10492 6197 10504 6249
rect 10556 6197 10568 6249
rect 10620 6197 10632 6249
rect 10684 6197 10716 6249
rect 10221 6176 10716 6197
<< via2 >>
rect 87 8209 112 8250
rect 112 8209 124 8250
rect 124 8209 176 8250
rect 176 8209 188 8250
rect 188 8209 240 8250
rect 240 8209 252 8250
rect 252 8209 304 8250
rect 304 8209 316 8250
rect 316 8209 368 8250
rect 368 8209 380 8250
rect 380 8209 432 8250
rect 432 8209 444 8250
rect 444 8209 496 8250
rect 496 8209 508 8250
rect 508 8209 560 8250
rect 560 8209 572 8250
rect 572 8209 623 8250
rect 87 8114 623 8209
rect 920 8200 1057 8250
rect 1057 8200 1109 8250
rect 1109 8200 1121 8250
rect 1121 8200 1173 8250
rect 1173 8200 1185 8250
rect 1185 8200 1237 8250
rect 1237 8200 1249 8250
rect 1249 8200 1301 8250
rect 1301 8200 1313 8250
rect 1313 8200 1365 8250
rect 1365 8200 1377 8250
rect 1377 8200 1429 8250
rect 1429 8200 1441 8250
rect 1441 8200 1493 8250
rect 1493 8200 1505 8250
rect 1505 8200 1557 8250
rect 1557 8200 1569 8250
rect 1569 8200 1621 8250
rect 1621 8200 1633 8250
rect 1633 8200 1685 8250
rect 1685 8200 1697 8250
rect 1697 8200 1749 8250
rect 1749 8200 1761 8250
rect 1761 8200 1813 8250
rect 1813 8200 1825 8250
rect 1825 8200 1877 8250
rect 1877 8200 1889 8250
rect 1889 8200 1941 8250
rect 1941 8200 1953 8250
rect 1953 8200 2005 8250
rect 2005 8200 2017 8250
rect 2017 8200 2069 8250
rect 2069 8200 2081 8250
rect 2081 8200 2133 8250
rect 2133 8200 2145 8250
rect 2145 8200 2197 8250
rect 2197 8200 2209 8250
rect 2209 8200 2261 8250
rect 2261 8200 2273 8250
rect 2273 8200 2325 8250
rect 2325 8200 2337 8250
rect 2337 8200 2389 8250
rect 2389 8200 2401 8250
rect 2401 8200 2453 8250
rect 2453 8200 2465 8250
rect 2465 8200 2517 8250
rect 2517 8200 2529 8250
rect 2529 8200 2581 8250
rect 2581 8200 2593 8250
rect 2593 8200 2645 8250
rect 2645 8200 2657 8250
rect 2657 8200 2709 8250
rect 2709 8200 2721 8250
rect 2721 8200 2773 8250
rect 2773 8200 2785 8250
rect 2785 8200 2837 8250
rect 2837 8200 2849 8250
rect 2849 8200 2901 8250
rect 2901 8200 2913 8250
rect 2913 8200 2965 8250
rect 2965 8200 2977 8250
rect 2977 8200 3029 8250
rect 3029 8200 3041 8250
rect 3041 8200 3093 8250
rect 3093 8200 3105 8250
rect 3105 8200 3157 8250
rect 3157 8200 3169 8250
rect 3169 8200 3221 8250
rect 3221 8200 3233 8250
rect 3233 8200 3285 8250
rect 3285 8200 3297 8250
rect 3297 8200 3349 8250
rect 3349 8200 3361 8250
rect 3361 8200 3413 8250
rect 3413 8200 3425 8250
rect 3425 8200 3477 8250
rect 3477 8200 3489 8250
rect 3489 8200 3541 8250
rect 3541 8200 3553 8250
rect 3553 8200 3605 8250
rect 3605 8200 3617 8250
rect 3617 8200 3669 8250
rect 3669 8200 3681 8250
rect 3681 8200 3733 8250
rect 3733 8200 3745 8250
rect 3745 8200 3797 8250
rect 3797 8200 3809 8250
rect 3809 8200 3861 8250
rect 3861 8200 3873 8250
rect 3873 8200 3925 8250
rect 3925 8200 3937 8250
rect 3937 8200 3989 8250
rect 3989 8200 4001 8250
rect 4001 8200 4053 8250
rect 4053 8200 4065 8250
rect 4065 8200 4117 8250
rect 4117 8200 4129 8250
rect 4129 8200 4181 8250
rect 4181 8200 4193 8250
rect 4193 8200 4245 8250
rect 4245 8200 4257 8250
rect 4257 8200 4309 8250
rect 4309 8200 4321 8250
rect 4321 8200 4373 8250
rect 4373 8200 4385 8250
rect 4385 8200 4437 8250
rect 4437 8200 4449 8250
rect 4449 8200 4501 8250
rect 4501 8200 4513 8250
rect 4513 8200 4565 8250
rect 4565 8200 4577 8250
rect 4577 8200 4629 8250
rect 4629 8200 4641 8250
rect 4641 8200 4693 8250
rect 4693 8200 4705 8250
rect 4705 8200 4757 8250
rect 4757 8200 4769 8250
rect 4769 8200 4821 8250
rect 4821 8200 4833 8250
rect 4833 8200 4885 8250
rect 4885 8200 4897 8250
rect 4897 8200 4949 8250
rect 4949 8200 4961 8250
rect 4961 8200 5013 8250
rect 5013 8200 5025 8250
rect 5025 8200 5077 8250
rect 5077 8200 5089 8250
rect 5089 8200 5141 8250
rect 5141 8200 5153 8250
rect 5153 8200 5205 8250
rect 5205 8200 5217 8250
rect 5217 8200 5269 8250
rect 5269 8200 5281 8250
rect 5281 8200 5333 8250
rect 5333 8200 5345 8250
rect 5345 8200 5397 8250
rect 5397 8200 5409 8250
rect 5409 8200 5461 8250
rect 5461 8200 5473 8250
rect 5473 8200 5525 8250
rect 5525 8200 5537 8250
rect 5537 8200 5589 8250
rect 5589 8200 5601 8250
rect 5601 8200 5653 8250
rect 5653 8200 5665 8250
rect 5665 8200 5717 8250
rect 5717 8200 5729 8250
rect 5729 8200 5781 8250
rect 5781 8200 5793 8250
rect 5793 8200 5845 8250
rect 5845 8200 5857 8250
rect 5857 8200 5909 8250
rect 5909 8200 5921 8250
rect 5921 8200 5973 8250
rect 5973 8200 5985 8250
rect 5985 8200 6037 8250
rect 6037 8200 6049 8250
rect 6049 8200 6101 8250
rect 6101 8200 6113 8250
rect 6113 8200 6165 8250
rect 6165 8200 6177 8250
rect 6177 8200 6229 8250
rect 6229 8200 6241 8250
rect 6241 8200 6293 8250
rect 6293 8200 6305 8250
rect 6305 8200 6357 8250
rect 6357 8200 6369 8250
rect 6369 8200 6421 8250
rect 6421 8200 6433 8250
rect 6433 8200 6485 8250
rect 6485 8200 6497 8250
rect 6497 8200 6549 8250
rect 6549 8200 6561 8250
rect 6561 8200 6613 8250
rect 6613 8200 6625 8250
rect 6625 8200 6677 8250
rect 6677 8200 6689 8250
rect 6689 8200 6741 8250
rect 6741 8200 6753 8250
rect 6753 8200 6805 8250
rect 6805 8200 6817 8250
rect 6817 8200 6869 8250
rect 6869 8200 6881 8250
rect 6881 8200 6933 8250
rect 6933 8200 6945 8250
rect 6945 8200 6997 8250
rect 6997 8200 7009 8250
rect 7009 8200 7056 8250
rect 920 8114 7056 8200
rect 7352 8228 7408 8230
rect 7432 8228 7488 8230
rect 7512 8228 7568 8230
rect 7592 8228 7648 8230
rect 7672 8228 7728 8230
rect 7752 8228 7808 8230
rect 7832 8228 7888 8230
rect 7912 8228 7968 8230
rect 7992 8228 8048 8230
rect 8072 8228 8128 8230
rect 8152 8228 8208 8230
rect 8232 8228 8288 8230
rect 8312 8228 8368 8230
rect 8392 8228 8448 8230
rect 8472 8228 8528 8230
rect 8552 8228 8608 8230
rect 8632 8228 8688 8230
rect 8712 8228 8768 8230
rect 8792 8228 8848 8230
rect 8872 8228 8928 8230
rect 8952 8228 9008 8230
rect 9032 8228 9088 8230
rect 9112 8228 9168 8230
rect 9192 8228 9248 8230
rect 9272 8228 9328 8230
rect 9352 8228 9408 8230
rect 9432 8228 9488 8230
rect 9512 8228 9568 8230
rect 9592 8228 9648 8230
rect 9672 8228 9728 8230
rect 9752 8228 9808 8230
rect 9832 8228 9888 8230
rect 9912 8228 9968 8230
rect 9992 8228 10048 8230
rect 10072 8228 10128 8230
rect 10152 8228 10208 8230
rect 10232 8228 10288 8230
rect 10312 8228 10368 8230
rect 10392 8228 10448 8230
rect 10472 8228 10528 8230
rect 10552 8228 10608 8230
rect 10632 8228 10688 8230
rect 10712 8228 10768 8230
rect 7352 8176 7390 8228
rect 7390 8176 7402 8228
rect 7402 8176 7408 8228
rect 7432 8176 7454 8228
rect 7454 8176 7466 8228
rect 7466 8176 7488 8228
rect 7512 8176 7518 8228
rect 7518 8176 7530 8228
rect 7530 8176 7568 8228
rect 7592 8176 7594 8228
rect 7594 8176 7646 8228
rect 7646 8176 7648 8228
rect 7672 8176 7710 8228
rect 7710 8176 7722 8228
rect 7722 8176 7728 8228
rect 7752 8176 7774 8228
rect 7774 8176 7786 8228
rect 7786 8176 7808 8228
rect 7832 8176 7838 8228
rect 7838 8176 7850 8228
rect 7850 8176 7888 8228
rect 7912 8176 7914 8228
rect 7914 8176 7966 8228
rect 7966 8176 7968 8228
rect 7992 8176 8030 8228
rect 8030 8176 8042 8228
rect 8042 8176 8048 8228
rect 8072 8176 8094 8228
rect 8094 8176 8106 8228
rect 8106 8176 8128 8228
rect 8152 8176 8158 8228
rect 8158 8176 8170 8228
rect 8170 8176 8208 8228
rect 8232 8176 8234 8228
rect 8234 8176 8286 8228
rect 8286 8176 8288 8228
rect 8312 8176 8350 8228
rect 8350 8176 8362 8228
rect 8362 8176 8368 8228
rect 8392 8176 8414 8228
rect 8414 8176 8426 8228
rect 8426 8176 8448 8228
rect 8472 8176 8478 8228
rect 8478 8176 8490 8228
rect 8490 8176 8528 8228
rect 8552 8176 8554 8228
rect 8554 8176 8606 8228
rect 8606 8176 8608 8228
rect 8632 8176 8670 8228
rect 8670 8176 8682 8228
rect 8682 8176 8688 8228
rect 8712 8176 8734 8228
rect 8734 8176 8746 8228
rect 8746 8176 8768 8228
rect 8792 8176 8798 8228
rect 8798 8176 8810 8228
rect 8810 8176 8848 8228
rect 8872 8176 8874 8228
rect 8874 8176 8926 8228
rect 8926 8176 8928 8228
rect 8952 8176 8990 8228
rect 8990 8176 9002 8228
rect 9002 8176 9008 8228
rect 9032 8176 9054 8228
rect 9054 8176 9066 8228
rect 9066 8176 9088 8228
rect 9112 8176 9118 8228
rect 9118 8176 9130 8228
rect 9130 8176 9168 8228
rect 9192 8176 9194 8228
rect 9194 8176 9246 8228
rect 9246 8176 9248 8228
rect 9272 8176 9310 8228
rect 9310 8176 9322 8228
rect 9322 8176 9328 8228
rect 9352 8176 9374 8228
rect 9374 8176 9386 8228
rect 9386 8176 9408 8228
rect 9432 8176 9438 8228
rect 9438 8176 9450 8228
rect 9450 8176 9488 8228
rect 9512 8176 9514 8228
rect 9514 8176 9566 8228
rect 9566 8176 9568 8228
rect 9592 8176 9630 8228
rect 9630 8176 9642 8228
rect 9642 8176 9648 8228
rect 9672 8176 9694 8228
rect 9694 8176 9706 8228
rect 9706 8176 9728 8228
rect 9752 8176 9758 8228
rect 9758 8176 9770 8228
rect 9770 8176 9808 8228
rect 9832 8176 9834 8228
rect 9834 8176 9886 8228
rect 9886 8176 9888 8228
rect 9912 8176 9950 8228
rect 9950 8176 9962 8228
rect 9962 8176 9968 8228
rect 9992 8176 10014 8228
rect 10014 8176 10026 8228
rect 10026 8176 10048 8228
rect 10072 8176 10078 8228
rect 10078 8176 10090 8228
rect 10090 8176 10128 8228
rect 10152 8176 10154 8228
rect 10154 8176 10206 8228
rect 10206 8176 10208 8228
rect 10232 8176 10270 8228
rect 10270 8176 10282 8228
rect 10282 8176 10288 8228
rect 10312 8176 10334 8228
rect 10334 8176 10346 8228
rect 10346 8176 10368 8228
rect 10392 8176 10398 8228
rect 10398 8176 10410 8228
rect 10410 8176 10448 8228
rect 10472 8176 10474 8228
rect 10474 8176 10526 8228
rect 10526 8176 10528 8228
rect 10552 8176 10590 8228
rect 10590 8176 10602 8228
rect 10602 8176 10608 8228
rect 10632 8176 10654 8228
rect 10654 8176 10666 8228
rect 10666 8176 10688 8228
rect 10712 8176 10718 8228
rect 10718 8176 10730 8228
rect 10730 8176 10768 8228
rect 7352 8174 7408 8176
rect 7432 8174 7488 8176
rect 7512 8174 7568 8176
rect 7592 8174 7648 8176
rect 7672 8174 7728 8176
rect 7752 8174 7808 8176
rect 7832 8174 7888 8176
rect 7912 8174 7968 8176
rect 7992 8174 8048 8176
rect 8072 8174 8128 8176
rect 8152 8174 8208 8176
rect 8232 8174 8288 8176
rect 8312 8174 8368 8176
rect 8392 8174 8448 8176
rect 8472 8174 8528 8176
rect 8552 8174 8608 8176
rect 8632 8174 8688 8176
rect 8712 8174 8768 8176
rect 8792 8174 8848 8176
rect 8872 8174 8928 8176
rect 8952 8174 9008 8176
rect 9032 8174 9088 8176
rect 9112 8174 9168 8176
rect 9192 8174 9248 8176
rect 9272 8174 9328 8176
rect 9352 8174 9408 8176
rect 9432 8174 9488 8176
rect 9512 8174 9568 8176
rect 9592 8174 9648 8176
rect 9672 8174 9728 8176
rect 9752 8174 9808 8176
rect 9832 8174 9888 8176
rect 9912 8174 9968 8176
rect 9992 8174 10048 8176
rect 10072 8174 10128 8176
rect 10152 8174 10208 8176
rect 10232 8174 10288 8176
rect 10312 8174 10368 8176
rect 10392 8174 10448 8176
rect 10472 8174 10528 8176
rect 10552 8174 10608 8176
rect 10632 8174 10688 8176
rect 10712 8174 10768 8176
rect 10146 8052 10202 8054
rect 10226 8052 10282 8054
rect 10146 8000 10156 8052
rect 10156 8000 10202 8052
rect 10226 8000 10272 8052
rect 10272 8000 10282 8052
rect 10146 7998 10202 8000
rect 10226 7998 10282 8000
rect 7316 7522 7372 7524
rect 7396 7522 7452 7524
rect 7476 7522 7532 7524
rect 7556 7522 7612 7524
rect 7636 7522 7692 7524
rect 7716 7522 7772 7524
rect 7796 7522 7852 7524
rect 7876 7522 7932 7524
rect 7956 7522 8012 7524
rect 8036 7522 8092 7524
rect 8116 7522 8172 7524
rect 8196 7522 8252 7524
rect 8276 7522 8332 7524
rect 7316 7470 7318 7522
rect 7318 7470 7370 7522
rect 7370 7470 7372 7522
rect 7396 7470 7434 7522
rect 7434 7470 7446 7522
rect 7446 7470 7452 7522
rect 7476 7470 7498 7522
rect 7498 7470 7510 7522
rect 7510 7470 7532 7522
rect 7556 7470 7562 7522
rect 7562 7470 7574 7522
rect 7574 7470 7612 7522
rect 7636 7470 7638 7522
rect 7638 7470 7690 7522
rect 7690 7470 7692 7522
rect 7716 7470 7754 7522
rect 7754 7470 7766 7522
rect 7766 7470 7772 7522
rect 7796 7470 7818 7522
rect 7818 7470 7830 7522
rect 7830 7470 7852 7522
rect 7876 7470 7882 7522
rect 7882 7470 7894 7522
rect 7894 7470 7932 7522
rect 7956 7470 7958 7522
rect 7958 7470 8010 7522
rect 8010 7470 8012 7522
rect 8036 7470 8074 7522
rect 8074 7470 8086 7522
rect 8086 7470 8092 7522
rect 8116 7470 8138 7522
rect 8138 7470 8150 7522
rect 8150 7470 8172 7522
rect 8196 7470 8202 7522
rect 8202 7470 8214 7522
rect 8214 7470 8252 7522
rect 8276 7470 8278 7522
rect 8278 7470 8330 7522
rect 8330 7470 8332 7522
rect 7316 7468 7372 7470
rect 7396 7468 7452 7470
rect 7476 7468 7532 7470
rect 7556 7468 7612 7470
rect 7636 7468 7692 7470
rect 7716 7468 7772 7470
rect 7796 7468 7852 7470
rect 7876 7468 7932 7470
rect 7956 7468 8012 7470
rect 8036 7468 8092 7470
rect 8116 7468 8172 7470
rect 8196 7468 8252 7470
rect 8276 7468 8332 7470
rect 6469 7015 6765 7017
rect 4336 6794 5272 6833
rect 4336 6537 4362 6794
rect 4362 6537 5246 6794
rect 5246 6537 5272 6794
rect 6469 6643 6765 7015
rect 10761 7727 10817 7729
rect 10841 7727 10897 7729
rect 10761 7675 10771 7727
rect 10771 7675 10817 7727
rect 10841 7675 10887 7727
rect 10887 7675 10897 7727
rect 10761 7673 10817 7675
rect 10841 7673 10897 7675
rect 8645 7522 8701 7524
rect 8725 7522 8781 7524
rect 8805 7522 8861 7524
rect 8885 7522 8941 7524
rect 8965 7522 9021 7524
rect 9045 7522 9101 7524
rect 9125 7522 9181 7524
rect 9205 7522 9261 7524
rect 9285 7522 9341 7524
rect 9365 7522 9421 7524
rect 9445 7522 9501 7524
rect 9525 7522 9581 7524
rect 9605 7522 9661 7524
rect 9685 7522 9741 7524
rect 9765 7522 9821 7524
rect 9845 7522 9901 7524
rect 9925 7522 9981 7524
rect 10005 7522 10061 7524
rect 10085 7522 10141 7524
rect 10165 7522 10221 7524
rect 10245 7522 10301 7524
rect 10325 7522 10381 7524
rect 10405 7522 10461 7524
rect 10485 7522 10541 7524
rect 10565 7522 10621 7524
rect 8645 7470 8647 7522
rect 8647 7470 8699 7522
rect 8699 7470 8701 7522
rect 8725 7470 8763 7522
rect 8763 7470 8775 7522
rect 8775 7470 8781 7522
rect 8805 7470 8827 7522
rect 8827 7470 8839 7522
rect 8839 7470 8861 7522
rect 8885 7470 8891 7522
rect 8891 7470 8903 7522
rect 8903 7470 8941 7522
rect 8965 7470 8967 7522
rect 8967 7470 9019 7522
rect 9019 7470 9021 7522
rect 9045 7470 9083 7522
rect 9083 7470 9095 7522
rect 9095 7470 9101 7522
rect 9125 7470 9147 7522
rect 9147 7470 9159 7522
rect 9159 7470 9181 7522
rect 9205 7470 9211 7522
rect 9211 7470 9223 7522
rect 9223 7470 9261 7522
rect 9285 7470 9287 7522
rect 9287 7470 9339 7522
rect 9339 7470 9341 7522
rect 9365 7470 9403 7522
rect 9403 7470 9415 7522
rect 9415 7470 9421 7522
rect 9445 7470 9467 7522
rect 9467 7470 9479 7522
rect 9479 7470 9501 7522
rect 9525 7470 9531 7522
rect 9531 7470 9543 7522
rect 9543 7470 9581 7522
rect 9605 7470 9607 7522
rect 9607 7470 9659 7522
rect 9659 7470 9661 7522
rect 9685 7470 9723 7522
rect 9723 7470 9735 7522
rect 9735 7470 9741 7522
rect 9765 7470 9787 7522
rect 9787 7470 9799 7522
rect 9799 7470 9821 7522
rect 9845 7470 9851 7522
rect 9851 7470 9863 7522
rect 9863 7470 9901 7522
rect 9925 7470 9927 7522
rect 9927 7470 9979 7522
rect 9979 7470 9981 7522
rect 10005 7470 10043 7522
rect 10043 7470 10055 7522
rect 10055 7470 10061 7522
rect 10085 7470 10107 7522
rect 10107 7470 10119 7522
rect 10119 7470 10141 7522
rect 10165 7470 10171 7522
rect 10171 7470 10183 7522
rect 10183 7470 10221 7522
rect 10245 7470 10247 7522
rect 10247 7470 10299 7522
rect 10299 7470 10301 7522
rect 10325 7470 10363 7522
rect 10363 7470 10375 7522
rect 10375 7470 10381 7522
rect 10405 7470 10427 7522
rect 10427 7470 10439 7522
rect 10439 7470 10461 7522
rect 10485 7470 10491 7522
rect 10491 7470 10503 7522
rect 10503 7470 10541 7522
rect 10565 7470 10567 7522
rect 10567 7470 10619 7522
rect 10619 7470 10621 7522
rect 8645 7468 8701 7470
rect 8725 7468 8781 7470
rect 8805 7468 8861 7470
rect 8885 7468 8941 7470
rect 8965 7468 9021 7470
rect 9045 7468 9101 7470
rect 9125 7468 9181 7470
rect 9205 7468 9261 7470
rect 9285 7468 9341 7470
rect 9365 7468 9421 7470
rect 9445 7468 9501 7470
rect 9525 7468 9581 7470
rect 9605 7468 9661 7470
rect 9685 7468 9741 7470
rect 9765 7468 9821 7470
rect 9845 7468 9901 7470
rect 9925 7468 9981 7470
rect 10005 7468 10061 7470
rect 10085 7468 10141 7470
rect 10165 7468 10221 7470
rect 10245 7468 10301 7470
rect 10325 7468 10381 7470
rect 10405 7468 10461 7470
rect 10485 7468 10541 7470
rect 10565 7468 10621 7470
rect 6469 6641 6765 6643
rect 10765 6771 10821 6827
rect 10845 6771 10901 6827
<< metal3 >>
rect 38 8250 7126 8283
rect 38 8114 87 8250
rect 623 8234 920 8250
rect 7056 8114 7126 8250
rect 7284 8234 10841 8278
rect 7284 8170 7348 8234
rect 7412 8170 7428 8234
rect 7492 8170 7508 8234
rect 7572 8170 7588 8234
rect 7652 8170 7668 8234
rect 7732 8170 7748 8234
rect 7812 8170 7828 8234
rect 7892 8170 7908 8234
rect 7972 8170 7988 8234
rect 8052 8170 8068 8234
rect 8132 8170 8148 8234
rect 8212 8170 8228 8234
rect 8292 8170 8308 8234
rect 8372 8170 8388 8234
rect 8452 8170 8468 8234
rect 8532 8170 8548 8234
rect 8612 8170 8628 8234
rect 8692 8170 8708 8234
rect 8772 8170 8788 8234
rect 8852 8170 8868 8234
rect 8932 8170 8948 8234
rect 9012 8170 9028 8234
rect 9092 8170 9108 8234
rect 9172 8170 9188 8234
rect 9252 8170 9268 8234
rect 9332 8170 9348 8234
rect 9412 8170 9428 8234
rect 9492 8170 9508 8234
rect 9572 8170 9588 8234
rect 9652 8170 9668 8234
rect 9732 8170 9748 8234
rect 9812 8170 9828 8234
rect 9892 8170 9908 8234
rect 9972 8170 9988 8234
rect 10052 8170 10068 8234
rect 10132 8170 10148 8234
rect 10212 8170 10228 8234
rect 10292 8170 10308 8234
rect 10372 8170 10388 8234
rect 10452 8170 10468 8234
rect 10532 8170 10548 8234
rect 10612 8170 10628 8234
rect 10692 8170 10708 8234
rect 10772 8170 10841 8234
rect 7284 8125 10841 8170
rect 38 8010 101 8114
rect 7045 8010 7126 8114
rect 38 7965 7126 8010
rect 10128 8056 10295 8064
rect 10128 8054 10431 8056
rect 10128 7998 10146 8054
rect 10202 7998 10226 8054
rect 10282 7998 10431 8054
rect 10128 7996 10431 7998
rect 10128 7991 10295 7996
rect 10371 7916 10431 7996
rect 10371 7856 11343 7916
rect 10743 7729 10910 7739
rect 10743 7673 10761 7729
rect 10817 7673 10841 7729
rect 10897 7673 10910 7729
rect 10743 7666 10910 7673
rect 7279 7528 10667 7570
rect 7279 7524 7345 7528
rect 7409 7524 7425 7528
rect 7489 7524 7505 7528
rect 7569 7524 7585 7528
rect 7649 7524 7665 7528
rect 7729 7524 7745 7528
rect 7809 7524 7825 7528
rect 7889 7524 7905 7528
rect 7969 7524 7985 7528
rect 8049 7524 8065 7528
rect 8129 7524 8145 7528
rect 8209 7524 8225 7528
rect 8289 7524 8305 7528
rect 7279 7468 7316 7524
rect 7279 7464 7345 7468
rect 7409 7464 7425 7468
rect 7489 7464 7505 7468
rect 7569 7464 7585 7468
rect 7649 7464 7665 7468
rect 7729 7464 7745 7468
rect 7809 7464 7825 7468
rect 7889 7464 7905 7468
rect 7969 7464 7985 7468
rect 8049 7464 8065 7468
rect 8129 7464 8145 7468
rect 8209 7464 8225 7468
rect 8289 7464 8305 7468
rect 8369 7464 8385 7528
rect 8449 7464 8465 7528
rect 8529 7464 8545 7528
rect 8609 7464 8625 7528
rect 8689 7524 8705 7528
rect 8769 7524 8785 7528
rect 8849 7524 8865 7528
rect 8929 7524 8945 7528
rect 9009 7524 9025 7528
rect 9089 7524 9105 7528
rect 9169 7524 9185 7528
rect 9249 7524 9265 7528
rect 9329 7524 9345 7528
rect 9409 7524 9425 7528
rect 9489 7524 9505 7528
rect 9569 7524 9585 7528
rect 9649 7524 9665 7528
rect 9729 7524 9745 7528
rect 9809 7524 9825 7528
rect 9889 7524 9905 7528
rect 9969 7524 9985 7528
rect 10049 7524 10065 7528
rect 10129 7524 10145 7528
rect 10209 7524 10225 7528
rect 10289 7524 10305 7528
rect 10369 7524 10385 7528
rect 10449 7524 10465 7528
rect 10529 7524 10545 7528
rect 10609 7524 10667 7528
rect 8701 7468 8705 7524
rect 8781 7468 8785 7524
rect 8861 7468 8865 7524
rect 8941 7468 8945 7524
rect 9021 7468 9025 7524
rect 9101 7468 9105 7524
rect 9181 7468 9185 7524
rect 9261 7468 9265 7524
rect 9341 7468 9345 7524
rect 9421 7468 9425 7524
rect 9501 7468 9505 7524
rect 9581 7468 9585 7524
rect 9661 7468 9665 7524
rect 9741 7468 9745 7524
rect 9821 7468 9825 7524
rect 9901 7468 9905 7524
rect 9981 7468 9985 7524
rect 10061 7468 10065 7524
rect 10141 7468 10145 7524
rect 10221 7468 10225 7524
rect 10301 7468 10305 7524
rect 10381 7468 10385 7524
rect 10461 7468 10465 7524
rect 10541 7468 10545 7524
rect 10621 7468 10667 7524
rect 10792 7551 10852 7666
rect 10792 7491 11344 7551
rect 8689 7464 8705 7468
rect 8769 7464 8785 7468
rect 8849 7464 8865 7468
rect 8929 7464 8945 7468
rect 9009 7464 9025 7468
rect 9089 7464 9105 7468
rect 9169 7464 9185 7468
rect 9249 7464 9265 7468
rect 9329 7464 9345 7468
rect 9409 7464 9425 7468
rect 9489 7464 9505 7468
rect 9569 7464 9585 7468
rect 9649 7464 9665 7468
rect 9729 7464 9745 7468
rect 9809 7464 9825 7468
rect 9889 7464 9905 7468
rect 9969 7464 9985 7468
rect 10049 7464 10065 7468
rect 10129 7464 10145 7468
rect 10209 7464 10225 7468
rect 10289 7464 10305 7468
rect 10369 7464 10385 7468
rect 10449 7464 10465 7468
rect 10529 7464 10545 7468
rect 10609 7464 10667 7468
rect 7279 7417 10667 7464
rect 4111 7269 5299 7317
rect 4111 6833 4377 7269
rect 5241 6833 5299 7269
rect 4111 6537 4336 6833
rect 5272 6537 5299 6833
rect 6408 7021 6825 7065
rect 6408 6637 6465 7021
rect 6769 6637 6825 7021
rect 10747 6834 10918 6840
rect 10747 6827 11342 6834
rect 10747 6771 10765 6827
rect 10821 6771 10845 6827
rect 10901 6771 11342 6827
rect 10747 6765 11342 6771
rect 10747 6758 10918 6765
rect 6408 6600 6825 6637
rect 4111 6494 5299 6537
rect 4111 6251 4307 6494
<< via3 >>
rect 101 8114 623 8234
rect 623 8114 920 8234
rect 920 8114 7045 8234
rect 7348 8230 7412 8234
rect 7348 8174 7352 8230
rect 7352 8174 7408 8230
rect 7408 8174 7412 8230
rect 7348 8170 7412 8174
rect 7428 8230 7492 8234
rect 7428 8174 7432 8230
rect 7432 8174 7488 8230
rect 7488 8174 7492 8230
rect 7428 8170 7492 8174
rect 7508 8230 7572 8234
rect 7508 8174 7512 8230
rect 7512 8174 7568 8230
rect 7568 8174 7572 8230
rect 7508 8170 7572 8174
rect 7588 8230 7652 8234
rect 7588 8174 7592 8230
rect 7592 8174 7648 8230
rect 7648 8174 7652 8230
rect 7588 8170 7652 8174
rect 7668 8230 7732 8234
rect 7668 8174 7672 8230
rect 7672 8174 7728 8230
rect 7728 8174 7732 8230
rect 7668 8170 7732 8174
rect 7748 8230 7812 8234
rect 7748 8174 7752 8230
rect 7752 8174 7808 8230
rect 7808 8174 7812 8230
rect 7748 8170 7812 8174
rect 7828 8230 7892 8234
rect 7828 8174 7832 8230
rect 7832 8174 7888 8230
rect 7888 8174 7892 8230
rect 7828 8170 7892 8174
rect 7908 8230 7972 8234
rect 7908 8174 7912 8230
rect 7912 8174 7968 8230
rect 7968 8174 7972 8230
rect 7908 8170 7972 8174
rect 7988 8230 8052 8234
rect 7988 8174 7992 8230
rect 7992 8174 8048 8230
rect 8048 8174 8052 8230
rect 7988 8170 8052 8174
rect 8068 8230 8132 8234
rect 8068 8174 8072 8230
rect 8072 8174 8128 8230
rect 8128 8174 8132 8230
rect 8068 8170 8132 8174
rect 8148 8230 8212 8234
rect 8148 8174 8152 8230
rect 8152 8174 8208 8230
rect 8208 8174 8212 8230
rect 8148 8170 8212 8174
rect 8228 8230 8292 8234
rect 8228 8174 8232 8230
rect 8232 8174 8288 8230
rect 8288 8174 8292 8230
rect 8228 8170 8292 8174
rect 8308 8230 8372 8234
rect 8308 8174 8312 8230
rect 8312 8174 8368 8230
rect 8368 8174 8372 8230
rect 8308 8170 8372 8174
rect 8388 8230 8452 8234
rect 8388 8174 8392 8230
rect 8392 8174 8448 8230
rect 8448 8174 8452 8230
rect 8388 8170 8452 8174
rect 8468 8230 8532 8234
rect 8468 8174 8472 8230
rect 8472 8174 8528 8230
rect 8528 8174 8532 8230
rect 8468 8170 8532 8174
rect 8548 8230 8612 8234
rect 8548 8174 8552 8230
rect 8552 8174 8608 8230
rect 8608 8174 8612 8230
rect 8548 8170 8612 8174
rect 8628 8230 8692 8234
rect 8628 8174 8632 8230
rect 8632 8174 8688 8230
rect 8688 8174 8692 8230
rect 8628 8170 8692 8174
rect 8708 8230 8772 8234
rect 8708 8174 8712 8230
rect 8712 8174 8768 8230
rect 8768 8174 8772 8230
rect 8708 8170 8772 8174
rect 8788 8230 8852 8234
rect 8788 8174 8792 8230
rect 8792 8174 8848 8230
rect 8848 8174 8852 8230
rect 8788 8170 8852 8174
rect 8868 8230 8932 8234
rect 8868 8174 8872 8230
rect 8872 8174 8928 8230
rect 8928 8174 8932 8230
rect 8868 8170 8932 8174
rect 8948 8230 9012 8234
rect 8948 8174 8952 8230
rect 8952 8174 9008 8230
rect 9008 8174 9012 8230
rect 8948 8170 9012 8174
rect 9028 8230 9092 8234
rect 9028 8174 9032 8230
rect 9032 8174 9088 8230
rect 9088 8174 9092 8230
rect 9028 8170 9092 8174
rect 9108 8230 9172 8234
rect 9108 8174 9112 8230
rect 9112 8174 9168 8230
rect 9168 8174 9172 8230
rect 9108 8170 9172 8174
rect 9188 8230 9252 8234
rect 9188 8174 9192 8230
rect 9192 8174 9248 8230
rect 9248 8174 9252 8230
rect 9188 8170 9252 8174
rect 9268 8230 9332 8234
rect 9268 8174 9272 8230
rect 9272 8174 9328 8230
rect 9328 8174 9332 8230
rect 9268 8170 9332 8174
rect 9348 8230 9412 8234
rect 9348 8174 9352 8230
rect 9352 8174 9408 8230
rect 9408 8174 9412 8230
rect 9348 8170 9412 8174
rect 9428 8230 9492 8234
rect 9428 8174 9432 8230
rect 9432 8174 9488 8230
rect 9488 8174 9492 8230
rect 9428 8170 9492 8174
rect 9508 8230 9572 8234
rect 9508 8174 9512 8230
rect 9512 8174 9568 8230
rect 9568 8174 9572 8230
rect 9508 8170 9572 8174
rect 9588 8230 9652 8234
rect 9588 8174 9592 8230
rect 9592 8174 9648 8230
rect 9648 8174 9652 8230
rect 9588 8170 9652 8174
rect 9668 8230 9732 8234
rect 9668 8174 9672 8230
rect 9672 8174 9728 8230
rect 9728 8174 9732 8230
rect 9668 8170 9732 8174
rect 9748 8230 9812 8234
rect 9748 8174 9752 8230
rect 9752 8174 9808 8230
rect 9808 8174 9812 8230
rect 9748 8170 9812 8174
rect 9828 8230 9892 8234
rect 9828 8174 9832 8230
rect 9832 8174 9888 8230
rect 9888 8174 9892 8230
rect 9828 8170 9892 8174
rect 9908 8230 9972 8234
rect 9908 8174 9912 8230
rect 9912 8174 9968 8230
rect 9968 8174 9972 8230
rect 9908 8170 9972 8174
rect 9988 8230 10052 8234
rect 9988 8174 9992 8230
rect 9992 8174 10048 8230
rect 10048 8174 10052 8230
rect 9988 8170 10052 8174
rect 10068 8230 10132 8234
rect 10068 8174 10072 8230
rect 10072 8174 10128 8230
rect 10128 8174 10132 8230
rect 10068 8170 10132 8174
rect 10148 8230 10212 8234
rect 10148 8174 10152 8230
rect 10152 8174 10208 8230
rect 10208 8174 10212 8230
rect 10148 8170 10212 8174
rect 10228 8230 10292 8234
rect 10228 8174 10232 8230
rect 10232 8174 10288 8230
rect 10288 8174 10292 8230
rect 10228 8170 10292 8174
rect 10308 8230 10372 8234
rect 10308 8174 10312 8230
rect 10312 8174 10368 8230
rect 10368 8174 10372 8230
rect 10308 8170 10372 8174
rect 10388 8230 10452 8234
rect 10388 8174 10392 8230
rect 10392 8174 10448 8230
rect 10448 8174 10452 8230
rect 10388 8170 10452 8174
rect 10468 8230 10532 8234
rect 10468 8174 10472 8230
rect 10472 8174 10528 8230
rect 10528 8174 10532 8230
rect 10468 8170 10532 8174
rect 10548 8230 10612 8234
rect 10548 8174 10552 8230
rect 10552 8174 10608 8230
rect 10608 8174 10612 8230
rect 10548 8170 10612 8174
rect 10628 8230 10692 8234
rect 10628 8174 10632 8230
rect 10632 8174 10688 8230
rect 10688 8174 10692 8230
rect 10628 8170 10692 8174
rect 10708 8230 10772 8234
rect 10708 8174 10712 8230
rect 10712 8174 10768 8230
rect 10768 8174 10772 8230
rect 10708 8170 10772 8174
rect 101 8010 7045 8114
rect 7345 7524 7409 7528
rect 7425 7524 7489 7528
rect 7505 7524 7569 7528
rect 7585 7524 7649 7528
rect 7665 7524 7729 7528
rect 7745 7524 7809 7528
rect 7825 7524 7889 7528
rect 7905 7524 7969 7528
rect 7985 7524 8049 7528
rect 8065 7524 8129 7528
rect 8145 7524 8209 7528
rect 8225 7524 8289 7528
rect 8305 7524 8369 7528
rect 7345 7468 7372 7524
rect 7372 7468 7396 7524
rect 7396 7468 7409 7524
rect 7425 7468 7452 7524
rect 7452 7468 7476 7524
rect 7476 7468 7489 7524
rect 7505 7468 7532 7524
rect 7532 7468 7556 7524
rect 7556 7468 7569 7524
rect 7585 7468 7612 7524
rect 7612 7468 7636 7524
rect 7636 7468 7649 7524
rect 7665 7468 7692 7524
rect 7692 7468 7716 7524
rect 7716 7468 7729 7524
rect 7745 7468 7772 7524
rect 7772 7468 7796 7524
rect 7796 7468 7809 7524
rect 7825 7468 7852 7524
rect 7852 7468 7876 7524
rect 7876 7468 7889 7524
rect 7905 7468 7932 7524
rect 7932 7468 7956 7524
rect 7956 7468 7969 7524
rect 7985 7468 8012 7524
rect 8012 7468 8036 7524
rect 8036 7468 8049 7524
rect 8065 7468 8092 7524
rect 8092 7468 8116 7524
rect 8116 7468 8129 7524
rect 8145 7468 8172 7524
rect 8172 7468 8196 7524
rect 8196 7468 8209 7524
rect 8225 7468 8252 7524
rect 8252 7468 8276 7524
rect 8276 7468 8289 7524
rect 8305 7468 8332 7524
rect 8332 7468 8369 7524
rect 7345 7464 7409 7468
rect 7425 7464 7489 7468
rect 7505 7464 7569 7468
rect 7585 7464 7649 7468
rect 7665 7464 7729 7468
rect 7745 7464 7809 7468
rect 7825 7464 7889 7468
rect 7905 7464 7969 7468
rect 7985 7464 8049 7468
rect 8065 7464 8129 7468
rect 8145 7464 8209 7468
rect 8225 7464 8289 7468
rect 8305 7464 8369 7468
rect 8385 7464 8449 7528
rect 8465 7464 8529 7528
rect 8545 7464 8609 7528
rect 8625 7524 8689 7528
rect 8705 7524 8769 7528
rect 8785 7524 8849 7528
rect 8865 7524 8929 7528
rect 8945 7524 9009 7528
rect 9025 7524 9089 7528
rect 9105 7524 9169 7528
rect 9185 7524 9249 7528
rect 9265 7524 9329 7528
rect 9345 7524 9409 7528
rect 9425 7524 9489 7528
rect 9505 7524 9569 7528
rect 9585 7524 9649 7528
rect 9665 7524 9729 7528
rect 9745 7524 9809 7528
rect 9825 7524 9889 7528
rect 9905 7524 9969 7528
rect 9985 7524 10049 7528
rect 10065 7524 10129 7528
rect 10145 7524 10209 7528
rect 10225 7524 10289 7528
rect 10305 7524 10369 7528
rect 10385 7524 10449 7528
rect 10465 7524 10529 7528
rect 10545 7524 10609 7528
rect 8625 7468 8645 7524
rect 8645 7468 8689 7524
rect 8705 7468 8725 7524
rect 8725 7468 8769 7524
rect 8785 7468 8805 7524
rect 8805 7468 8849 7524
rect 8865 7468 8885 7524
rect 8885 7468 8929 7524
rect 8945 7468 8965 7524
rect 8965 7468 9009 7524
rect 9025 7468 9045 7524
rect 9045 7468 9089 7524
rect 9105 7468 9125 7524
rect 9125 7468 9169 7524
rect 9185 7468 9205 7524
rect 9205 7468 9249 7524
rect 9265 7468 9285 7524
rect 9285 7468 9329 7524
rect 9345 7468 9365 7524
rect 9365 7468 9409 7524
rect 9425 7468 9445 7524
rect 9445 7468 9489 7524
rect 9505 7468 9525 7524
rect 9525 7468 9569 7524
rect 9585 7468 9605 7524
rect 9605 7468 9649 7524
rect 9665 7468 9685 7524
rect 9685 7468 9729 7524
rect 9745 7468 9765 7524
rect 9765 7468 9809 7524
rect 9825 7468 9845 7524
rect 9845 7468 9889 7524
rect 9905 7468 9925 7524
rect 9925 7468 9969 7524
rect 9985 7468 10005 7524
rect 10005 7468 10049 7524
rect 10065 7468 10085 7524
rect 10085 7468 10129 7524
rect 10145 7468 10165 7524
rect 10165 7468 10209 7524
rect 10225 7468 10245 7524
rect 10245 7468 10289 7524
rect 10305 7468 10325 7524
rect 10325 7468 10369 7524
rect 10385 7468 10405 7524
rect 10405 7468 10449 7524
rect 10465 7468 10485 7524
rect 10485 7468 10529 7524
rect 10545 7468 10565 7524
rect 10565 7468 10609 7524
rect 8625 7464 8689 7468
rect 8705 7464 8769 7468
rect 8785 7464 8849 7468
rect 8865 7464 8929 7468
rect 8945 7464 9009 7468
rect 9025 7464 9089 7468
rect 9105 7464 9169 7468
rect 9185 7464 9249 7468
rect 9265 7464 9329 7468
rect 9345 7464 9409 7468
rect 9425 7464 9489 7468
rect 9505 7464 9569 7468
rect 9585 7464 9649 7468
rect 9665 7464 9729 7468
rect 9745 7464 9809 7468
rect 9825 7464 9889 7468
rect 9905 7464 9969 7468
rect 9985 7464 10049 7468
rect 10065 7464 10129 7468
rect 10145 7464 10209 7468
rect 10225 7464 10289 7468
rect 10305 7464 10369 7468
rect 10385 7464 10449 7468
rect 10465 7464 10529 7468
rect 10545 7464 10609 7468
rect 4377 6833 5241 7269
rect 4377 6565 5241 6833
rect 6465 7017 6769 7021
rect 6465 6641 6469 7017
rect 6469 6641 6765 7017
rect 6765 6641 6769 7017
rect 6465 6637 6769 6641
<< metal4 >>
rect 38 8234 7126 8283
rect 38 8010 101 8234
rect 7045 8010 7126 8234
rect 38 7965 7126 8010
rect 7241 8234 11180 8291
rect 7241 8170 7348 8234
rect 7412 8170 7428 8234
rect 7492 8170 7508 8234
rect 7572 8170 7588 8234
rect 7652 8170 7668 8234
rect 7732 8170 7748 8234
rect 7812 8170 7828 8234
rect 7892 8170 7908 8234
rect 7972 8170 7988 8234
rect 8052 8170 8068 8234
rect 8132 8170 8148 8234
rect 8212 8170 8228 8234
rect 8292 8170 8308 8234
rect 8372 8170 8388 8234
rect 8452 8170 8468 8234
rect 8532 8170 8548 8234
rect 8612 8170 8628 8234
rect 8692 8170 8708 8234
rect 8772 8170 8788 8234
rect 8852 8170 8868 8234
rect 8932 8170 8948 8234
rect 9012 8170 9028 8234
rect 9092 8170 9108 8234
rect 9172 8170 9188 8234
rect 9252 8170 9268 8234
rect 9332 8170 9348 8234
rect 9412 8170 9428 8234
rect 9492 8170 9508 8234
rect 9572 8170 9588 8234
rect 9652 8170 9668 8234
rect 9732 8170 9748 8234
rect 9812 8170 9828 8234
rect 9892 8170 9908 8234
rect 9972 8170 9988 8234
rect 10052 8170 10068 8234
rect 10132 8170 10148 8234
rect 10212 8170 10228 8234
rect 10292 8170 10308 8234
rect 10372 8170 10388 8234
rect 10452 8170 10468 8234
rect 10532 8170 10548 8234
rect 10612 8170 10628 8234
rect 10692 8170 10708 8234
rect 10772 8170 11180 8234
rect 7241 7962 11180 8170
rect 38 7528 10667 7655
rect 38 7464 7345 7528
rect 7409 7464 7425 7528
rect 7489 7464 7505 7528
rect 7569 7464 7585 7528
rect 7649 7464 7665 7528
rect 7729 7464 7745 7528
rect 7809 7464 7825 7528
rect 7889 7464 7905 7528
rect 7969 7464 7985 7528
rect 8049 7464 8065 7528
rect 8129 7464 8145 7528
rect 8209 7464 8225 7528
rect 8289 7464 8305 7528
rect 8369 7464 8385 7528
rect 8449 7464 8465 7528
rect 8529 7464 8545 7528
rect 8609 7464 8625 7528
rect 8689 7464 8705 7528
rect 8769 7464 8785 7528
rect 8849 7464 8865 7528
rect 8929 7464 8945 7528
rect 9009 7464 9025 7528
rect 9089 7464 9105 7528
rect 9169 7464 9185 7528
rect 9249 7464 9265 7528
rect 9329 7464 9345 7528
rect 9409 7464 9425 7528
rect 9489 7464 9505 7528
rect 9569 7464 9585 7528
rect 9649 7464 9665 7528
rect 9729 7464 9745 7528
rect 9809 7464 9825 7528
rect 9889 7464 9905 7528
rect 9969 7464 9985 7528
rect 10049 7464 10065 7528
rect 10129 7464 10145 7528
rect 10209 7464 10225 7528
rect 10289 7464 10305 7528
rect 10369 7464 10385 7528
rect 10449 7464 10465 7528
rect 10529 7464 10545 7528
rect 10609 7464 10667 7528
rect 38 7269 10667 7464
rect 38 7255 4377 7269
rect 3817 7180 4377 7255
rect 5241 7255 10667 7269
rect 10843 7623 11178 7774
rect 10843 7387 10894 7623
rect 11130 7387 11178 7623
rect 10843 7303 11178 7387
rect 5241 7180 5299 7255
rect 3817 6624 4371 7180
rect 5247 6624 5299 7180
rect 10843 7074 10894 7303
rect 3817 6565 4377 6624
rect 5241 6565 5299 6624
rect 6386 7067 10894 7074
rect 11130 7067 11178 7303
rect 6386 7021 11178 7067
rect 6386 6637 6465 7021
rect 6769 6983 11178 7021
rect 6769 6747 10894 6983
rect 11130 6747 11178 6983
rect 6769 6637 11178 6747
rect 6386 6591 11178 6637
rect 3817 6522 5299 6565
rect 3817 51 4011 6522
rect 4101 51 4793 6251
<< via4 >>
rect 10894 7387 11130 7623
rect 4371 6624 4377 7180
rect 4377 6624 5241 7180
rect 5241 6624 5247 7180
rect 10894 7067 11130 7303
rect 10894 6747 11130 6983
<< metal5 >>
rect 10851 7623 11171 7779
rect 10851 7387 10894 7623
rect 11130 7387 11171 7623
rect 4313 7180 5299 7317
rect 4313 6624 4371 7180
rect 5247 6624 5299 7180
rect 4313 6494 5299 6624
rect 4507 6135 5299 6494
rect 10851 7303 11171 7387
rect 10851 7067 10894 7303
rect 11130 7067 11171 7303
rect 10851 6983 11171 7067
rect 10851 6747 10894 6983
rect 11130 6747 11171 6983
rect 10851 6242 11171 6747
use sky130_fd_pr__cap_mim_m3_1_WRT4AW  sky130_fd_pr__cap_mim_m3_1_WRT4AW_0
timestamp 1698351692
transform -1 0 7027 0 1 3151
box -3136 -3100 3136 3100
use sky130_fd_pr__cap_mim_m3_2_W5U4AW  sky130_fd_pr__cap_mim_m3_2_W5U4AW_0
timestamp 1698351692
transform 1 0 7970 0 1 3151
box -3179 -3101 3201 3101
use sky130_fd_pr__nfet_g5v0d10v5_PKVMTM  sky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0
timestamp 1698351692
transform 1 0 2660 0 1 6770
box -298 -448 298 448
use sky130_fd_pr__nfet_g5v0d10v5_TGFUGS  sky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0
timestamp 1698351692
transform 1 0 1515 0 1 6769
box -952 -448 952 448
use sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC  sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_0
timestamp 1698351692
transform -1 0 371 0 1 6769
box -298 -448 298 448
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0
timestamp 1698351692
transform 1 0 6644 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1
timestamp 1698351692
transform 1 0 3392 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2
timestamp 1698351692
transform 1 0 3878 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3
timestamp 1698351692
transform 1 0 408 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YEUEBV  sky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0
timestamp 1698351692
transform 1 0 5018 0 1 7841
box -992 -497 992 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPBG  sky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0
timestamp 1698351692
transform 1 0 2906 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPXE  sky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0
timestamp 1698351692
transform 1 0 6158 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ  sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0
timestamp 1698351692
transform 1 0 1657 0 1 7841
box -1101 -497 1101 497
use sky130_fd_pr__res_xhigh_po_0p69_S5N9F3  sky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0
timestamp 1698351692
transform 1 0 5446 0 1 3098
box -5436 -3088 5436 3088
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_0
timestamp 1698351692
transform 1 0 8523 0 1 6404
box -66 -43 1986 897
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_1
timestamp 1698351692
transform 1 0 7477 0 1 7438
box -66 -43 1986 897
use sky130_fd_sc_hvl__fill_4  sky130_fd_sc_hvl__fill_4_0
timestamp 1698351692
transform 1 0 10443 0 1 6404
box -66 -43 450 897
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_0
timestamp 1698351692
transform 1 0 9397 0 1 7438
box -66 -43 1506 897
use sky130_fd_sc_hvl__schmittbuf_1  sky130_fd_sc_hvl__schmittbuf_1_0
timestamp 1698351692
transform 1 0 7467 0 1 6404
box -66 -43 1122 897
<< labels >>
flabel metal4 s 38 7965 73 8283 0 FreeSans 400 0 0 0 vdd3v3
port 1 nsew
flabel metal4 s 10974 7962 11180 8291 0 FreeSans 400 0 0 0 vdd1v8
port 2 nsew
flabel metal4 s 38 7255 232 7655 0 FreeSans 400 0 0 0 vss
port 3 nsew
flabel metal3 s 10969 6765 11342 6834 0 FreeSans 400 0 0 0 porb_h
port 4 nsew
flabel metal3 s 11189 7491 11344 7551 0 FreeSans 400 0 0 0 por_l
port 5 nsew
flabel metal3 s 11188 7856 11343 7916 0 FreeSans 400 0 0 0 porb_l
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 11344 8338
<< end >>
