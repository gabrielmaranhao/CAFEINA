magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< nwell >>
rect 3549 -998 4227 -608
<< pmoshvt >>
rect 3663 -876 3863 -676
rect 3921 -876 4121 -676
<< pdiff >>
rect 3605 -691 3663 -676
rect 3605 -725 3617 -691
rect 3651 -725 3663 -691
rect 3605 -759 3663 -725
rect 3605 -793 3617 -759
rect 3651 -793 3663 -759
rect 3605 -827 3663 -793
rect 3605 -861 3617 -827
rect 3651 -861 3663 -827
rect 3605 -876 3663 -861
rect 3863 -876 3921 -676
rect 4121 -691 4179 -676
rect 4121 -725 4133 -691
rect 4167 -725 4179 -691
rect 4121 -759 4179 -725
rect 4121 -793 4133 -759
rect 4167 -793 4179 -759
rect 4121 -827 4179 -793
rect 4121 -861 4133 -827
rect 4167 -861 4179 -827
rect 4121 -876 4179 -861
<< pdiffc >>
rect 3617 -725 3651 -691
rect 3617 -793 3651 -759
rect 3617 -861 3651 -827
rect 4133 -725 4167 -691
rect 4133 -793 4167 -759
rect 4133 -861 4167 -827
<< poly >>
rect 3663 -676 3863 -650
rect 3921 -676 4121 -650
rect 3663 -923 3863 -876
rect 3663 -957 3712 -923
rect 3746 -957 3780 -923
rect 3814 -957 3863 -923
rect 3663 -973 3863 -957
rect 3921 -923 4121 -876
rect 3921 -957 3970 -923
rect 4004 -957 4038 -923
rect 4072 -957 4121 -923
rect 3921 -973 4121 -957
<< polycont >>
rect 3712 -957 3746 -923
rect 3780 -957 3814 -923
rect 3970 -957 4004 -923
rect 4038 -957 4072 -923
<< locali >>
rect 3617 -691 3651 -672
rect 3617 -759 3651 -757
rect 3617 -795 3651 -793
rect 3617 -880 3651 -861
rect 4133 -691 4167 -672
rect 4133 -759 4167 -757
rect 4133 -795 4167 -793
rect 4133 -880 4167 -861
rect 3663 -957 3710 -923
rect 3746 -957 3780 -923
rect 3816 -957 3863 -923
rect 3921 -957 3968 -923
rect 4004 -957 4038 -923
rect 4074 -957 4121 -923
<< viali >>
rect 3617 -725 3651 -723
rect 3617 -757 3651 -725
rect 3617 -827 3651 -795
rect 3617 -829 3651 -827
rect 4133 -725 4167 -723
rect 4133 -757 4167 -725
rect 4133 -827 4167 -795
rect 4133 -829 4167 -827
rect 3710 -957 3712 -923
rect 3712 -957 3744 -923
rect 3782 -957 3814 -923
rect 3814 -957 3816 -923
rect 3968 -957 3970 -923
rect 3970 -957 4002 -923
rect 4040 -957 4072 -923
rect 4072 -957 4074 -923
<< metal1 >>
rect 3611 -723 3657 -676
rect 3611 -757 3617 -723
rect 3651 -757 3657 -723
rect 3611 -795 3657 -757
rect 3611 -829 3617 -795
rect 3651 -829 3657 -795
rect 3611 -876 3657 -829
rect 4127 -723 4173 -676
rect 4127 -757 4133 -723
rect 4167 -757 4173 -723
rect 4127 -795 4173 -757
rect 4127 -829 4133 -795
rect 4167 -829 4173 -795
rect 4127 -876 4173 -829
rect 3667 -923 3859 -917
rect 3667 -957 3710 -923
rect 3744 -957 3782 -923
rect 3816 -957 3859 -923
rect 3667 -963 3859 -957
rect 3925 -923 4117 -917
rect 3925 -957 3968 -923
rect 4002 -957 4040 -923
rect 4074 -957 4117 -923
rect 3925 -963 4117 -957
<< end >>
