magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< pwell >>
rect -270 592 3355 1015
rect -270 398 -184 592
rect 3269 398 3355 592
rect -270 312 3355 398
rect -270 118 -184 312
rect 3269 118 3355 312
rect -270 -134 3355 118
rect -270 -555 -184 -134
rect 3269 -555 3355 -134
rect -270 -807 3355 -555
rect -270 -1000 -184 -807
rect 3269 -1000 3355 -807
rect -270 -1086 3355 -1000
rect -270 -1279 -184 -1086
rect 3269 -1279 3355 -1086
rect -270 -1531 3355 -1279
rect -270 -1952 -184 -1531
rect 3269 -1952 3355 -1531
rect -270 -2204 3355 -1952
rect -270 -2398 -184 -2204
rect 3269 -2398 3355 -2204
rect -270 -2484 3355 -2398
rect -270 -2678 -184 -2484
rect 3269 -2678 3355 -2484
rect -270 -3101 3355 -2678
<< nmos >>
rect -84 618 116 818
rect 421 618 621 818
rect 679 618 879 818
rect 1184 618 1384 818
rect 1442 618 1642 818
rect 1700 618 1900 818
rect 2205 618 2405 818
rect 2463 618 2663 818
rect 2969 618 3169 818
rect -84 -108 116 92
rect 421 -108 621 92
rect 679 -108 879 92
rect 1184 -108 1384 92
rect 1442 -108 1642 92
rect 1700 -108 1900 92
rect 2205 -108 2405 92
rect 2463 -108 2663 92
rect 2969 -108 3169 92
rect -84 -781 116 -581
rect 421 -781 621 -581
rect 679 -781 879 -581
rect 1184 -781 1384 -581
rect 1442 -781 1642 -581
rect 1700 -781 1900 -581
rect 2205 -781 2405 -581
rect 2463 -781 2663 -581
rect 2969 -781 3169 -581
rect -84 -1505 116 -1305
rect 421 -1505 621 -1305
rect 679 -1505 879 -1305
rect 1184 -1505 1384 -1305
rect 1442 -1505 1642 -1305
rect 1700 -1505 1900 -1305
rect 2205 -1505 2405 -1305
rect 2463 -1505 2663 -1305
rect 2969 -1505 3169 -1305
rect -84 -2178 116 -1978
rect 421 -2178 621 -1978
rect 679 -2178 879 -1978
rect 1184 -2178 1384 -1978
rect 1442 -2178 1642 -1978
rect 1700 -2178 1900 -1978
rect 2205 -2178 2405 -1978
rect 2463 -2178 2663 -1978
rect 2969 -2178 3169 -1978
rect -84 -2904 116 -2704
rect 421 -2904 621 -2704
rect 679 -2904 879 -2704
rect 1184 -2904 1384 -2704
rect 1442 -2904 1642 -2704
rect 1700 -2904 1900 -2704
rect 2205 -2904 2405 -2704
rect 2463 -2904 2663 -2704
rect 2969 -2904 3169 -2704
<< ndiff >>
rect -142 803 -84 818
rect -142 769 -130 803
rect -96 769 -84 803
rect -142 735 -84 769
rect -142 701 -130 735
rect -96 701 -84 735
rect -142 667 -84 701
rect -142 633 -130 667
rect -96 633 -84 667
rect -142 618 -84 633
rect 116 803 174 818
rect 116 769 128 803
rect 162 769 174 803
rect 116 735 174 769
rect 116 701 128 735
rect 162 701 174 735
rect 116 667 174 701
rect 116 633 128 667
rect 162 633 174 667
rect 116 618 174 633
rect 363 803 421 818
rect 363 769 375 803
rect 409 769 421 803
rect 363 735 421 769
rect 363 701 375 735
rect 409 701 421 735
rect 363 667 421 701
rect 363 633 375 667
rect 409 633 421 667
rect 363 618 421 633
rect 621 803 679 818
rect 621 769 633 803
rect 667 769 679 803
rect 621 735 679 769
rect 621 701 633 735
rect 667 701 679 735
rect 621 667 679 701
rect 621 633 633 667
rect 667 633 679 667
rect 621 618 679 633
rect 879 803 937 818
rect 879 769 891 803
rect 925 769 937 803
rect 879 735 937 769
rect 879 701 891 735
rect 925 701 937 735
rect 879 667 937 701
rect 879 633 891 667
rect 925 633 937 667
rect 879 618 937 633
rect 1126 803 1184 818
rect 1126 769 1138 803
rect 1172 769 1184 803
rect 1126 735 1184 769
rect 1126 701 1138 735
rect 1172 701 1184 735
rect 1126 667 1184 701
rect 1126 633 1138 667
rect 1172 633 1184 667
rect 1126 618 1184 633
rect 1384 803 1442 818
rect 1384 769 1396 803
rect 1430 769 1442 803
rect 1384 735 1442 769
rect 1384 701 1396 735
rect 1430 701 1442 735
rect 1384 667 1442 701
rect 1384 633 1396 667
rect 1430 633 1442 667
rect 1384 618 1442 633
rect 1642 803 1700 818
rect 1642 769 1654 803
rect 1688 769 1700 803
rect 1642 735 1700 769
rect 1642 701 1654 735
rect 1688 701 1700 735
rect 1642 667 1700 701
rect 1642 633 1654 667
rect 1688 633 1700 667
rect 1642 618 1700 633
rect 1900 803 1958 818
rect 1900 769 1912 803
rect 1946 769 1958 803
rect 1900 735 1958 769
rect 1900 701 1912 735
rect 1946 701 1958 735
rect 1900 667 1958 701
rect 1900 633 1912 667
rect 1946 633 1958 667
rect 1900 618 1958 633
rect 2147 803 2205 818
rect 2147 769 2159 803
rect 2193 769 2205 803
rect 2147 735 2205 769
rect 2147 701 2159 735
rect 2193 701 2205 735
rect 2147 667 2205 701
rect 2147 633 2159 667
rect 2193 633 2205 667
rect 2147 618 2205 633
rect 2405 803 2463 818
rect 2405 769 2417 803
rect 2451 769 2463 803
rect 2405 735 2463 769
rect 2405 701 2417 735
rect 2451 701 2463 735
rect 2405 667 2463 701
rect 2405 633 2417 667
rect 2451 633 2463 667
rect 2405 618 2463 633
rect 2663 803 2721 818
rect 2663 769 2675 803
rect 2709 769 2721 803
rect 2663 735 2721 769
rect 2663 701 2675 735
rect 2709 701 2721 735
rect 2663 667 2721 701
rect 2663 633 2675 667
rect 2709 633 2721 667
rect 2663 618 2721 633
rect 2911 803 2969 818
rect 2911 769 2923 803
rect 2957 769 2969 803
rect 2911 735 2969 769
rect 2911 701 2923 735
rect 2957 701 2969 735
rect 2911 667 2969 701
rect 2911 633 2923 667
rect 2957 633 2969 667
rect 2911 618 2969 633
rect 3169 803 3227 818
rect 3169 769 3181 803
rect 3215 769 3227 803
rect 3169 735 3227 769
rect 3169 701 3181 735
rect 3215 701 3227 735
rect 3169 667 3227 701
rect 3169 633 3181 667
rect 3215 633 3227 667
rect 3169 618 3227 633
rect -142 77 -84 92
rect -142 43 -130 77
rect -96 43 -84 77
rect -142 9 -84 43
rect -142 -25 -130 9
rect -96 -25 -84 9
rect -142 -59 -84 -25
rect -142 -93 -130 -59
rect -96 -93 -84 -59
rect -142 -108 -84 -93
rect 116 77 174 92
rect 116 43 128 77
rect 162 43 174 77
rect 116 9 174 43
rect 116 -25 128 9
rect 162 -25 174 9
rect 116 -59 174 -25
rect 116 -93 128 -59
rect 162 -93 174 -59
rect 116 -108 174 -93
rect 363 77 421 92
rect 363 43 375 77
rect 409 43 421 77
rect 363 9 421 43
rect 363 -25 375 9
rect 409 -25 421 9
rect 363 -59 421 -25
rect 363 -93 375 -59
rect 409 -93 421 -59
rect 363 -108 421 -93
rect 621 77 679 92
rect 621 43 633 77
rect 667 43 679 77
rect 621 9 679 43
rect 621 -25 633 9
rect 667 -25 679 9
rect 621 -59 679 -25
rect 621 -93 633 -59
rect 667 -93 679 -59
rect 621 -108 679 -93
rect 879 77 937 92
rect 879 43 891 77
rect 925 43 937 77
rect 879 9 937 43
rect 879 -25 891 9
rect 925 -25 937 9
rect 879 -59 937 -25
rect 879 -93 891 -59
rect 925 -93 937 -59
rect 879 -108 937 -93
rect 1126 77 1184 92
rect 1126 43 1138 77
rect 1172 43 1184 77
rect 1126 9 1184 43
rect 1126 -25 1138 9
rect 1172 -25 1184 9
rect 1126 -59 1184 -25
rect 1126 -93 1138 -59
rect 1172 -93 1184 -59
rect 1126 -108 1184 -93
rect 1384 77 1442 92
rect 1384 43 1396 77
rect 1430 43 1442 77
rect 1384 9 1442 43
rect 1384 -25 1396 9
rect 1430 -25 1442 9
rect 1384 -59 1442 -25
rect 1384 -93 1396 -59
rect 1430 -93 1442 -59
rect 1384 -108 1442 -93
rect 1642 77 1700 92
rect 1642 43 1654 77
rect 1688 43 1700 77
rect 1642 9 1700 43
rect 1642 -25 1654 9
rect 1688 -25 1700 9
rect 1642 -59 1700 -25
rect 1642 -93 1654 -59
rect 1688 -93 1700 -59
rect 1642 -108 1700 -93
rect 1900 77 1958 92
rect 1900 43 1912 77
rect 1946 43 1958 77
rect 1900 9 1958 43
rect 1900 -25 1912 9
rect 1946 -25 1958 9
rect 1900 -59 1958 -25
rect 1900 -93 1912 -59
rect 1946 -93 1958 -59
rect 1900 -108 1958 -93
rect 2147 77 2205 92
rect 2147 43 2159 77
rect 2193 43 2205 77
rect 2147 9 2205 43
rect 2147 -25 2159 9
rect 2193 -25 2205 9
rect 2147 -59 2205 -25
rect 2147 -93 2159 -59
rect 2193 -93 2205 -59
rect 2147 -108 2205 -93
rect 2405 77 2463 92
rect 2405 43 2417 77
rect 2451 43 2463 77
rect 2405 9 2463 43
rect 2405 -25 2417 9
rect 2451 -25 2463 9
rect 2405 -59 2463 -25
rect 2405 -93 2417 -59
rect 2451 -93 2463 -59
rect 2405 -108 2463 -93
rect 2663 77 2721 92
rect 2663 43 2675 77
rect 2709 43 2721 77
rect 2663 9 2721 43
rect 2663 -25 2675 9
rect 2709 -25 2721 9
rect 2663 -59 2721 -25
rect 2663 -93 2675 -59
rect 2709 -93 2721 -59
rect 2663 -108 2721 -93
rect 2911 77 2969 92
rect 2911 43 2923 77
rect 2957 43 2969 77
rect 2911 9 2969 43
rect 2911 -25 2923 9
rect 2957 -25 2969 9
rect 2911 -59 2969 -25
rect 2911 -93 2923 -59
rect 2957 -93 2969 -59
rect 2911 -108 2969 -93
rect 3169 77 3227 92
rect 3169 43 3181 77
rect 3215 43 3227 77
rect 3169 9 3227 43
rect 3169 -25 3181 9
rect 3215 -25 3227 9
rect 3169 -59 3227 -25
rect 3169 -93 3181 -59
rect 3215 -93 3227 -59
rect 3169 -108 3227 -93
rect -142 -596 -84 -581
rect -142 -630 -130 -596
rect -96 -630 -84 -596
rect -142 -664 -84 -630
rect -142 -698 -130 -664
rect -96 -698 -84 -664
rect -142 -732 -84 -698
rect -142 -766 -130 -732
rect -96 -766 -84 -732
rect -142 -781 -84 -766
rect 116 -596 174 -581
rect 116 -630 128 -596
rect 162 -630 174 -596
rect 116 -664 174 -630
rect 116 -698 128 -664
rect 162 -698 174 -664
rect 116 -732 174 -698
rect 116 -766 128 -732
rect 162 -766 174 -732
rect 116 -781 174 -766
rect 363 -596 421 -581
rect 363 -630 375 -596
rect 409 -630 421 -596
rect 363 -664 421 -630
rect 363 -698 375 -664
rect 409 -698 421 -664
rect 363 -732 421 -698
rect 363 -766 375 -732
rect 409 -766 421 -732
rect 363 -781 421 -766
rect 621 -596 679 -581
rect 621 -630 633 -596
rect 667 -630 679 -596
rect 621 -664 679 -630
rect 621 -698 633 -664
rect 667 -698 679 -664
rect 621 -732 679 -698
rect 621 -766 633 -732
rect 667 -766 679 -732
rect 621 -781 679 -766
rect 879 -596 937 -581
rect 879 -630 891 -596
rect 925 -630 937 -596
rect 879 -664 937 -630
rect 879 -698 891 -664
rect 925 -698 937 -664
rect 879 -732 937 -698
rect 879 -766 891 -732
rect 925 -766 937 -732
rect 879 -781 937 -766
rect 1126 -596 1184 -581
rect 1126 -630 1138 -596
rect 1172 -630 1184 -596
rect 1126 -664 1184 -630
rect 1126 -698 1138 -664
rect 1172 -698 1184 -664
rect 1126 -732 1184 -698
rect 1126 -766 1138 -732
rect 1172 -766 1184 -732
rect 1126 -781 1184 -766
rect 1384 -596 1442 -581
rect 1384 -630 1396 -596
rect 1430 -630 1442 -596
rect 1384 -664 1442 -630
rect 1384 -698 1396 -664
rect 1430 -698 1442 -664
rect 1384 -732 1442 -698
rect 1384 -766 1396 -732
rect 1430 -766 1442 -732
rect 1384 -781 1442 -766
rect 1642 -596 1700 -581
rect 1642 -630 1654 -596
rect 1688 -630 1700 -596
rect 1642 -664 1700 -630
rect 1642 -698 1654 -664
rect 1688 -698 1700 -664
rect 1642 -732 1700 -698
rect 1642 -766 1654 -732
rect 1688 -766 1700 -732
rect 1642 -781 1700 -766
rect 1900 -596 1958 -581
rect 1900 -630 1912 -596
rect 1946 -630 1958 -596
rect 1900 -664 1958 -630
rect 1900 -698 1912 -664
rect 1946 -698 1958 -664
rect 1900 -732 1958 -698
rect 1900 -766 1912 -732
rect 1946 -766 1958 -732
rect 1900 -781 1958 -766
rect 2147 -596 2205 -581
rect 2147 -630 2159 -596
rect 2193 -630 2205 -596
rect 2147 -664 2205 -630
rect 2147 -698 2159 -664
rect 2193 -698 2205 -664
rect 2147 -732 2205 -698
rect 2147 -766 2159 -732
rect 2193 -766 2205 -732
rect 2147 -781 2205 -766
rect 2405 -596 2463 -581
rect 2405 -630 2417 -596
rect 2451 -630 2463 -596
rect 2405 -664 2463 -630
rect 2405 -698 2417 -664
rect 2451 -698 2463 -664
rect 2405 -732 2463 -698
rect 2405 -766 2417 -732
rect 2451 -766 2463 -732
rect 2405 -781 2463 -766
rect 2663 -596 2721 -581
rect 2663 -630 2675 -596
rect 2709 -630 2721 -596
rect 2663 -664 2721 -630
rect 2663 -698 2675 -664
rect 2709 -698 2721 -664
rect 2663 -732 2721 -698
rect 2663 -766 2675 -732
rect 2709 -766 2721 -732
rect 2663 -781 2721 -766
rect 2911 -596 2969 -581
rect 2911 -630 2923 -596
rect 2957 -630 2969 -596
rect 2911 -664 2969 -630
rect 2911 -698 2923 -664
rect 2957 -698 2969 -664
rect 2911 -732 2969 -698
rect 2911 -766 2923 -732
rect 2957 -766 2969 -732
rect 2911 -781 2969 -766
rect 3169 -596 3227 -581
rect 3169 -630 3181 -596
rect 3215 -630 3227 -596
rect 3169 -664 3227 -630
rect 3169 -698 3181 -664
rect 3215 -698 3227 -664
rect 3169 -732 3227 -698
rect 3169 -766 3181 -732
rect 3215 -766 3227 -732
rect 3169 -781 3227 -766
rect -142 -1320 -84 -1305
rect -142 -1354 -130 -1320
rect -96 -1354 -84 -1320
rect -142 -1388 -84 -1354
rect -142 -1422 -130 -1388
rect -96 -1422 -84 -1388
rect -142 -1456 -84 -1422
rect -142 -1490 -130 -1456
rect -96 -1490 -84 -1456
rect -142 -1505 -84 -1490
rect 116 -1320 174 -1305
rect 116 -1354 128 -1320
rect 162 -1354 174 -1320
rect 116 -1388 174 -1354
rect 116 -1422 128 -1388
rect 162 -1422 174 -1388
rect 116 -1456 174 -1422
rect 116 -1490 128 -1456
rect 162 -1490 174 -1456
rect 116 -1505 174 -1490
rect 363 -1320 421 -1305
rect 363 -1354 375 -1320
rect 409 -1354 421 -1320
rect 363 -1388 421 -1354
rect 363 -1422 375 -1388
rect 409 -1422 421 -1388
rect 363 -1456 421 -1422
rect 363 -1490 375 -1456
rect 409 -1490 421 -1456
rect 363 -1505 421 -1490
rect 621 -1320 679 -1305
rect 621 -1354 633 -1320
rect 667 -1354 679 -1320
rect 621 -1388 679 -1354
rect 621 -1422 633 -1388
rect 667 -1422 679 -1388
rect 621 -1456 679 -1422
rect 621 -1490 633 -1456
rect 667 -1490 679 -1456
rect 621 -1505 679 -1490
rect 879 -1320 937 -1305
rect 879 -1354 891 -1320
rect 925 -1354 937 -1320
rect 879 -1388 937 -1354
rect 879 -1422 891 -1388
rect 925 -1422 937 -1388
rect 879 -1456 937 -1422
rect 879 -1490 891 -1456
rect 925 -1490 937 -1456
rect 879 -1505 937 -1490
rect 1126 -1320 1184 -1305
rect 1126 -1354 1138 -1320
rect 1172 -1354 1184 -1320
rect 1126 -1388 1184 -1354
rect 1126 -1422 1138 -1388
rect 1172 -1422 1184 -1388
rect 1126 -1456 1184 -1422
rect 1126 -1490 1138 -1456
rect 1172 -1490 1184 -1456
rect 1126 -1505 1184 -1490
rect 1384 -1320 1442 -1305
rect 1384 -1354 1396 -1320
rect 1430 -1354 1442 -1320
rect 1384 -1388 1442 -1354
rect 1384 -1422 1396 -1388
rect 1430 -1422 1442 -1388
rect 1384 -1456 1442 -1422
rect 1384 -1490 1396 -1456
rect 1430 -1490 1442 -1456
rect 1384 -1505 1442 -1490
rect 1642 -1320 1700 -1305
rect 1642 -1354 1654 -1320
rect 1688 -1354 1700 -1320
rect 1642 -1388 1700 -1354
rect 1642 -1422 1654 -1388
rect 1688 -1422 1700 -1388
rect 1642 -1456 1700 -1422
rect 1642 -1490 1654 -1456
rect 1688 -1490 1700 -1456
rect 1642 -1505 1700 -1490
rect 1900 -1320 1958 -1305
rect 1900 -1354 1912 -1320
rect 1946 -1354 1958 -1320
rect 1900 -1388 1958 -1354
rect 1900 -1422 1912 -1388
rect 1946 -1422 1958 -1388
rect 1900 -1456 1958 -1422
rect 1900 -1490 1912 -1456
rect 1946 -1490 1958 -1456
rect 1900 -1505 1958 -1490
rect 2147 -1320 2205 -1305
rect 2147 -1354 2159 -1320
rect 2193 -1354 2205 -1320
rect 2147 -1388 2205 -1354
rect 2147 -1422 2159 -1388
rect 2193 -1422 2205 -1388
rect 2147 -1456 2205 -1422
rect 2147 -1490 2159 -1456
rect 2193 -1490 2205 -1456
rect 2147 -1505 2205 -1490
rect 2405 -1320 2463 -1305
rect 2405 -1354 2417 -1320
rect 2451 -1354 2463 -1320
rect 2405 -1388 2463 -1354
rect 2405 -1422 2417 -1388
rect 2451 -1422 2463 -1388
rect 2405 -1456 2463 -1422
rect 2405 -1490 2417 -1456
rect 2451 -1490 2463 -1456
rect 2405 -1505 2463 -1490
rect 2663 -1320 2721 -1305
rect 2663 -1354 2675 -1320
rect 2709 -1354 2721 -1320
rect 2663 -1388 2721 -1354
rect 2663 -1422 2675 -1388
rect 2709 -1422 2721 -1388
rect 2663 -1456 2721 -1422
rect 2663 -1490 2675 -1456
rect 2709 -1490 2721 -1456
rect 2663 -1505 2721 -1490
rect 2911 -1320 2969 -1305
rect 2911 -1354 2923 -1320
rect 2957 -1354 2969 -1320
rect 2911 -1388 2969 -1354
rect 2911 -1422 2923 -1388
rect 2957 -1422 2969 -1388
rect 2911 -1456 2969 -1422
rect 2911 -1490 2923 -1456
rect 2957 -1490 2969 -1456
rect 2911 -1505 2969 -1490
rect 3169 -1320 3227 -1305
rect 3169 -1354 3181 -1320
rect 3215 -1354 3227 -1320
rect 3169 -1388 3227 -1354
rect 3169 -1422 3181 -1388
rect 3215 -1422 3227 -1388
rect 3169 -1456 3227 -1422
rect 3169 -1490 3181 -1456
rect 3215 -1490 3227 -1456
rect 3169 -1505 3227 -1490
rect -142 -1993 -84 -1978
rect -142 -2027 -130 -1993
rect -96 -2027 -84 -1993
rect -142 -2061 -84 -2027
rect -142 -2095 -130 -2061
rect -96 -2095 -84 -2061
rect -142 -2129 -84 -2095
rect -142 -2163 -130 -2129
rect -96 -2163 -84 -2129
rect -142 -2178 -84 -2163
rect 116 -1993 174 -1978
rect 116 -2027 128 -1993
rect 162 -2027 174 -1993
rect 116 -2061 174 -2027
rect 116 -2095 128 -2061
rect 162 -2095 174 -2061
rect 116 -2129 174 -2095
rect 116 -2163 128 -2129
rect 162 -2163 174 -2129
rect 116 -2178 174 -2163
rect 363 -1993 421 -1978
rect 363 -2027 375 -1993
rect 409 -2027 421 -1993
rect 363 -2061 421 -2027
rect 363 -2095 375 -2061
rect 409 -2095 421 -2061
rect 363 -2129 421 -2095
rect 363 -2163 375 -2129
rect 409 -2163 421 -2129
rect 363 -2178 421 -2163
rect 621 -1993 679 -1978
rect 621 -2027 633 -1993
rect 667 -2027 679 -1993
rect 621 -2061 679 -2027
rect 621 -2095 633 -2061
rect 667 -2095 679 -2061
rect 621 -2129 679 -2095
rect 621 -2163 633 -2129
rect 667 -2163 679 -2129
rect 621 -2178 679 -2163
rect 879 -1993 937 -1978
rect 879 -2027 891 -1993
rect 925 -2027 937 -1993
rect 879 -2061 937 -2027
rect 879 -2095 891 -2061
rect 925 -2095 937 -2061
rect 879 -2129 937 -2095
rect 879 -2163 891 -2129
rect 925 -2163 937 -2129
rect 879 -2178 937 -2163
rect 1126 -1993 1184 -1978
rect 1126 -2027 1138 -1993
rect 1172 -2027 1184 -1993
rect 1126 -2061 1184 -2027
rect 1126 -2095 1138 -2061
rect 1172 -2095 1184 -2061
rect 1126 -2129 1184 -2095
rect 1126 -2163 1138 -2129
rect 1172 -2163 1184 -2129
rect 1126 -2178 1184 -2163
rect 1384 -1993 1442 -1978
rect 1384 -2027 1396 -1993
rect 1430 -2027 1442 -1993
rect 1384 -2061 1442 -2027
rect 1384 -2095 1396 -2061
rect 1430 -2095 1442 -2061
rect 1384 -2129 1442 -2095
rect 1384 -2163 1396 -2129
rect 1430 -2163 1442 -2129
rect 1384 -2178 1442 -2163
rect 1642 -1993 1700 -1978
rect 1642 -2027 1654 -1993
rect 1688 -2027 1700 -1993
rect 1642 -2061 1700 -2027
rect 1642 -2095 1654 -2061
rect 1688 -2095 1700 -2061
rect 1642 -2129 1700 -2095
rect 1642 -2163 1654 -2129
rect 1688 -2163 1700 -2129
rect 1642 -2178 1700 -2163
rect 1900 -1993 1958 -1978
rect 1900 -2027 1912 -1993
rect 1946 -2027 1958 -1993
rect 1900 -2061 1958 -2027
rect 1900 -2095 1912 -2061
rect 1946 -2095 1958 -2061
rect 1900 -2129 1958 -2095
rect 1900 -2163 1912 -2129
rect 1946 -2163 1958 -2129
rect 1900 -2178 1958 -2163
rect 2147 -1993 2205 -1978
rect 2147 -2027 2159 -1993
rect 2193 -2027 2205 -1993
rect 2147 -2061 2205 -2027
rect 2147 -2095 2159 -2061
rect 2193 -2095 2205 -2061
rect 2147 -2129 2205 -2095
rect 2147 -2163 2159 -2129
rect 2193 -2163 2205 -2129
rect 2147 -2178 2205 -2163
rect 2405 -1993 2463 -1978
rect 2405 -2027 2417 -1993
rect 2451 -2027 2463 -1993
rect 2405 -2061 2463 -2027
rect 2405 -2095 2417 -2061
rect 2451 -2095 2463 -2061
rect 2405 -2129 2463 -2095
rect 2405 -2163 2417 -2129
rect 2451 -2163 2463 -2129
rect 2405 -2178 2463 -2163
rect 2663 -1993 2721 -1978
rect 2663 -2027 2675 -1993
rect 2709 -2027 2721 -1993
rect 2663 -2061 2721 -2027
rect 2663 -2095 2675 -2061
rect 2709 -2095 2721 -2061
rect 2663 -2129 2721 -2095
rect 2663 -2163 2675 -2129
rect 2709 -2163 2721 -2129
rect 2663 -2178 2721 -2163
rect 2911 -1993 2969 -1978
rect 2911 -2027 2923 -1993
rect 2957 -2027 2969 -1993
rect 2911 -2061 2969 -2027
rect 2911 -2095 2923 -2061
rect 2957 -2095 2969 -2061
rect 2911 -2129 2969 -2095
rect 2911 -2163 2923 -2129
rect 2957 -2163 2969 -2129
rect 2911 -2178 2969 -2163
rect 3169 -1993 3227 -1978
rect 3169 -2027 3181 -1993
rect 3215 -2027 3227 -1993
rect 3169 -2061 3227 -2027
rect 3169 -2095 3181 -2061
rect 3215 -2095 3227 -2061
rect 3169 -2129 3227 -2095
rect 3169 -2163 3181 -2129
rect 3215 -2163 3227 -2129
rect 3169 -2178 3227 -2163
rect -142 -2719 -84 -2704
rect -142 -2753 -130 -2719
rect -96 -2753 -84 -2719
rect -142 -2787 -84 -2753
rect -142 -2821 -130 -2787
rect -96 -2821 -84 -2787
rect -142 -2855 -84 -2821
rect -142 -2889 -130 -2855
rect -96 -2889 -84 -2855
rect -142 -2904 -84 -2889
rect 116 -2719 174 -2704
rect 116 -2753 128 -2719
rect 162 -2753 174 -2719
rect 116 -2787 174 -2753
rect 116 -2821 128 -2787
rect 162 -2821 174 -2787
rect 116 -2855 174 -2821
rect 116 -2889 128 -2855
rect 162 -2889 174 -2855
rect 116 -2904 174 -2889
rect 363 -2719 421 -2704
rect 363 -2753 375 -2719
rect 409 -2753 421 -2719
rect 363 -2787 421 -2753
rect 363 -2821 375 -2787
rect 409 -2821 421 -2787
rect 363 -2855 421 -2821
rect 363 -2889 375 -2855
rect 409 -2889 421 -2855
rect 363 -2904 421 -2889
rect 621 -2719 679 -2704
rect 621 -2753 633 -2719
rect 667 -2753 679 -2719
rect 621 -2787 679 -2753
rect 621 -2821 633 -2787
rect 667 -2821 679 -2787
rect 621 -2855 679 -2821
rect 621 -2889 633 -2855
rect 667 -2889 679 -2855
rect 621 -2904 679 -2889
rect 879 -2719 937 -2704
rect 879 -2753 891 -2719
rect 925 -2753 937 -2719
rect 879 -2787 937 -2753
rect 879 -2821 891 -2787
rect 925 -2821 937 -2787
rect 879 -2855 937 -2821
rect 879 -2889 891 -2855
rect 925 -2889 937 -2855
rect 879 -2904 937 -2889
rect 1126 -2719 1184 -2704
rect 1126 -2753 1138 -2719
rect 1172 -2753 1184 -2719
rect 1126 -2787 1184 -2753
rect 1126 -2821 1138 -2787
rect 1172 -2821 1184 -2787
rect 1126 -2855 1184 -2821
rect 1126 -2889 1138 -2855
rect 1172 -2889 1184 -2855
rect 1126 -2904 1184 -2889
rect 1384 -2719 1442 -2704
rect 1384 -2753 1396 -2719
rect 1430 -2753 1442 -2719
rect 1384 -2787 1442 -2753
rect 1384 -2821 1396 -2787
rect 1430 -2821 1442 -2787
rect 1384 -2855 1442 -2821
rect 1384 -2889 1396 -2855
rect 1430 -2889 1442 -2855
rect 1384 -2904 1442 -2889
rect 1642 -2719 1700 -2704
rect 1642 -2753 1654 -2719
rect 1688 -2753 1700 -2719
rect 1642 -2787 1700 -2753
rect 1642 -2821 1654 -2787
rect 1688 -2821 1700 -2787
rect 1642 -2855 1700 -2821
rect 1642 -2889 1654 -2855
rect 1688 -2889 1700 -2855
rect 1642 -2904 1700 -2889
rect 1900 -2719 1958 -2704
rect 1900 -2753 1912 -2719
rect 1946 -2753 1958 -2719
rect 1900 -2787 1958 -2753
rect 1900 -2821 1912 -2787
rect 1946 -2821 1958 -2787
rect 1900 -2855 1958 -2821
rect 1900 -2889 1912 -2855
rect 1946 -2889 1958 -2855
rect 1900 -2904 1958 -2889
rect 2147 -2719 2205 -2704
rect 2147 -2753 2159 -2719
rect 2193 -2753 2205 -2719
rect 2147 -2787 2205 -2753
rect 2147 -2821 2159 -2787
rect 2193 -2821 2205 -2787
rect 2147 -2855 2205 -2821
rect 2147 -2889 2159 -2855
rect 2193 -2889 2205 -2855
rect 2147 -2904 2205 -2889
rect 2405 -2719 2463 -2704
rect 2405 -2753 2417 -2719
rect 2451 -2753 2463 -2719
rect 2405 -2787 2463 -2753
rect 2405 -2821 2417 -2787
rect 2451 -2821 2463 -2787
rect 2405 -2855 2463 -2821
rect 2405 -2889 2417 -2855
rect 2451 -2889 2463 -2855
rect 2405 -2904 2463 -2889
rect 2663 -2719 2721 -2704
rect 2663 -2753 2675 -2719
rect 2709 -2753 2721 -2719
rect 2663 -2787 2721 -2753
rect 2663 -2821 2675 -2787
rect 2709 -2821 2721 -2787
rect 2663 -2855 2721 -2821
rect 2663 -2889 2675 -2855
rect 2709 -2889 2721 -2855
rect 2663 -2904 2721 -2889
rect 2911 -2719 2969 -2704
rect 2911 -2753 2923 -2719
rect 2957 -2753 2969 -2719
rect 2911 -2787 2969 -2753
rect 2911 -2821 2923 -2787
rect 2957 -2821 2969 -2787
rect 2911 -2855 2969 -2821
rect 2911 -2889 2923 -2855
rect 2957 -2889 2969 -2855
rect 2911 -2904 2969 -2889
rect 3169 -2719 3227 -2704
rect 3169 -2753 3181 -2719
rect 3215 -2753 3227 -2719
rect 3169 -2787 3227 -2753
rect 3169 -2821 3181 -2787
rect 3215 -2821 3227 -2787
rect 3169 -2855 3227 -2821
rect 3169 -2889 3181 -2855
rect 3215 -2889 3227 -2855
rect 3169 -2904 3227 -2889
<< ndiffc >>
rect -130 769 -96 803
rect -130 701 -96 735
rect -130 633 -96 667
rect 128 769 162 803
rect 128 701 162 735
rect 128 633 162 667
rect 375 769 409 803
rect 375 701 409 735
rect 375 633 409 667
rect 633 769 667 803
rect 633 701 667 735
rect 633 633 667 667
rect 891 769 925 803
rect 891 701 925 735
rect 891 633 925 667
rect 1138 769 1172 803
rect 1138 701 1172 735
rect 1138 633 1172 667
rect 1396 769 1430 803
rect 1396 701 1430 735
rect 1396 633 1430 667
rect 1654 769 1688 803
rect 1654 701 1688 735
rect 1654 633 1688 667
rect 1912 769 1946 803
rect 1912 701 1946 735
rect 1912 633 1946 667
rect 2159 769 2193 803
rect 2159 701 2193 735
rect 2159 633 2193 667
rect 2417 769 2451 803
rect 2417 701 2451 735
rect 2417 633 2451 667
rect 2675 769 2709 803
rect 2675 701 2709 735
rect 2675 633 2709 667
rect 2923 769 2957 803
rect 2923 701 2957 735
rect 2923 633 2957 667
rect 3181 769 3215 803
rect 3181 701 3215 735
rect 3181 633 3215 667
rect -130 43 -96 77
rect -130 -25 -96 9
rect -130 -93 -96 -59
rect 128 43 162 77
rect 128 -25 162 9
rect 128 -93 162 -59
rect 375 43 409 77
rect 375 -25 409 9
rect 375 -93 409 -59
rect 633 43 667 77
rect 633 -25 667 9
rect 633 -93 667 -59
rect 891 43 925 77
rect 891 -25 925 9
rect 891 -93 925 -59
rect 1138 43 1172 77
rect 1138 -25 1172 9
rect 1138 -93 1172 -59
rect 1396 43 1430 77
rect 1396 -25 1430 9
rect 1396 -93 1430 -59
rect 1654 43 1688 77
rect 1654 -25 1688 9
rect 1654 -93 1688 -59
rect 1912 43 1946 77
rect 1912 -25 1946 9
rect 1912 -93 1946 -59
rect 2159 43 2193 77
rect 2159 -25 2193 9
rect 2159 -93 2193 -59
rect 2417 43 2451 77
rect 2417 -25 2451 9
rect 2417 -93 2451 -59
rect 2675 43 2709 77
rect 2675 -25 2709 9
rect 2675 -93 2709 -59
rect 2923 43 2957 77
rect 2923 -25 2957 9
rect 2923 -93 2957 -59
rect 3181 43 3215 77
rect 3181 -25 3215 9
rect 3181 -93 3215 -59
rect -130 -630 -96 -596
rect -130 -698 -96 -664
rect -130 -766 -96 -732
rect 128 -630 162 -596
rect 128 -698 162 -664
rect 128 -766 162 -732
rect 375 -630 409 -596
rect 375 -698 409 -664
rect 375 -766 409 -732
rect 633 -630 667 -596
rect 633 -698 667 -664
rect 633 -766 667 -732
rect 891 -630 925 -596
rect 891 -698 925 -664
rect 891 -766 925 -732
rect 1138 -630 1172 -596
rect 1138 -698 1172 -664
rect 1138 -766 1172 -732
rect 1396 -630 1430 -596
rect 1396 -698 1430 -664
rect 1396 -766 1430 -732
rect 1654 -630 1688 -596
rect 1654 -698 1688 -664
rect 1654 -766 1688 -732
rect 1912 -630 1946 -596
rect 1912 -698 1946 -664
rect 1912 -766 1946 -732
rect 2159 -630 2193 -596
rect 2159 -698 2193 -664
rect 2159 -766 2193 -732
rect 2417 -630 2451 -596
rect 2417 -698 2451 -664
rect 2417 -766 2451 -732
rect 2675 -630 2709 -596
rect 2675 -698 2709 -664
rect 2675 -766 2709 -732
rect 2923 -630 2957 -596
rect 2923 -698 2957 -664
rect 2923 -766 2957 -732
rect 3181 -630 3215 -596
rect 3181 -698 3215 -664
rect 3181 -766 3215 -732
rect -130 -1354 -96 -1320
rect -130 -1422 -96 -1388
rect -130 -1490 -96 -1456
rect 128 -1354 162 -1320
rect 128 -1422 162 -1388
rect 128 -1490 162 -1456
rect 375 -1354 409 -1320
rect 375 -1422 409 -1388
rect 375 -1490 409 -1456
rect 633 -1354 667 -1320
rect 633 -1422 667 -1388
rect 633 -1490 667 -1456
rect 891 -1354 925 -1320
rect 891 -1422 925 -1388
rect 891 -1490 925 -1456
rect 1138 -1354 1172 -1320
rect 1138 -1422 1172 -1388
rect 1138 -1490 1172 -1456
rect 1396 -1354 1430 -1320
rect 1396 -1422 1430 -1388
rect 1396 -1490 1430 -1456
rect 1654 -1354 1688 -1320
rect 1654 -1422 1688 -1388
rect 1654 -1490 1688 -1456
rect 1912 -1354 1946 -1320
rect 1912 -1422 1946 -1388
rect 1912 -1490 1946 -1456
rect 2159 -1354 2193 -1320
rect 2159 -1422 2193 -1388
rect 2159 -1490 2193 -1456
rect 2417 -1354 2451 -1320
rect 2417 -1422 2451 -1388
rect 2417 -1490 2451 -1456
rect 2675 -1354 2709 -1320
rect 2675 -1422 2709 -1388
rect 2675 -1490 2709 -1456
rect 2923 -1354 2957 -1320
rect 2923 -1422 2957 -1388
rect 2923 -1490 2957 -1456
rect 3181 -1354 3215 -1320
rect 3181 -1422 3215 -1388
rect 3181 -1490 3215 -1456
rect -130 -2027 -96 -1993
rect -130 -2095 -96 -2061
rect -130 -2163 -96 -2129
rect 128 -2027 162 -1993
rect 128 -2095 162 -2061
rect 128 -2163 162 -2129
rect 375 -2027 409 -1993
rect 375 -2095 409 -2061
rect 375 -2163 409 -2129
rect 633 -2027 667 -1993
rect 633 -2095 667 -2061
rect 633 -2163 667 -2129
rect 891 -2027 925 -1993
rect 891 -2095 925 -2061
rect 891 -2163 925 -2129
rect 1138 -2027 1172 -1993
rect 1138 -2095 1172 -2061
rect 1138 -2163 1172 -2129
rect 1396 -2027 1430 -1993
rect 1396 -2095 1430 -2061
rect 1396 -2163 1430 -2129
rect 1654 -2027 1688 -1993
rect 1654 -2095 1688 -2061
rect 1654 -2163 1688 -2129
rect 1912 -2027 1946 -1993
rect 1912 -2095 1946 -2061
rect 1912 -2163 1946 -2129
rect 2159 -2027 2193 -1993
rect 2159 -2095 2193 -2061
rect 2159 -2163 2193 -2129
rect 2417 -2027 2451 -1993
rect 2417 -2095 2451 -2061
rect 2417 -2163 2451 -2129
rect 2675 -2027 2709 -1993
rect 2675 -2095 2709 -2061
rect 2675 -2163 2709 -2129
rect 2923 -2027 2957 -1993
rect 2923 -2095 2957 -2061
rect 2923 -2163 2957 -2129
rect 3181 -2027 3215 -1993
rect 3181 -2095 3215 -2061
rect 3181 -2163 3215 -2129
rect -130 -2753 -96 -2719
rect -130 -2821 -96 -2787
rect -130 -2889 -96 -2855
rect 128 -2753 162 -2719
rect 128 -2821 162 -2787
rect 128 -2889 162 -2855
rect 375 -2753 409 -2719
rect 375 -2821 409 -2787
rect 375 -2889 409 -2855
rect 633 -2753 667 -2719
rect 633 -2821 667 -2787
rect 633 -2889 667 -2855
rect 891 -2753 925 -2719
rect 891 -2821 925 -2787
rect 891 -2889 925 -2855
rect 1138 -2753 1172 -2719
rect 1138 -2821 1172 -2787
rect 1138 -2889 1172 -2855
rect 1396 -2753 1430 -2719
rect 1396 -2821 1430 -2787
rect 1396 -2889 1430 -2855
rect 1654 -2753 1688 -2719
rect 1654 -2821 1688 -2787
rect 1654 -2889 1688 -2855
rect 1912 -2753 1946 -2719
rect 1912 -2821 1946 -2787
rect 1912 -2889 1946 -2855
rect 2159 -2753 2193 -2719
rect 2159 -2821 2193 -2787
rect 2159 -2889 2193 -2855
rect 2417 -2753 2451 -2719
rect 2417 -2821 2451 -2787
rect 2417 -2889 2451 -2855
rect 2675 -2753 2709 -2719
rect 2675 -2821 2709 -2787
rect 2675 -2889 2709 -2855
rect 2923 -2753 2957 -2719
rect 2923 -2821 2957 -2787
rect 2923 -2889 2957 -2855
rect 3181 -2753 3215 -2719
rect 3181 -2821 3215 -2787
rect 3181 -2889 3215 -2855
<< psubdiff >>
rect -244 955 -59 989
rect -25 955 9 989
rect 43 955 77 989
rect 111 955 145 989
rect 179 955 213 989
rect 247 955 281 989
rect 315 955 349 989
rect 383 955 417 989
rect 451 955 485 989
rect 519 955 553 989
rect 587 955 621 989
rect 655 955 689 989
rect 723 955 757 989
rect 791 955 825 989
rect 859 955 893 989
rect 927 955 961 989
rect 995 955 1029 989
rect 1063 955 1097 989
rect 1131 955 1165 989
rect 1199 955 1233 989
rect 1267 955 1301 989
rect 1335 955 1369 989
rect 1403 955 1437 989
rect 1471 955 1505 989
rect 1539 955 1573 989
rect 1607 955 1641 989
rect 1675 955 1709 989
rect 1743 955 1777 989
rect 1811 955 1845 989
rect 1879 955 1913 989
rect 1947 955 1981 989
rect 2015 955 2049 989
rect 2083 955 2117 989
rect 2151 955 2185 989
rect 2219 955 2253 989
rect 2287 955 2321 989
rect 2355 955 2389 989
rect 2423 955 2457 989
rect 2491 955 2525 989
rect 2559 955 2593 989
rect 2627 955 2661 989
rect 2695 955 2729 989
rect 2763 955 2797 989
rect 2831 955 2865 989
rect 2899 955 2933 989
rect 2967 955 3001 989
rect 3035 955 3069 989
rect 3103 955 3137 989
rect 3171 955 3329 989
rect -244 848 -210 955
rect 3295 848 3329 955
rect -244 780 -210 814
rect -244 712 -210 746
rect -244 644 -210 678
rect 3295 780 3329 814
rect 3295 712 3329 746
rect 3295 644 3329 678
rect -244 576 -210 610
rect -244 508 -210 542
rect -244 440 -210 474
rect -244 372 -210 406
rect 3295 576 3329 610
rect 3295 508 3329 542
rect 3295 440 3329 474
rect 3295 372 3329 406
rect -210 338 -59 372
rect -25 338 9 372
rect 43 338 77 372
rect 111 338 145 372
rect 179 338 213 372
rect 247 338 281 372
rect 315 338 349 372
rect 383 338 417 372
rect 451 338 485 372
rect 519 338 553 372
rect 587 338 621 372
rect 655 338 689 372
rect 723 338 757 372
rect 791 338 825 372
rect 859 338 893 372
rect 927 338 961 372
rect 995 338 1029 372
rect 1063 338 1097 372
rect 1131 338 1165 372
rect 1199 338 1233 372
rect 1267 338 1301 372
rect 1335 338 1369 372
rect 1403 338 1437 372
rect 1471 338 1505 372
rect 1539 338 1573 372
rect 1607 338 1641 372
rect 1675 338 1709 372
rect 1743 338 1777 372
rect 1811 338 1845 372
rect 1879 338 1913 372
rect 1947 338 1981 372
rect 2015 338 2049 372
rect 2083 338 2117 372
rect 2151 338 2185 372
rect 2219 338 2253 372
rect 2287 338 2321 372
rect 2355 338 2389 372
rect 2423 338 2457 372
rect 2491 338 2525 372
rect 2559 338 2593 372
rect 2627 338 2661 372
rect 2695 338 2729 372
rect 2763 338 2797 372
rect 2831 338 2865 372
rect 2899 338 2933 372
rect 2967 338 3001 372
rect 3035 338 3069 372
rect 3103 338 3137 372
rect 3171 338 3295 372
rect -244 304 -210 338
rect -244 236 -210 270
rect -244 168 -210 202
rect -244 100 -210 134
rect 3295 304 3329 338
rect 3295 236 3329 270
rect 3295 168 3329 202
rect 3295 100 3329 134
rect -244 32 -210 66
rect -244 -36 -210 -2
rect -244 -104 -210 -70
rect 3295 32 3329 66
rect 3295 -36 3329 -2
rect 3295 -104 3329 -70
rect -244 -172 -210 -138
rect 3295 -172 3329 -138
rect -244 -240 -210 -206
rect -244 -308 -210 -274
rect -244 -376 -210 -342
rect -244 -444 -210 -410
rect -244 -512 -210 -478
rect 3295 -240 3329 -206
rect 3295 -308 3329 -274
rect 3295 -376 3329 -342
rect 3295 -444 3329 -410
rect -244 -580 -210 -546
rect 3295 -512 3329 -478
rect 3295 -580 3329 -546
rect -244 -648 -210 -614
rect -244 -716 -210 -682
rect -244 -784 -210 -750
rect 3295 -648 3329 -614
rect 3295 -716 3329 -682
rect 3295 -784 3329 -750
rect -244 -852 -210 -818
rect -244 -1026 -210 -886
rect 3295 -852 3329 -818
rect 3295 -1026 3329 -886
rect -244 -1060 -59 -1026
rect -25 -1060 9 -1026
rect 43 -1060 77 -1026
rect 111 -1060 145 -1026
rect 179 -1060 213 -1026
rect 247 -1060 281 -1026
rect 315 -1060 349 -1026
rect 383 -1060 417 -1026
rect 451 -1060 485 -1026
rect 519 -1060 553 -1026
rect 587 -1060 621 -1026
rect 655 -1060 689 -1026
rect 723 -1060 757 -1026
rect 791 -1060 825 -1026
rect 859 -1060 893 -1026
rect 927 -1060 961 -1026
rect 995 -1060 1029 -1026
rect 1063 -1060 1097 -1026
rect 1131 -1060 1165 -1026
rect 1199 -1060 1233 -1026
rect 1267 -1060 1301 -1026
rect 1335 -1060 1369 -1026
rect 1403 -1060 1437 -1026
rect 1471 -1060 1505 -1026
rect 1539 -1060 1573 -1026
rect 1607 -1060 1641 -1026
rect 1675 -1060 1709 -1026
rect 1743 -1060 1777 -1026
rect 1811 -1060 1845 -1026
rect 1879 -1060 1913 -1026
rect 1947 -1060 1981 -1026
rect 2015 -1060 2049 -1026
rect 2083 -1060 2117 -1026
rect 2151 -1060 2185 -1026
rect 2219 -1060 2253 -1026
rect 2287 -1060 2321 -1026
rect 2355 -1060 2389 -1026
rect 2423 -1060 2457 -1026
rect 2491 -1060 2525 -1026
rect 2559 -1060 2593 -1026
rect 2627 -1060 2661 -1026
rect 2695 -1060 2729 -1026
rect 2763 -1060 2797 -1026
rect 2831 -1060 2865 -1026
rect 2899 -1060 2933 -1026
rect 2967 -1060 3001 -1026
rect 3035 -1060 3069 -1026
rect 3103 -1060 3137 -1026
rect 3171 -1060 3329 -1026
rect -244 -1200 -210 -1060
rect -244 -1268 -210 -1234
rect 3295 -1200 3329 -1060
rect 3295 -1268 3329 -1234
rect -244 -1336 -210 -1302
rect -244 -1404 -210 -1370
rect -244 -1472 -210 -1438
rect 3295 -1336 3329 -1302
rect 3295 -1404 3329 -1370
rect 3295 -1472 3329 -1438
rect -244 -1540 -210 -1506
rect -244 -1608 -210 -1574
rect 3295 -1540 3329 -1506
rect -244 -1676 -210 -1642
rect -244 -1744 -210 -1710
rect -244 -1812 -210 -1778
rect -244 -1880 -210 -1846
rect 3295 -1608 3329 -1574
rect 3295 -1676 3329 -1642
rect 3295 -1744 3329 -1710
rect 3295 -1812 3329 -1778
rect 3295 -1880 3329 -1846
rect -244 -1948 -210 -1914
rect 3295 -1948 3329 -1914
rect -244 -2016 -210 -1982
rect -244 -2084 -210 -2050
rect -244 -2152 -210 -2118
rect 3295 -2016 3329 -1982
rect 3295 -2084 3329 -2050
rect 3295 -2152 3329 -2118
rect -244 -2220 -210 -2186
rect -244 -2288 -210 -2254
rect -244 -2356 -210 -2322
rect -244 -2424 -210 -2390
rect 3295 -2220 3329 -2186
rect 3295 -2288 3329 -2254
rect 3295 -2356 3329 -2322
rect 3295 -2424 3329 -2390
rect -210 -2458 -59 -2424
rect -25 -2458 9 -2424
rect 43 -2458 77 -2424
rect 111 -2458 145 -2424
rect 179 -2458 213 -2424
rect 247 -2458 281 -2424
rect 315 -2458 349 -2424
rect 383 -2458 417 -2424
rect 451 -2458 485 -2424
rect 519 -2458 553 -2424
rect 587 -2458 621 -2424
rect 655 -2458 689 -2424
rect 723 -2458 757 -2424
rect 791 -2458 825 -2424
rect 859 -2458 893 -2424
rect 927 -2458 961 -2424
rect 995 -2458 1029 -2424
rect 1063 -2458 1097 -2424
rect 1131 -2458 1165 -2424
rect 1199 -2458 1233 -2424
rect 1267 -2458 1301 -2424
rect 1335 -2458 1369 -2424
rect 1403 -2458 1437 -2424
rect 1471 -2458 1505 -2424
rect 1539 -2458 1573 -2424
rect 1607 -2458 1641 -2424
rect 1675 -2458 1709 -2424
rect 1743 -2458 1777 -2424
rect 1811 -2458 1845 -2424
rect 1879 -2458 1913 -2424
rect 1947 -2458 1981 -2424
rect 2015 -2458 2049 -2424
rect 2083 -2458 2117 -2424
rect 2151 -2458 2185 -2424
rect 2219 -2458 2253 -2424
rect 2287 -2458 2321 -2424
rect 2355 -2458 2389 -2424
rect 2423 -2458 2457 -2424
rect 2491 -2458 2525 -2424
rect 2559 -2458 2593 -2424
rect 2627 -2458 2661 -2424
rect 2695 -2458 2729 -2424
rect 2763 -2458 2797 -2424
rect 2831 -2458 2865 -2424
rect 2899 -2458 2933 -2424
rect 2967 -2458 3001 -2424
rect 3035 -2458 3069 -2424
rect 3103 -2458 3137 -2424
rect 3171 -2458 3295 -2424
rect -244 -2492 -210 -2458
rect -244 -2560 -210 -2526
rect -244 -2628 -210 -2594
rect -244 -2696 -210 -2662
rect 3295 -2492 3329 -2458
rect 3295 -2560 3329 -2526
rect 3295 -2628 3329 -2594
rect 3295 -2696 3329 -2662
rect -244 -2764 -210 -2730
rect -244 -2832 -210 -2798
rect -244 -2900 -210 -2866
rect 3295 -2764 3329 -2730
rect 3295 -2832 3329 -2798
rect 3295 -2900 3329 -2866
rect -244 -3041 -210 -2934
rect 3295 -3041 3329 -2934
rect -244 -3075 -59 -3041
rect -25 -3075 9 -3041
rect 43 -3075 77 -3041
rect 111 -3075 145 -3041
rect 179 -3075 213 -3041
rect 247 -3075 281 -3041
rect 315 -3075 349 -3041
rect 383 -3075 417 -3041
rect 451 -3075 485 -3041
rect 519 -3075 553 -3041
rect 587 -3075 621 -3041
rect 655 -3075 689 -3041
rect 723 -3075 757 -3041
rect 791 -3075 825 -3041
rect 859 -3075 893 -3041
rect 927 -3075 961 -3041
rect 995 -3075 1029 -3041
rect 1063 -3075 1097 -3041
rect 1131 -3075 1165 -3041
rect 1199 -3075 1233 -3041
rect 1267 -3075 1301 -3041
rect 1335 -3075 1369 -3041
rect 1403 -3075 1437 -3041
rect 1471 -3075 1505 -3041
rect 1539 -3075 1573 -3041
rect 1607 -3075 1641 -3041
rect 1675 -3075 1709 -3041
rect 1743 -3075 1777 -3041
rect 1811 -3075 1845 -3041
rect 1879 -3075 1913 -3041
rect 1947 -3075 1981 -3041
rect 2015 -3075 2049 -3041
rect 2083 -3075 2117 -3041
rect 2151 -3075 2185 -3041
rect 2219 -3075 2253 -3041
rect 2287 -3075 2321 -3041
rect 2355 -3075 2389 -3041
rect 2423 -3075 2457 -3041
rect 2491 -3075 2525 -3041
rect 2559 -3075 2593 -3041
rect 2627 -3075 2661 -3041
rect 2695 -3075 2729 -3041
rect 2763 -3075 2797 -3041
rect 2831 -3075 2865 -3041
rect 2899 -3075 2933 -3041
rect 2967 -3075 3001 -3041
rect 3035 -3075 3069 -3041
rect 3103 -3075 3137 -3041
rect 3171 -3075 3329 -3041
<< psubdiffcont >>
rect -59 955 -25 989
rect 9 955 43 989
rect 77 955 111 989
rect 145 955 179 989
rect 213 955 247 989
rect 281 955 315 989
rect 349 955 383 989
rect 417 955 451 989
rect 485 955 519 989
rect 553 955 587 989
rect 621 955 655 989
rect 689 955 723 989
rect 757 955 791 989
rect 825 955 859 989
rect 893 955 927 989
rect 961 955 995 989
rect 1029 955 1063 989
rect 1097 955 1131 989
rect 1165 955 1199 989
rect 1233 955 1267 989
rect 1301 955 1335 989
rect 1369 955 1403 989
rect 1437 955 1471 989
rect 1505 955 1539 989
rect 1573 955 1607 989
rect 1641 955 1675 989
rect 1709 955 1743 989
rect 1777 955 1811 989
rect 1845 955 1879 989
rect 1913 955 1947 989
rect 1981 955 2015 989
rect 2049 955 2083 989
rect 2117 955 2151 989
rect 2185 955 2219 989
rect 2253 955 2287 989
rect 2321 955 2355 989
rect 2389 955 2423 989
rect 2457 955 2491 989
rect 2525 955 2559 989
rect 2593 955 2627 989
rect 2661 955 2695 989
rect 2729 955 2763 989
rect 2797 955 2831 989
rect 2865 955 2899 989
rect 2933 955 2967 989
rect 3001 955 3035 989
rect 3069 955 3103 989
rect 3137 955 3171 989
rect -244 814 -210 848
rect -244 746 -210 780
rect -244 678 -210 712
rect -244 610 -210 644
rect 3295 814 3329 848
rect 3295 746 3329 780
rect 3295 678 3329 712
rect 3295 610 3329 644
rect -244 542 -210 576
rect -244 474 -210 508
rect -244 406 -210 440
rect 3295 542 3329 576
rect 3295 474 3329 508
rect 3295 406 3329 440
rect -244 338 -210 372
rect -59 338 -25 372
rect 9 338 43 372
rect 77 338 111 372
rect 145 338 179 372
rect 213 338 247 372
rect 281 338 315 372
rect 349 338 383 372
rect 417 338 451 372
rect 485 338 519 372
rect 553 338 587 372
rect 621 338 655 372
rect 689 338 723 372
rect 757 338 791 372
rect 825 338 859 372
rect 893 338 927 372
rect 961 338 995 372
rect 1029 338 1063 372
rect 1097 338 1131 372
rect 1165 338 1199 372
rect 1233 338 1267 372
rect 1301 338 1335 372
rect 1369 338 1403 372
rect 1437 338 1471 372
rect 1505 338 1539 372
rect 1573 338 1607 372
rect 1641 338 1675 372
rect 1709 338 1743 372
rect 1777 338 1811 372
rect 1845 338 1879 372
rect 1913 338 1947 372
rect 1981 338 2015 372
rect 2049 338 2083 372
rect 2117 338 2151 372
rect 2185 338 2219 372
rect 2253 338 2287 372
rect 2321 338 2355 372
rect 2389 338 2423 372
rect 2457 338 2491 372
rect 2525 338 2559 372
rect 2593 338 2627 372
rect 2661 338 2695 372
rect 2729 338 2763 372
rect 2797 338 2831 372
rect 2865 338 2899 372
rect 2933 338 2967 372
rect 3001 338 3035 372
rect 3069 338 3103 372
rect 3137 338 3171 372
rect 3295 338 3329 372
rect -244 270 -210 304
rect -244 202 -210 236
rect -244 134 -210 168
rect 3295 270 3329 304
rect 3295 202 3329 236
rect 3295 134 3329 168
rect -244 66 -210 100
rect -244 -2 -210 32
rect -244 -70 -210 -36
rect -244 -138 -210 -104
rect 3295 66 3329 100
rect 3295 -2 3329 32
rect 3295 -70 3329 -36
rect -244 -206 -210 -172
rect 3295 -138 3329 -104
rect -244 -274 -210 -240
rect -244 -342 -210 -308
rect -244 -410 -210 -376
rect -244 -478 -210 -444
rect 3295 -206 3329 -172
rect 3295 -274 3329 -240
rect 3295 -342 3329 -308
rect 3295 -410 3329 -376
rect 3295 -478 3329 -444
rect -244 -546 -210 -512
rect -244 -614 -210 -580
rect 3295 -546 3329 -512
rect -244 -682 -210 -648
rect -244 -750 -210 -716
rect 3295 -614 3329 -580
rect 3295 -682 3329 -648
rect 3295 -750 3329 -716
rect -244 -818 -210 -784
rect -244 -886 -210 -852
rect 3295 -818 3329 -784
rect 3295 -886 3329 -852
rect -59 -1060 -25 -1026
rect 9 -1060 43 -1026
rect 77 -1060 111 -1026
rect 145 -1060 179 -1026
rect 213 -1060 247 -1026
rect 281 -1060 315 -1026
rect 349 -1060 383 -1026
rect 417 -1060 451 -1026
rect 485 -1060 519 -1026
rect 553 -1060 587 -1026
rect 621 -1060 655 -1026
rect 689 -1060 723 -1026
rect 757 -1060 791 -1026
rect 825 -1060 859 -1026
rect 893 -1060 927 -1026
rect 961 -1060 995 -1026
rect 1029 -1060 1063 -1026
rect 1097 -1060 1131 -1026
rect 1165 -1060 1199 -1026
rect 1233 -1060 1267 -1026
rect 1301 -1060 1335 -1026
rect 1369 -1060 1403 -1026
rect 1437 -1060 1471 -1026
rect 1505 -1060 1539 -1026
rect 1573 -1060 1607 -1026
rect 1641 -1060 1675 -1026
rect 1709 -1060 1743 -1026
rect 1777 -1060 1811 -1026
rect 1845 -1060 1879 -1026
rect 1913 -1060 1947 -1026
rect 1981 -1060 2015 -1026
rect 2049 -1060 2083 -1026
rect 2117 -1060 2151 -1026
rect 2185 -1060 2219 -1026
rect 2253 -1060 2287 -1026
rect 2321 -1060 2355 -1026
rect 2389 -1060 2423 -1026
rect 2457 -1060 2491 -1026
rect 2525 -1060 2559 -1026
rect 2593 -1060 2627 -1026
rect 2661 -1060 2695 -1026
rect 2729 -1060 2763 -1026
rect 2797 -1060 2831 -1026
rect 2865 -1060 2899 -1026
rect 2933 -1060 2967 -1026
rect 3001 -1060 3035 -1026
rect 3069 -1060 3103 -1026
rect 3137 -1060 3171 -1026
rect -244 -1234 -210 -1200
rect -244 -1302 -210 -1268
rect 3295 -1234 3329 -1200
rect 3295 -1302 3329 -1268
rect -244 -1370 -210 -1336
rect -244 -1438 -210 -1404
rect -244 -1506 -210 -1472
rect 3295 -1370 3329 -1336
rect 3295 -1438 3329 -1404
rect -244 -1574 -210 -1540
rect 3295 -1506 3329 -1472
rect 3295 -1574 3329 -1540
rect -244 -1642 -210 -1608
rect -244 -1710 -210 -1676
rect -244 -1778 -210 -1744
rect -244 -1846 -210 -1812
rect -244 -1914 -210 -1880
rect 3295 -1642 3329 -1608
rect 3295 -1710 3329 -1676
rect 3295 -1778 3329 -1744
rect 3295 -1846 3329 -1812
rect -244 -1982 -210 -1948
rect 3295 -1914 3329 -1880
rect -244 -2050 -210 -2016
rect -244 -2118 -210 -2084
rect -244 -2186 -210 -2152
rect 3295 -1982 3329 -1948
rect 3295 -2050 3329 -2016
rect 3295 -2118 3329 -2084
rect 3295 -2186 3329 -2152
rect -244 -2254 -210 -2220
rect -244 -2322 -210 -2288
rect -244 -2390 -210 -2356
rect 3295 -2254 3329 -2220
rect 3295 -2322 3329 -2288
rect 3295 -2390 3329 -2356
rect -244 -2458 -210 -2424
rect -59 -2458 -25 -2424
rect 9 -2458 43 -2424
rect 77 -2458 111 -2424
rect 145 -2458 179 -2424
rect 213 -2458 247 -2424
rect 281 -2458 315 -2424
rect 349 -2458 383 -2424
rect 417 -2458 451 -2424
rect 485 -2458 519 -2424
rect 553 -2458 587 -2424
rect 621 -2458 655 -2424
rect 689 -2458 723 -2424
rect 757 -2458 791 -2424
rect 825 -2458 859 -2424
rect 893 -2458 927 -2424
rect 961 -2458 995 -2424
rect 1029 -2458 1063 -2424
rect 1097 -2458 1131 -2424
rect 1165 -2458 1199 -2424
rect 1233 -2458 1267 -2424
rect 1301 -2458 1335 -2424
rect 1369 -2458 1403 -2424
rect 1437 -2458 1471 -2424
rect 1505 -2458 1539 -2424
rect 1573 -2458 1607 -2424
rect 1641 -2458 1675 -2424
rect 1709 -2458 1743 -2424
rect 1777 -2458 1811 -2424
rect 1845 -2458 1879 -2424
rect 1913 -2458 1947 -2424
rect 1981 -2458 2015 -2424
rect 2049 -2458 2083 -2424
rect 2117 -2458 2151 -2424
rect 2185 -2458 2219 -2424
rect 2253 -2458 2287 -2424
rect 2321 -2458 2355 -2424
rect 2389 -2458 2423 -2424
rect 2457 -2458 2491 -2424
rect 2525 -2458 2559 -2424
rect 2593 -2458 2627 -2424
rect 2661 -2458 2695 -2424
rect 2729 -2458 2763 -2424
rect 2797 -2458 2831 -2424
rect 2865 -2458 2899 -2424
rect 2933 -2458 2967 -2424
rect 3001 -2458 3035 -2424
rect 3069 -2458 3103 -2424
rect 3137 -2458 3171 -2424
rect 3295 -2458 3329 -2424
rect -244 -2526 -210 -2492
rect -244 -2594 -210 -2560
rect -244 -2662 -210 -2628
rect 3295 -2526 3329 -2492
rect 3295 -2594 3329 -2560
rect 3295 -2662 3329 -2628
rect -244 -2730 -210 -2696
rect -244 -2798 -210 -2764
rect -244 -2866 -210 -2832
rect -244 -2934 -210 -2900
rect 3295 -2730 3329 -2696
rect 3295 -2798 3329 -2764
rect 3295 -2866 3329 -2832
rect 3295 -2934 3329 -2900
rect -59 -3075 -25 -3041
rect 9 -3075 43 -3041
rect 77 -3075 111 -3041
rect 145 -3075 179 -3041
rect 213 -3075 247 -3041
rect 281 -3075 315 -3041
rect 349 -3075 383 -3041
rect 417 -3075 451 -3041
rect 485 -3075 519 -3041
rect 553 -3075 587 -3041
rect 621 -3075 655 -3041
rect 689 -3075 723 -3041
rect 757 -3075 791 -3041
rect 825 -3075 859 -3041
rect 893 -3075 927 -3041
rect 961 -3075 995 -3041
rect 1029 -3075 1063 -3041
rect 1097 -3075 1131 -3041
rect 1165 -3075 1199 -3041
rect 1233 -3075 1267 -3041
rect 1301 -3075 1335 -3041
rect 1369 -3075 1403 -3041
rect 1437 -3075 1471 -3041
rect 1505 -3075 1539 -3041
rect 1573 -3075 1607 -3041
rect 1641 -3075 1675 -3041
rect 1709 -3075 1743 -3041
rect 1777 -3075 1811 -3041
rect 1845 -3075 1879 -3041
rect 1913 -3075 1947 -3041
rect 1981 -3075 2015 -3041
rect 2049 -3075 2083 -3041
rect 2117 -3075 2151 -3041
rect 2185 -3075 2219 -3041
rect 2253 -3075 2287 -3041
rect 2321 -3075 2355 -3041
rect 2389 -3075 2423 -3041
rect 2457 -3075 2491 -3041
rect 2525 -3075 2559 -3041
rect 2593 -3075 2627 -3041
rect 2661 -3075 2695 -3041
rect 2729 -3075 2763 -3041
rect 2797 -3075 2831 -3041
rect 2865 -3075 2899 -3041
rect 2933 -3075 2967 -3041
rect 3001 -3075 3035 -3041
rect 3069 -3075 3103 -3041
rect 3137 -3075 3171 -3041
<< poly >>
rect -84 890 116 906
rect -84 856 -35 890
rect -1 856 33 890
rect 67 856 116 890
rect -84 818 116 856
rect 421 890 621 906
rect 421 856 470 890
rect 504 856 538 890
rect 572 856 621 890
rect 421 818 621 856
rect 679 890 879 906
rect 679 856 728 890
rect 762 856 796 890
rect 830 856 879 890
rect 679 818 879 856
rect 1184 890 1384 906
rect 1184 856 1233 890
rect 1267 856 1301 890
rect 1335 856 1384 890
rect 1184 818 1384 856
rect 1442 890 1642 906
rect 1442 856 1491 890
rect 1525 856 1559 890
rect 1593 856 1642 890
rect 1442 818 1642 856
rect 1700 890 1900 906
rect 1700 856 1749 890
rect 1783 856 1817 890
rect 1851 856 1900 890
rect 1700 818 1900 856
rect 2205 890 2405 906
rect 2205 856 2254 890
rect 2288 856 2322 890
rect 2356 856 2405 890
rect 2205 818 2405 856
rect 2463 890 2663 906
rect 2463 856 2512 890
rect 2546 856 2580 890
rect 2614 856 2663 890
rect 2463 818 2663 856
rect 2969 890 3169 906
rect 2969 856 3018 890
rect 3052 856 3086 890
rect 3120 856 3169 890
rect 2969 818 3169 856
rect -84 592 116 618
rect 421 592 621 618
rect 679 592 879 618
rect 1184 592 1384 618
rect 1442 592 1642 618
rect 1700 592 1900 618
rect 2205 592 2405 618
rect 2463 592 2663 618
rect 2969 592 3169 618
rect -84 92 116 118
rect 421 92 621 118
rect 679 92 879 118
rect 1184 92 1384 118
rect 1442 92 1642 118
rect 1700 92 1900 118
rect 2205 92 2405 118
rect 2463 92 2663 118
rect 2969 92 3169 118
rect -84 -146 116 -108
rect -84 -180 -35 -146
rect -1 -180 33 -146
rect 67 -180 116 -146
rect -84 -196 116 -180
rect 421 -146 621 -108
rect 421 -180 470 -146
rect 504 -180 538 -146
rect 572 -180 621 -146
rect 421 -196 621 -180
rect 679 -146 879 -108
rect 679 -180 728 -146
rect 762 -180 796 -146
rect 830 -180 879 -146
rect 679 -196 879 -180
rect 1184 -146 1384 -108
rect 1184 -180 1233 -146
rect 1267 -180 1301 -146
rect 1335 -180 1384 -146
rect 1184 -196 1384 -180
rect 1442 -146 1642 -108
rect 1442 -180 1491 -146
rect 1525 -180 1559 -146
rect 1593 -180 1642 -146
rect 1442 -196 1642 -180
rect 1700 -146 1900 -108
rect 1700 -180 1749 -146
rect 1783 -180 1817 -146
rect 1851 -180 1900 -146
rect 1700 -196 1900 -180
rect 2205 -146 2405 -108
rect 2205 -180 2254 -146
rect 2288 -180 2322 -146
rect 2356 -180 2405 -146
rect 2205 -196 2405 -180
rect 2463 -146 2663 -108
rect 2463 -180 2512 -146
rect 2546 -180 2580 -146
rect 2614 -180 2663 -146
rect 2463 -196 2663 -180
rect 2969 -146 3169 -108
rect 2969 -180 3018 -146
rect 3052 -180 3086 -146
rect 3120 -180 3169 -146
rect 2969 -196 3169 -180
rect -84 -509 116 -493
rect -84 -543 -35 -509
rect -1 -543 33 -509
rect 67 -543 116 -509
rect -84 -581 116 -543
rect 421 -509 621 -493
rect 421 -543 470 -509
rect 504 -543 538 -509
rect 572 -543 621 -509
rect 421 -581 621 -543
rect 679 -509 879 -493
rect 679 -543 728 -509
rect 762 -543 796 -509
rect 830 -543 879 -509
rect 679 -581 879 -543
rect 1184 -509 1384 -493
rect 1184 -543 1233 -509
rect 1267 -543 1301 -509
rect 1335 -543 1384 -509
rect 1184 -581 1384 -543
rect 1442 -509 1642 -493
rect 1442 -543 1491 -509
rect 1525 -543 1559 -509
rect 1593 -543 1642 -509
rect 1442 -581 1642 -543
rect 1700 -509 1900 -493
rect 1700 -543 1749 -509
rect 1783 -543 1817 -509
rect 1851 -543 1900 -509
rect 1700 -581 1900 -543
rect 2205 -509 2405 -493
rect 2205 -543 2254 -509
rect 2288 -543 2322 -509
rect 2356 -543 2405 -509
rect 2205 -581 2405 -543
rect 2463 -509 2663 -493
rect 2463 -543 2512 -509
rect 2546 -543 2580 -509
rect 2614 -543 2663 -509
rect 2463 -581 2663 -543
rect 2969 -509 3169 -493
rect 2969 -543 3018 -509
rect 3052 -543 3086 -509
rect 3120 -543 3169 -509
rect 2969 -581 3169 -543
rect -84 -807 116 -781
rect 421 -807 621 -781
rect 679 -807 879 -781
rect 1184 -807 1384 -781
rect 1442 -807 1642 -781
rect 1700 -807 1900 -781
rect 2205 -807 2405 -781
rect 2463 -807 2663 -781
rect 2969 -807 3169 -781
rect -84 -1305 116 -1279
rect 421 -1305 621 -1279
rect 679 -1305 879 -1279
rect 1184 -1305 1384 -1279
rect 1442 -1305 1642 -1279
rect 1700 -1305 1900 -1279
rect 2205 -1305 2405 -1279
rect 2463 -1305 2663 -1279
rect 2969 -1305 3169 -1279
rect -84 -1543 116 -1505
rect -84 -1577 -35 -1543
rect -1 -1577 33 -1543
rect 67 -1577 116 -1543
rect -84 -1593 116 -1577
rect 421 -1543 621 -1505
rect 421 -1577 470 -1543
rect 504 -1577 538 -1543
rect 572 -1577 621 -1543
rect 421 -1593 621 -1577
rect 679 -1543 879 -1505
rect 679 -1577 728 -1543
rect 762 -1577 796 -1543
rect 830 -1577 879 -1543
rect 679 -1593 879 -1577
rect 1184 -1543 1384 -1505
rect 1184 -1577 1233 -1543
rect 1267 -1577 1301 -1543
rect 1335 -1577 1384 -1543
rect 1184 -1593 1384 -1577
rect 1442 -1543 1642 -1505
rect 1442 -1577 1491 -1543
rect 1525 -1577 1559 -1543
rect 1593 -1577 1642 -1543
rect 1442 -1593 1642 -1577
rect 1700 -1543 1900 -1505
rect 1700 -1577 1749 -1543
rect 1783 -1577 1817 -1543
rect 1851 -1577 1900 -1543
rect 1700 -1593 1900 -1577
rect 2205 -1543 2405 -1505
rect 2205 -1577 2254 -1543
rect 2288 -1577 2322 -1543
rect 2356 -1577 2405 -1543
rect 2205 -1593 2405 -1577
rect 2463 -1543 2663 -1505
rect 2463 -1577 2512 -1543
rect 2546 -1577 2580 -1543
rect 2614 -1577 2663 -1543
rect 2463 -1593 2663 -1577
rect 2969 -1543 3169 -1505
rect 2969 -1577 3018 -1543
rect 3052 -1577 3086 -1543
rect 3120 -1577 3169 -1543
rect 2969 -1593 3169 -1577
rect -84 -1906 116 -1890
rect -84 -1940 -35 -1906
rect -1 -1940 33 -1906
rect 67 -1940 116 -1906
rect -84 -1978 116 -1940
rect 421 -1906 621 -1890
rect 421 -1940 470 -1906
rect 504 -1940 538 -1906
rect 572 -1940 621 -1906
rect 421 -1978 621 -1940
rect 679 -1906 879 -1890
rect 679 -1940 728 -1906
rect 762 -1940 796 -1906
rect 830 -1940 879 -1906
rect 679 -1978 879 -1940
rect 1184 -1906 1384 -1890
rect 1184 -1940 1233 -1906
rect 1267 -1940 1301 -1906
rect 1335 -1940 1384 -1906
rect 1184 -1978 1384 -1940
rect 1442 -1906 1642 -1890
rect 1442 -1940 1491 -1906
rect 1525 -1940 1559 -1906
rect 1593 -1940 1642 -1906
rect 1442 -1978 1642 -1940
rect 1700 -1906 1900 -1890
rect 1700 -1940 1749 -1906
rect 1783 -1940 1817 -1906
rect 1851 -1940 1900 -1906
rect 1700 -1978 1900 -1940
rect 2205 -1906 2405 -1890
rect 2205 -1940 2254 -1906
rect 2288 -1940 2322 -1906
rect 2356 -1940 2405 -1906
rect 2205 -1978 2405 -1940
rect 2463 -1906 2663 -1890
rect 2463 -1940 2512 -1906
rect 2546 -1940 2580 -1906
rect 2614 -1940 2663 -1906
rect 2463 -1978 2663 -1940
rect 2969 -1906 3169 -1890
rect 2969 -1940 3018 -1906
rect 3052 -1940 3086 -1906
rect 3120 -1940 3169 -1906
rect 2969 -1978 3169 -1940
rect -84 -2204 116 -2178
rect 421 -2204 621 -2178
rect 679 -2204 879 -2178
rect 1184 -2204 1384 -2178
rect 1442 -2204 1642 -2178
rect 1700 -2204 1900 -2178
rect 2205 -2204 2405 -2178
rect 2463 -2204 2663 -2178
rect 2969 -2204 3169 -2178
rect -84 -2704 116 -2678
rect 421 -2704 621 -2678
rect 679 -2704 879 -2678
rect 1184 -2704 1384 -2678
rect 1442 -2704 1642 -2678
rect 1700 -2704 1900 -2678
rect 2205 -2704 2405 -2678
rect 2463 -2704 2663 -2678
rect 2969 -2704 3169 -2678
rect -84 -2942 116 -2904
rect -84 -2976 -35 -2942
rect -1 -2976 33 -2942
rect 67 -2976 116 -2942
rect -84 -2992 116 -2976
rect 421 -2942 621 -2904
rect 421 -2976 470 -2942
rect 504 -2976 538 -2942
rect 572 -2976 621 -2942
rect 421 -2992 621 -2976
rect 679 -2942 879 -2904
rect 679 -2976 728 -2942
rect 762 -2976 796 -2942
rect 830 -2976 879 -2942
rect 679 -2992 879 -2976
rect 1184 -2942 1384 -2904
rect 1184 -2976 1233 -2942
rect 1267 -2976 1301 -2942
rect 1335 -2976 1384 -2942
rect 1184 -2992 1384 -2976
rect 1442 -2942 1642 -2904
rect 1442 -2976 1491 -2942
rect 1525 -2976 1559 -2942
rect 1593 -2976 1642 -2942
rect 1442 -2992 1642 -2976
rect 1700 -2942 1900 -2904
rect 1700 -2976 1749 -2942
rect 1783 -2976 1817 -2942
rect 1851 -2976 1900 -2942
rect 1700 -2992 1900 -2976
rect 2205 -2942 2405 -2904
rect 2205 -2976 2254 -2942
rect 2288 -2976 2322 -2942
rect 2356 -2976 2405 -2942
rect 2205 -2992 2405 -2976
rect 2463 -2942 2663 -2904
rect 2463 -2976 2512 -2942
rect 2546 -2976 2580 -2942
rect 2614 -2976 2663 -2942
rect 2463 -2992 2663 -2976
rect 2969 -2942 3169 -2904
rect 2969 -2976 3018 -2942
rect 3052 -2976 3086 -2942
rect 3120 -2976 3169 -2942
rect 2969 -2992 3169 -2976
<< polycont >>
rect -35 856 -1 890
rect 33 856 67 890
rect 470 856 504 890
rect 538 856 572 890
rect 728 856 762 890
rect 796 856 830 890
rect 1233 856 1267 890
rect 1301 856 1335 890
rect 1491 856 1525 890
rect 1559 856 1593 890
rect 1749 856 1783 890
rect 1817 856 1851 890
rect 2254 856 2288 890
rect 2322 856 2356 890
rect 2512 856 2546 890
rect 2580 856 2614 890
rect 3018 856 3052 890
rect 3086 856 3120 890
rect -35 -180 -1 -146
rect 33 -180 67 -146
rect 470 -180 504 -146
rect 538 -180 572 -146
rect 728 -180 762 -146
rect 796 -180 830 -146
rect 1233 -180 1267 -146
rect 1301 -180 1335 -146
rect 1491 -180 1525 -146
rect 1559 -180 1593 -146
rect 1749 -180 1783 -146
rect 1817 -180 1851 -146
rect 2254 -180 2288 -146
rect 2322 -180 2356 -146
rect 2512 -180 2546 -146
rect 2580 -180 2614 -146
rect 3018 -180 3052 -146
rect 3086 -180 3120 -146
rect -35 -543 -1 -509
rect 33 -543 67 -509
rect 470 -543 504 -509
rect 538 -543 572 -509
rect 728 -543 762 -509
rect 796 -543 830 -509
rect 1233 -543 1267 -509
rect 1301 -543 1335 -509
rect 1491 -543 1525 -509
rect 1559 -543 1593 -509
rect 1749 -543 1783 -509
rect 1817 -543 1851 -509
rect 2254 -543 2288 -509
rect 2322 -543 2356 -509
rect 2512 -543 2546 -509
rect 2580 -543 2614 -509
rect 3018 -543 3052 -509
rect 3086 -543 3120 -509
rect -35 -1577 -1 -1543
rect 33 -1577 67 -1543
rect 470 -1577 504 -1543
rect 538 -1577 572 -1543
rect 728 -1577 762 -1543
rect 796 -1577 830 -1543
rect 1233 -1577 1267 -1543
rect 1301 -1577 1335 -1543
rect 1491 -1577 1525 -1543
rect 1559 -1577 1593 -1543
rect 1749 -1577 1783 -1543
rect 1817 -1577 1851 -1543
rect 2254 -1577 2288 -1543
rect 2322 -1577 2356 -1543
rect 2512 -1577 2546 -1543
rect 2580 -1577 2614 -1543
rect 3018 -1577 3052 -1543
rect 3086 -1577 3120 -1543
rect -35 -1940 -1 -1906
rect 33 -1940 67 -1906
rect 470 -1940 504 -1906
rect 538 -1940 572 -1906
rect 728 -1940 762 -1906
rect 796 -1940 830 -1906
rect 1233 -1940 1267 -1906
rect 1301 -1940 1335 -1906
rect 1491 -1940 1525 -1906
rect 1559 -1940 1593 -1906
rect 1749 -1940 1783 -1906
rect 1817 -1940 1851 -1906
rect 2254 -1940 2288 -1906
rect 2322 -1940 2356 -1906
rect 2512 -1940 2546 -1906
rect 2580 -1940 2614 -1906
rect 3018 -1940 3052 -1906
rect 3086 -1940 3120 -1906
rect -35 -2976 -1 -2942
rect 33 -2976 67 -2942
rect 470 -2976 504 -2942
rect 538 -2976 572 -2942
rect 728 -2976 762 -2942
rect 796 -2976 830 -2942
rect 1233 -2976 1267 -2942
rect 1301 -2976 1335 -2942
rect 1491 -2976 1525 -2942
rect 1559 -2976 1593 -2942
rect 1749 -2976 1783 -2942
rect 1817 -2976 1851 -2942
rect 2254 -2976 2288 -2942
rect 2322 -2976 2356 -2942
rect 2512 -2976 2546 -2942
rect 2580 -2976 2614 -2942
rect 3018 -2976 3052 -2942
rect 3086 -2976 3120 -2942
<< locali >>
rect -244 955 -80 989
rect -25 955 -8 989
rect 43 955 64 989
rect 111 955 136 989
rect 179 955 208 989
rect 247 955 280 989
rect 315 955 349 989
rect 386 955 417 989
rect 458 955 485 989
rect 530 955 553 989
rect 602 955 621 989
rect 674 955 689 989
rect 746 955 757 989
rect 818 955 825 989
rect 890 955 893 989
rect 927 955 928 989
rect 995 955 1000 989
rect 1063 955 1072 989
rect 1131 955 1144 989
rect 1199 955 1216 989
rect 1267 955 1288 989
rect 1335 955 1360 989
rect 1403 955 1432 989
rect 1471 955 1504 989
rect 1539 955 1573 989
rect 1610 955 1641 989
rect 1682 955 1709 989
rect 1754 955 1777 989
rect 1826 955 1845 989
rect 1898 955 1913 989
rect 1970 955 1981 989
rect 2042 955 2049 989
rect 2114 955 2117 989
rect 2151 955 2152 989
rect 2219 955 2224 989
rect 2287 955 2296 989
rect 2355 955 2368 989
rect 2423 955 2440 989
rect 2491 955 2512 989
rect 2559 955 2584 989
rect 2627 955 2656 989
rect 2695 955 2728 989
rect 2763 955 2797 989
rect 2834 955 2865 989
rect 2906 955 2933 989
rect 2978 955 3001 989
rect 3050 955 3069 989
rect 3122 955 3137 989
rect 3194 955 3329 989
rect -244 882 -210 955
rect -84 856 -37 890
rect -1 856 33 890
rect 69 856 116 890
rect 421 856 468 890
rect 504 856 538 890
rect 574 856 621 890
rect 679 856 726 890
rect 762 856 796 890
rect 832 856 879 890
rect 1184 856 1231 890
rect 1267 856 1301 890
rect 1337 856 1384 890
rect 1442 856 1489 890
rect 1525 856 1559 890
rect 1595 856 1642 890
rect 1700 856 1747 890
rect 1783 856 1817 890
rect 1853 856 1900 890
rect 2205 856 2252 890
rect 2288 856 2322 890
rect 2358 856 2405 890
rect 2463 856 2510 890
rect 2546 856 2580 890
rect 2616 856 2663 890
rect 2969 856 3016 890
rect 3052 856 3086 890
rect 3122 856 3169 890
rect 3295 882 3329 955
rect -244 810 -210 814
rect -244 738 -210 746
rect -244 666 -210 678
rect -130 803 -96 822
rect -130 735 -96 737
rect -130 699 -96 701
rect -130 614 -96 633
rect 128 803 162 822
rect 128 735 162 737
rect 128 699 162 701
rect 128 614 162 633
rect 375 803 409 822
rect 375 735 409 737
rect 375 699 409 701
rect 375 614 409 633
rect 633 803 667 822
rect 633 735 667 737
rect 633 699 667 701
rect 633 614 667 633
rect 891 803 925 822
rect 891 735 925 737
rect 891 699 925 701
rect 891 614 925 633
rect 1138 803 1172 822
rect 1138 735 1172 737
rect 1138 699 1172 701
rect 1138 614 1172 633
rect 1396 803 1430 822
rect 1396 735 1430 737
rect 1396 699 1430 701
rect 1396 614 1430 633
rect 1654 803 1688 822
rect 1654 735 1688 737
rect 1654 699 1688 701
rect 1654 614 1688 633
rect 1912 803 1946 822
rect 1912 735 1946 737
rect 1912 699 1946 701
rect 1912 614 1946 633
rect 2159 803 2193 822
rect 2159 735 2193 737
rect 2159 699 2193 701
rect 2159 614 2193 633
rect 2417 803 2451 822
rect 2417 735 2451 737
rect 2417 699 2451 701
rect 2417 614 2451 633
rect 2675 803 2709 822
rect 2675 735 2709 737
rect 2675 699 2709 701
rect 2675 614 2709 633
rect 2923 803 2957 822
rect 2923 735 2957 737
rect 2923 699 2957 701
rect 2923 614 2957 633
rect 3181 803 3215 822
rect 3181 735 3215 737
rect 3181 699 3215 701
rect 3181 614 3215 633
rect 3295 810 3329 814
rect 3295 738 3329 746
rect 3295 666 3329 678
rect -244 594 -210 610
rect -244 522 -210 542
rect -244 450 -210 474
rect -244 378 -210 406
rect 3295 594 3329 610
rect 3295 522 3329 542
rect 3295 450 3329 474
rect 3295 378 3329 406
rect -210 338 -59 372
rect -25 338 9 372
rect 43 338 77 372
rect 111 338 145 372
rect 179 338 213 372
rect 247 338 281 372
rect 315 338 349 372
rect 383 338 417 372
rect 451 338 485 372
rect 519 338 553 372
rect 587 338 621 372
rect 655 338 689 372
rect 723 338 757 372
rect 791 338 825 372
rect 859 338 893 372
rect 927 338 961 372
rect 995 338 1029 372
rect 1063 338 1097 372
rect 1131 338 1165 372
rect 1199 338 1233 372
rect 1267 338 1301 372
rect 1335 338 1369 372
rect 1403 338 1437 372
rect 1471 338 1505 372
rect 1539 338 1573 372
rect 1607 338 1641 372
rect 1675 338 1709 372
rect 1743 338 1777 372
rect 1811 338 1845 372
rect 1879 338 1913 372
rect 1947 338 1981 372
rect 2015 338 2049 372
rect 2083 338 2117 372
rect 2151 338 2185 372
rect 2219 338 2253 372
rect 2287 338 2321 372
rect 2355 338 2389 372
rect 2423 338 2457 372
rect 2491 338 2525 372
rect 2559 338 2593 372
rect 2627 338 2661 372
rect 2695 338 2729 372
rect 2763 338 2797 372
rect 2831 338 2865 372
rect 2899 338 2933 372
rect 2967 338 3001 372
rect 3035 338 3069 372
rect 3103 338 3137 372
rect 3171 338 3295 372
rect -244 306 -210 338
rect -244 236 -210 270
rect -244 168 -210 200
rect -244 100 -210 128
rect 3295 306 3329 338
rect 3295 236 3329 270
rect 3295 168 3329 200
rect 3295 100 3329 128
rect -244 32 -210 56
rect -244 -36 -210 -16
rect -244 -104 -210 -88
rect -130 77 -96 96
rect -130 9 -96 11
rect -130 -27 -96 -25
rect -130 -112 -96 -93
rect 128 77 162 96
rect 128 9 162 11
rect 128 -27 162 -25
rect 128 -112 162 -93
rect 375 77 409 96
rect 375 9 409 11
rect 375 -27 409 -25
rect 375 -112 409 -93
rect 633 77 667 96
rect 633 9 667 11
rect 633 -27 667 -25
rect 633 -112 667 -93
rect 891 77 925 96
rect 891 9 925 11
rect 891 -27 925 -25
rect 891 -112 925 -93
rect 1138 77 1172 96
rect 1138 9 1172 11
rect 1138 -27 1172 -25
rect 1138 -112 1172 -93
rect 1396 77 1430 96
rect 1396 9 1430 11
rect 1396 -27 1430 -25
rect 1396 -112 1430 -93
rect 1654 77 1688 96
rect 1654 9 1688 11
rect 1654 -27 1688 -25
rect 1654 -112 1688 -93
rect 1912 77 1946 96
rect 1912 9 1946 11
rect 1912 -27 1946 -25
rect 1912 -112 1946 -93
rect 2159 77 2193 96
rect 2159 9 2193 11
rect 2159 -27 2193 -25
rect 2159 -112 2193 -93
rect 2417 77 2451 96
rect 2417 9 2451 11
rect 2417 -27 2451 -25
rect 2417 -112 2451 -93
rect 2675 77 2709 96
rect 2675 9 2709 11
rect 2675 -27 2709 -25
rect 2675 -112 2709 -93
rect 2923 77 2957 96
rect 2923 9 2957 11
rect 2923 -27 2957 -25
rect 2923 -112 2957 -93
rect 3181 77 3215 96
rect 3181 9 3215 11
rect 3181 -27 3215 -25
rect 3181 -112 3215 -93
rect 3295 32 3329 56
rect 3295 -36 3329 -16
rect 3295 -104 3329 -88
rect -244 -172 -210 -160
rect -84 -180 -37 -146
rect -1 -180 33 -146
rect 69 -180 116 -146
rect 421 -180 468 -146
rect 504 -180 538 -146
rect 574 -180 621 -146
rect 679 -180 726 -146
rect 762 -180 796 -146
rect 832 -180 879 -146
rect 1184 -180 1231 -146
rect 1267 -180 1301 -146
rect 1337 -180 1384 -146
rect 1442 -180 1489 -146
rect 1525 -180 1559 -146
rect 1595 -180 1642 -146
rect 1700 -180 1747 -146
rect 1783 -180 1817 -146
rect 1853 -180 1900 -146
rect 2205 -180 2252 -146
rect 2288 -180 2322 -146
rect 2358 -180 2405 -146
rect 2463 -180 2510 -146
rect 2546 -180 2580 -146
rect 2616 -180 2663 -146
rect 2969 -180 3016 -146
rect 3052 -180 3086 -146
rect 3122 -180 3169 -146
rect 3295 -172 3329 -160
rect -244 -240 -210 -232
rect -244 -308 -210 -304
rect -244 -414 -210 -410
rect -244 -486 -210 -478
rect 3295 -240 3329 -232
rect 3295 -308 3329 -304
rect 3295 -414 3329 -410
rect 3295 -486 3329 -478
rect -84 -543 -37 -509
rect -1 -543 33 -509
rect 69 -543 116 -509
rect 421 -543 468 -509
rect 504 -543 538 -509
rect 574 -543 621 -509
rect 679 -543 726 -509
rect 762 -543 796 -509
rect 832 -543 879 -509
rect 1184 -543 1231 -509
rect 1267 -543 1301 -509
rect 1337 -543 1384 -509
rect 1442 -543 1489 -509
rect 1525 -543 1559 -509
rect 1595 -543 1642 -509
rect 1700 -543 1747 -509
rect 1783 -543 1817 -509
rect 1853 -543 1900 -509
rect 2205 -543 2252 -509
rect 2288 -543 2322 -509
rect 2358 -543 2405 -509
rect 2463 -543 2510 -509
rect 2546 -543 2580 -509
rect 2616 -543 2663 -509
rect 2969 -543 3016 -509
rect 3052 -543 3086 -509
rect 3122 -543 3169 -509
rect -244 -558 -210 -546
rect 3295 -558 3329 -546
rect -244 -630 -210 -614
rect -244 -702 -210 -682
rect -244 -774 -210 -750
rect -130 -596 -96 -577
rect -130 -664 -96 -662
rect -130 -700 -96 -698
rect -130 -785 -96 -766
rect 128 -596 162 -577
rect 128 -664 162 -662
rect 128 -700 162 -698
rect 128 -785 162 -766
rect 375 -596 409 -577
rect 375 -664 409 -662
rect 375 -700 409 -698
rect 375 -785 409 -766
rect 633 -596 667 -577
rect 633 -664 667 -662
rect 633 -700 667 -698
rect 633 -785 667 -766
rect 891 -596 925 -577
rect 891 -664 925 -662
rect 891 -700 925 -698
rect 891 -785 925 -766
rect 1138 -596 1172 -577
rect 1138 -664 1172 -662
rect 1138 -700 1172 -698
rect 1138 -785 1172 -766
rect 1396 -596 1430 -577
rect 1396 -664 1430 -662
rect 1396 -700 1430 -698
rect 1396 -785 1430 -766
rect 1654 -596 1688 -577
rect 1654 -664 1688 -662
rect 1654 -700 1688 -698
rect 1654 -785 1688 -766
rect 1912 -596 1946 -577
rect 1912 -664 1946 -662
rect 1912 -700 1946 -698
rect 1912 -785 1946 -766
rect 2159 -596 2193 -577
rect 2159 -664 2193 -662
rect 2159 -700 2193 -698
rect 2159 -785 2193 -766
rect 2417 -596 2451 -577
rect 2417 -664 2451 -662
rect 2417 -700 2451 -698
rect 2417 -785 2451 -766
rect 2675 -596 2709 -577
rect 2675 -664 2709 -662
rect 2675 -700 2709 -698
rect 2675 -785 2709 -766
rect 2923 -596 2957 -577
rect 2923 -664 2957 -662
rect 2923 -700 2957 -698
rect 2923 -785 2957 -766
rect 3181 -596 3215 -577
rect 3181 -664 3215 -662
rect 3181 -700 3215 -698
rect 3181 -785 3215 -766
rect 3295 -630 3329 -614
rect 3295 -702 3329 -682
rect 3295 -774 3329 -750
rect -244 -846 -210 -818
rect -244 -918 -210 -886
rect -244 -990 -210 -952
rect -244 -1026 -210 -1024
rect 3295 -846 3329 -818
rect 3295 -918 3329 -886
rect 3295 -990 3329 -952
rect 3295 -1026 3329 -1024
rect -244 -1060 -59 -1026
rect -25 -1060 9 -1026
rect 43 -1060 77 -1026
rect 111 -1060 145 -1026
rect 179 -1060 213 -1026
rect 247 -1060 281 -1026
rect 315 -1060 349 -1026
rect 383 -1060 417 -1026
rect 451 -1060 485 -1026
rect 519 -1060 553 -1026
rect 587 -1060 621 -1026
rect 655 -1060 689 -1026
rect 723 -1060 757 -1026
rect 791 -1060 825 -1026
rect 859 -1060 893 -1026
rect 927 -1060 961 -1026
rect 995 -1060 1029 -1026
rect 1063 -1060 1097 -1026
rect 1131 -1060 1165 -1026
rect 1199 -1060 1233 -1026
rect 1267 -1060 1301 -1026
rect 1335 -1060 1369 -1026
rect 1403 -1060 1437 -1026
rect 1471 -1060 1505 -1026
rect 1539 -1060 1573 -1026
rect 1607 -1060 1641 -1026
rect 1675 -1060 1709 -1026
rect 1743 -1060 1777 -1026
rect 1811 -1060 1845 -1026
rect 1879 -1060 1913 -1026
rect 1947 -1060 1981 -1026
rect 2015 -1060 2049 -1026
rect 2083 -1060 2117 -1026
rect 2151 -1060 2185 -1026
rect 2219 -1060 2253 -1026
rect 2287 -1060 2321 -1026
rect 2355 -1060 2389 -1026
rect 2423 -1060 2457 -1026
rect 2491 -1060 2525 -1026
rect 2559 -1060 2593 -1026
rect 2627 -1060 2661 -1026
rect 2695 -1060 2729 -1026
rect 2763 -1060 2797 -1026
rect 2831 -1060 2865 -1026
rect 2899 -1060 2933 -1026
rect 2967 -1060 3001 -1026
rect 3035 -1060 3069 -1026
rect 3103 -1060 3137 -1026
rect 3171 -1060 3329 -1026
rect -244 -1062 -210 -1060
rect -244 -1134 -210 -1096
rect -244 -1200 -210 -1168
rect -244 -1268 -210 -1240
rect 3295 -1062 3329 -1060
rect 3295 -1134 3329 -1096
rect 3295 -1200 3329 -1168
rect 3295 -1268 3329 -1240
rect -244 -1336 -210 -1312
rect -244 -1404 -210 -1384
rect -244 -1472 -210 -1456
rect -130 -1320 -96 -1301
rect -130 -1388 -96 -1386
rect -130 -1424 -96 -1422
rect -130 -1509 -96 -1490
rect 128 -1320 162 -1301
rect 128 -1388 162 -1386
rect 128 -1424 162 -1422
rect 128 -1509 162 -1490
rect 375 -1320 409 -1301
rect 375 -1388 409 -1386
rect 375 -1424 409 -1422
rect 375 -1509 409 -1490
rect 633 -1320 667 -1301
rect 633 -1388 667 -1386
rect 633 -1424 667 -1422
rect 633 -1509 667 -1490
rect 891 -1320 925 -1301
rect 891 -1388 925 -1386
rect 891 -1424 925 -1422
rect 891 -1509 925 -1490
rect 1138 -1320 1172 -1301
rect 1138 -1388 1172 -1386
rect 1138 -1424 1172 -1422
rect 1138 -1509 1172 -1490
rect 1396 -1320 1430 -1301
rect 1396 -1388 1430 -1386
rect 1396 -1424 1430 -1422
rect 1396 -1509 1430 -1490
rect 1654 -1320 1688 -1301
rect 1654 -1388 1688 -1386
rect 1654 -1424 1688 -1422
rect 1654 -1509 1688 -1490
rect 1912 -1320 1946 -1301
rect 1912 -1388 1946 -1386
rect 1912 -1424 1946 -1422
rect 1912 -1509 1946 -1490
rect 2159 -1320 2193 -1301
rect 2159 -1388 2193 -1386
rect 2159 -1424 2193 -1422
rect 2159 -1509 2193 -1490
rect 2417 -1320 2451 -1301
rect 2417 -1388 2451 -1386
rect 2417 -1424 2451 -1422
rect 2417 -1509 2451 -1490
rect 2675 -1320 2709 -1301
rect 2675 -1388 2709 -1386
rect 2675 -1424 2709 -1422
rect 2675 -1509 2709 -1490
rect 2923 -1320 2957 -1301
rect 2923 -1388 2957 -1386
rect 2923 -1424 2957 -1422
rect 2923 -1509 2957 -1490
rect 3181 -1320 3215 -1301
rect 3181 -1388 3215 -1386
rect 3181 -1424 3215 -1422
rect 3181 -1509 3215 -1490
rect 3295 -1336 3329 -1312
rect 3295 -1404 3329 -1384
rect 3295 -1472 3329 -1456
rect -244 -1540 -210 -1528
rect 3295 -1540 3329 -1528
rect -84 -1577 -37 -1543
rect -1 -1577 33 -1543
rect 69 -1577 116 -1543
rect 421 -1577 468 -1543
rect 504 -1577 538 -1543
rect 574 -1577 621 -1543
rect 679 -1577 726 -1543
rect 762 -1577 796 -1543
rect 832 -1577 879 -1543
rect 1184 -1577 1231 -1543
rect 1267 -1577 1301 -1543
rect 1337 -1577 1384 -1543
rect 1442 -1577 1489 -1543
rect 1525 -1577 1559 -1543
rect 1595 -1577 1642 -1543
rect 1700 -1577 1747 -1543
rect 1783 -1577 1817 -1543
rect 1853 -1577 1900 -1543
rect 2205 -1577 2252 -1543
rect 2288 -1577 2322 -1543
rect 2358 -1577 2405 -1543
rect 2463 -1577 2510 -1543
rect 2546 -1577 2580 -1543
rect 2616 -1577 2663 -1543
rect 2969 -1577 3016 -1543
rect 3052 -1577 3086 -1543
rect 3122 -1577 3169 -1543
rect -244 -1608 -210 -1600
rect -244 -1676 -210 -1672
rect -244 -1782 -210 -1778
rect -244 -1854 -210 -1846
rect 3295 -1608 3329 -1600
rect 3295 -1676 3329 -1672
rect 3295 -1782 3329 -1778
rect 3295 -1854 3329 -1846
rect -244 -1926 -210 -1914
rect -84 -1940 -37 -1906
rect -1 -1940 33 -1906
rect 69 -1940 116 -1906
rect 421 -1940 468 -1906
rect 504 -1940 538 -1906
rect 574 -1940 621 -1906
rect 679 -1940 726 -1906
rect 762 -1940 796 -1906
rect 832 -1940 879 -1906
rect 1184 -1940 1231 -1906
rect 1267 -1940 1301 -1906
rect 1337 -1940 1384 -1906
rect 1442 -1940 1489 -1906
rect 1525 -1940 1559 -1906
rect 1595 -1940 1642 -1906
rect 1700 -1940 1747 -1906
rect 1783 -1940 1817 -1906
rect 1853 -1940 1900 -1906
rect 2205 -1940 2252 -1906
rect 2288 -1940 2322 -1906
rect 2358 -1940 2405 -1906
rect 2463 -1940 2510 -1906
rect 2546 -1940 2580 -1906
rect 2616 -1940 2663 -1906
rect 2969 -1940 3016 -1906
rect 3052 -1940 3086 -1906
rect 3122 -1940 3169 -1906
rect 3295 -1926 3329 -1914
rect -244 -1998 -210 -1982
rect -244 -2070 -210 -2050
rect -244 -2142 -210 -2118
rect -130 -1993 -96 -1974
rect -130 -2061 -96 -2059
rect -130 -2097 -96 -2095
rect -130 -2182 -96 -2163
rect 128 -1993 162 -1974
rect 128 -2061 162 -2059
rect 128 -2097 162 -2095
rect 128 -2182 162 -2163
rect 375 -1993 409 -1974
rect 375 -2061 409 -2059
rect 375 -2097 409 -2095
rect 375 -2182 409 -2163
rect 633 -1993 667 -1974
rect 633 -2061 667 -2059
rect 633 -2097 667 -2095
rect 633 -2182 667 -2163
rect 891 -1993 925 -1974
rect 891 -2061 925 -2059
rect 891 -2097 925 -2095
rect 891 -2182 925 -2163
rect 1138 -1993 1172 -1974
rect 1138 -2061 1172 -2059
rect 1138 -2097 1172 -2095
rect 1138 -2182 1172 -2163
rect 1396 -1993 1430 -1974
rect 1396 -2061 1430 -2059
rect 1396 -2097 1430 -2095
rect 1396 -2182 1430 -2163
rect 1654 -1993 1688 -1974
rect 1654 -2061 1688 -2059
rect 1654 -2097 1688 -2095
rect 1654 -2182 1688 -2163
rect 1912 -1993 1946 -1974
rect 1912 -2061 1946 -2059
rect 1912 -2097 1946 -2095
rect 1912 -2182 1946 -2163
rect 2159 -1993 2193 -1974
rect 2159 -2061 2193 -2059
rect 2159 -2097 2193 -2095
rect 2159 -2182 2193 -2163
rect 2417 -1993 2451 -1974
rect 2417 -2061 2451 -2059
rect 2417 -2097 2451 -2095
rect 2417 -2182 2451 -2163
rect 2675 -1993 2709 -1974
rect 2675 -2061 2709 -2059
rect 2675 -2097 2709 -2095
rect 2675 -2182 2709 -2163
rect 2923 -1993 2957 -1974
rect 2923 -2061 2957 -2059
rect 2923 -2097 2957 -2095
rect 2923 -2182 2957 -2163
rect 3181 -1993 3215 -1974
rect 3181 -2061 3215 -2059
rect 3181 -2097 3215 -2095
rect 3181 -2182 3215 -2163
rect 3295 -1998 3329 -1982
rect 3295 -2070 3329 -2050
rect 3295 -2142 3329 -2118
rect -244 -2214 -210 -2186
rect -244 -2286 -210 -2254
rect -244 -2356 -210 -2322
rect -244 -2424 -210 -2392
rect 3295 -2214 3329 -2186
rect 3295 -2286 3329 -2254
rect 3295 -2356 3329 -2322
rect 3295 -2424 3329 -2392
rect -210 -2458 -59 -2424
rect -25 -2458 9 -2424
rect 43 -2458 77 -2424
rect 111 -2458 145 -2424
rect 179 -2458 213 -2424
rect 247 -2458 281 -2424
rect 315 -2458 349 -2424
rect 383 -2458 417 -2424
rect 451 -2458 485 -2424
rect 519 -2458 553 -2424
rect 587 -2458 621 -2424
rect 655 -2458 689 -2424
rect 723 -2458 757 -2424
rect 791 -2458 825 -2424
rect 859 -2458 893 -2424
rect 927 -2458 961 -2424
rect 995 -2458 1029 -2424
rect 1063 -2458 1097 -2424
rect 1131 -2458 1165 -2424
rect 1199 -2458 1233 -2424
rect 1267 -2458 1301 -2424
rect 1335 -2458 1369 -2424
rect 1403 -2458 1437 -2424
rect 1471 -2458 1505 -2424
rect 1539 -2458 1573 -2424
rect 1607 -2458 1641 -2424
rect 1675 -2458 1709 -2424
rect 1743 -2458 1777 -2424
rect 1811 -2458 1845 -2424
rect 1879 -2458 1913 -2424
rect 1947 -2458 1981 -2424
rect 2015 -2458 2049 -2424
rect 2083 -2458 2117 -2424
rect 2151 -2458 2185 -2424
rect 2219 -2458 2253 -2424
rect 2287 -2458 2321 -2424
rect 2355 -2458 2389 -2424
rect 2423 -2458 2457 -2424
rect 2491 -2458 2525 -2424
rect 2559 -2458 2593 -2424
rect 2627 -2458 2661 -2424
rect 2695 -2458 2729 -2424
rect 2763 -2458 2797 -2424
rect 2831 -2458 2865 -2424
rect 2899 -2458 2933 -2424
rect 2967 -2458 3001 -2424
rect 3035 -2458 3069 -2424
rect 3103 -2458 3137 -2424
rect 3171 -2458 3295 -2424
rect -244 -2492 -210 -2464
rect -244 -2560 -210 -2536
rect -244 -2628 -210 -2608
rect -244 -2696 -210 -2680
rect 3295 -2492 3329 -2464
rect 3295 -2560 3329 -2536
rect 3295 -2628 3329 -2608
rect 3295 -2696 3329 -2680
rect -244 -2764 -210 -2752
rect -244 -2832 -210 -2824
rect -244 -2900 -210 -2896
rect -130 -2719 -96 -2700
rect -130 -2787 -96 -2785
rect -130 -2823 -96 -2821
rect -130 -2908 -96 -2889
rect 128 -2719 162 -2700
rect 128 -2787 162 -2785
rect 128 -2823 162 -2821
rect 128 -2908 162 -2889
rect 375 -2719 409 -2700
rect 375 -2787 409 -2785
rect 375 -2823 409 -2821
rect 375 -2908 409 -2889
rect 633 -2719 667 -2700
rect 633 -2787 667 -2785
rect 633 -2823 667 -2821
rect 633 -2908 667 -2889
rect 891 -2719 925 -2700
rect 891 -2787 925 -2785
rect 891 -2823 925 -2821
rect 891 -2908 925 -2889
rect 1138 -2719 1172 -2700
rect 1138 -2787 1172 -2785
rect 1138 -2823 1172 -2821
rect 1138 -2908 1172 -2889
rect 1396 -2719 1430 -2700
rect 1396 -2787 1430 -2785
rect 1396 -2823 1430 -2821
rect 1396 -2908 1430 -2889
rect 1654 -2719 1688 -2700
rect 1654 -2787 1688 -2785
rect 1654 -2823 1688 -2821
rect 1654 -2908 1688 -2889
rect 1912 -2719 1946 -2700
rect 1912 -2787 1946 -2785
rect 1912 -2823 1946 -2821
rect 1912 -2908 1946 -2889
rect 2159 -2719 2193 -2700
rect 2159 -2787 2193 -2785
rect 2159 -2823 2193 -2821
rect 2159 -2908 2193 -2889
rect 2417 -2719 2451 -2700
rect 2417 -2787 2451 -2785
rect 2417 -2823 2451 -2821
rect 2417 -2908 2451 -2889
rect 2675 -2719 2709 -2700
rect 2675 -2787 2709 -2785
rect 2675 -2823 2709 -2821
rect 2675 -2908 2709 -2889
rect 2923 -2719 2957 -2700
rect 2923 -2787 2957 -2785
rect 2923 -2823 2957 -2821
rect 2923 -2908 2957 -2889
rect 3181 -2719 3215 -2700
rect 3181 -2787 3215 -2785
rect 3181 -2823 3215 -2821
rect 3181 -2908 3215 -2889
rect 3295 -2764 3329 -2752
rect 3295 -2832 3329 -2824
rect 3295 -2900 3329 -2896
rect -244 -3041 -210 -2968
rect -84 -2976 -37 -2942
rect -1 -2976 33 -2942
rect 69 -2976 116 -2942
rect 421 -2976 468 -2942
rect 504 -2976 538 -2942
rect 574 -2976 621 -2942
rect 679 -2976 726 -2942
rect 762 -2976 796 -2942
rect 832 -2976 879 -2942
rect 1184 -2976 1231 -2942
rect 1267 -2976 1301 -2942
rect 1337 -2976 1384 -2942
rect 1442 -2976 1489 -2942
rect 1525 -2976 1559 -2942
rect 1595 -2976 1642 -2942
rect 1700 -2976 1747 -2942
rect 1783 -2976 1817 -2942
rect 1853 -2976 1900 -2942
rect 2205 -2976 2252 -2942
rect 2288 -2976 2322 -2942
rect 2358 -2976 2405 -2942
rect 2463 -2976 2510 -2942
rect 2546 -2976 2580 -2942
rect 2616 -2976 2663 -2942
rect 2969 -2976 3016 -2942
rect 3052 -2976 3086 -2942
rect 3122 -2976 3169 -2942
rect 3295 -3041 3329 -2968
rect -244 -3075 -80 -3041
rect -25 -3075 -8 -3041
rect 43 -3075 64 -3041
rect 111 -3075 136 -3041
rect 179 -3075 208 -3041
rect 247 -3075 280 -3041
rect 315 -3075 349 -3041
rect 386 -3075 417 -3041
rect 458 -3075 485 -3041
rect 530 -3075 553 -3041
rect 602 -3075 621 -3041
rect 674 -3075 689 -3041
rect 746 -3075 757 -3041
rect 818 -3075 825 -3041
rect 890 -3075 893 -3041
rect 927 -3075 928 -3041
rect 995 -3075 1000 -3041
rect 1063 -3075 1072 -3041
rect 1131 -3075 1144 -3041
rect 1199 -3075 1216 -3041
rect 1267 -3075 1288 -3041
rect 1335 -3075 1360 -3041
rect 1403 -3075 1432 -3041
rect 1471 -3075 1504 -3041
rect 1539 -3075 1573 -3041
rect 1610 -3075 1641 -3041
rect 1682 -3075 1709 -3041
rect 1754 -3075 1777 -3041
rect 1826 -3075 1845 -3041
rect 1898 -3075 1913 -3041
rect 1970 -3075 1981 -3041
rect 2042 -3075 2049 -3041
rect 2114 -3075 2117 -3041
rect 2151 -3075 2152 -3041
rect 2219 -3075 2224 -3041
rect 2287 -3075 2296 -3041
rect 2355 -3075 2368 -3041
rect 2423 -3075 2440 -3041
rect 2491 -3075 2512 -3041
rect 2559 -3075 2584 -3041
rect 2627 -3075 2656 -3041
rect 2695 -3075 2728 -3041
rect 2763 -3075 2797 -3041
rect 2834 -3075 2865 -3041
rect 2906 -3075 2933 -3041
rect 2978 -3075 3001 -3041
rect 3050 -3075 3069 -3041
rect 3122 -3075 3137 -3041
rect 3194 -3075 3329 -3041
<< viali >>
rect -80 955 -59 989
rect -59 955 -46 989
rect -8 955 9 989
rect 9 955 26 989
rect 64 955 77 989
rect 77 955 98 989
rect 136 955 145 989
rect 145 955 170 989
rect 208 955 213 989
rect 213 955 242 989
rect 280 955 281 989
rect 281 955 314 989
rect 352 955 383 989
rect 383 955 386 989
rect 424 955 451 989
rect 451 955 458 989
rect 496 955 519 989
rect 519 955 530 989
rect 568 955 587 989
rect 587 955 602 989
rect 640 955 655 989
rect 655 955 674 989
rect 712 955 723 989
rect 723 955 746 989
rect 784 955 791 989
rect 791 955 818 989
rect 856 955 859 989
rect 859 955 890 989
rect 928 955 961 989
rect 961 955 962 989
rect 1000 955 1029 989
rect 1029 955 1034 989
rect 1072 955 1097 989
rect 1097 955 1106 989
rect 1144 955 1165 989
rect 1165 955 1178 989
rect 1216 955 1233 989
rect 1233 955 1250 989
rect 1288 955 1301 989
rect 1301 955 1322 989
rect 1360 955 1369 989
rect 1369 955 1394 989
rect 1432 955 1437 989
rect 1437 955 1466 989
rect 1504 955 1505 989
rect 1505 955 1538 989
rect 1576 955 1607 989
rect 1607 955 1610 989
rect 1648 955 1675 989
rect 1675 955 1682 989
rect 1720 955 1743 989
rect 1743 955 1754 989
rect 1792 955 1811 989
rect 1811 955 1826 989
rect 1864 955 1879 989
rect 1879 955 1898 989
rect 1936 955 1947 989
rect 1947 955 1970 989
rect 2008 955 2015 989
rect 2015 955 2042 989
rect 2080 955 2083 989
rect 2083 955 2114 989
rect 2152 955 2185 989
rect 2185 955 2186 989
rect 2224 955 2253 989
rect 2253 955 2258 989
rect 2296 955 2321 989
rect 2321 955 2330 989
rect 2368 955 2389 989
rect 2389 955 2402 989
rect 2440 955 2457 989
rect 2457 955 2474 989
rect 2512 955 2525 989
rect 2525 955 2546 989
rect 2584 955 2593 989
rect 2593 955 2618 989
rect 2656 955 2661 989
rect 2661 955 2690 989
rect 2728 955 2729 989
rect 2729 955 2762 989
rect 2800 955 2831 989
rect 2831 955 2834 989
rect 2872 955 2899 989
rect 2899 955 2906 989
rect 2944 955 2967 989
rect 2967 955 2978 989
rect 3016 955 3035 989
rect 3035 955 3050 989
rect 3088 955 3103 989
rect 3103 955 3122 989
rect 3160 955 3171 989
rect 3171 955 3194 989
rect -244 848 -210 882
rect -37 856 -35 890
rect -35 856 -3 890
rect 35 856 67 890
rect 67 856 69 890
rect 468 856 470 890
rect 470 856 502 890
rect 540 856 572 890
rect 572 856 574 890
rect 726 856 728 890
rect 728 856 760 890
rect 798 856 830 890
rect 830 856 832 890
rect 1231 856 1233 890
rect 1233 856 1265 890
rect 1303 856 1335 890
rect 1335 856 1337 890
rect 1489 856 1491 890
rect 1491 856 1523 890
rect 1561 856 1593 890
rect 1593 856 1595 890
rect 1747 856 1749 890
rect 1749 856 1781 890
rect 1819 856 1851 890
rect 1851 856 1853 890
rect 2252 856 2254 890
rect 2254 856 2286 890
rect 2324 856 2356 890
rect 2356 856 2358 890
rect 2510 856 2512 890
rect 2512 856 2544 890
rect 2582 856 2614 890
rect 2614 856 2616 890
rect 3016 856 3018 890
rect 3018 856 3050 890
rect 3088 856 3120 890
rect 3120 856 3122 890
rect 3295 848 3329 882
rect -244 780 -210 810
rect -244 776 -210 780
rect -244 712 -210 738
rect -244 704 -210 712
rect -244 644 -210 666
rect -244 632 -210 644
rect -130 769 -96 771
rect -130 737 -96 769
rect -130 667 -96 699
rect -130 665 -96 667
rect 128 769 162 771
rect 128 737 162 769
rect 128 667 162 699
rect 128 665 162 667
rect 375 769 409 771
rect 375 737 409 769
rect 375 667 409 699
rect 375 665 409 667
rect 633 769 667 771
rect 633 737 667 769
rect 633 667 667 699
rect 633 665 667 667
rect 891 769 925 771
rect 891 737 925 769
rect 891 667 925 699
rect 891 665 925 667
rect 1138 769 1172 771
rect 1138 737 1172 769
rect 1138 667 1172 699
rect 1138 665 1172 667
rect 1396 769 1430 771
rect 1396 737 1430 769
rect 1396 667 1430 699
rect 1396 665 1430 667
rect 1654 769 1688 771
rect 1654 737 1688 769
rect 1654 667 1688 699
rect 1654 665 1688 667
rect 1912 769 1946 771
rect 1912 737 1946 769
rect 1912 667 1946 699
rect 1912 665 1946 667
rect 2159 769 2193 771
rect 2159 737 2193 769
rect 2159 667 2193 699
rect 2159 665 2193 667
rect 2417 769 2451 771
rect 2417 737 2451 769
rect 2417 667 2451 699
rect 2417 665 2451 667
rect 2675 769 2709 771
rect 2675 737 2709 769
rect 2675 667 2709 699
rect 2675 665 2709 667
rect 2923 769 2957 771
rect 2923 737 2957 769
rect 2923 667 2957 699
rect 2923 665 2957 667
rect 3181 769 3215 771
rect 3181 737 3215 769
rect 3181 667 3215 699
rect 3181 665 3215 667
rect 3295 780 3329 810
rect 3295 776 3329 780
rect 3295 712 3329 738
rect 3295 704 3329 712
rect 3295 644 3329 666
rect 3295 632 3329 644
rect -244 576 -210 594
rect -244 560 -210 576
rect -244 508 -210 522
rect -244 488 -210 508
rect -244 440 -210 450
rect -244 416 -210 440
rect -244 372 -210 378
rect 3295 576 3329 594
rect 3295 560 3329 576
rect 3295 508 3329 522
rect 3295 488 3329 508
rect 3295 440 3329 450
rect 3295 416 3329 440
rect 3295 372 3329 378
rect -244 344 -210 372
rect 3295 344 3329 372
rect -244 304 -210 306
rect -244 272 -210 304
rect -244 202 -210 234
rect -244 200 -210 202
rect -244 134 -210 162
rect -244 128 -210 134
rect 3295 304 3329 306
rect 3295 272 3329 304
rect 3295 202 3329 234
rect 3295 200 3329 202
rect 3295 134 3329 162
rect 3295 128 3329 134
rect -244 66 -210 90
rect -244 56 -210 66
rect -244 -2 -210 18
rect -244 -16 -210 -2
rect -244 -70 -210 -54
rect -244 -88 -210 -70
rect -130 43 -96 45
rect -130 11 -96 43
rect -130 -59 -96 -27
rect -130 -61 -96 -59
rect 128 43 162 45
rect 128 11 162 43
rect 128 -59 162 -27
rect 128 -61 162 -59
rect 375 43 409 45
rect 375 11 409 43
rect 375 -59 409 -27
rect 375 -61 409 -59
rect 633 43 667 45
rect 633 11 667 43
rect 633 -59 667 -27
rect 633 -61 667 -59
rect 891 43 925 45
rect 891 11 925 43
rect 891 -59 925 -27
rect 891 -61 925 -59
rect 1138 43 1172 45
rect 1138 11 1172 43
rect 1138 -59 1172 -27
rect 1138 -61 1172 -59
rect 1396 43 1430 45
rect 1396 11 1430 43
rect 1396 -59 1430 -27
rect 1396 -61 1430 -59
rect 1654 43 1688 45
rect 1654 11 1688 43
rect 1654 -59 1688 -27
rect 1654 -61 1688 -59
rect 1912 43 1946 45
rect 1912 11 1946 43
rect 1912 -59 1946 -27
rect 1912 -61 1946 -59
rect 2159 43 2193 45
rect 2159 11 2193 43
rect 2159 -59 2193 -27
rect 2159 -61 2193 -59
rect 2417 43 2451 45
rect 2417 11 2451 43
rect 2417 -59 2451 -27
rect 2417 -61 2451 -59
rect 2675 43 2709 45
rect 2675 11 2709 43
rect 2675 -59 2709 -27
rect 2675 -61 2709 -59
rect 2923 43 2957 45
rect 2923 11 2957 43
rect 2923 -59 2957 -27
rect 2923 -61 2957 -59
rect 3181 43 3215 45
rect 3181 11 3215 43
rect 3181 -59 3215 -27
rect 3181 -61 3215 -59
rect 3295 66 3329 90
rect 3295 56 3329 66
rect 3295 -2 3329 18
rect 3295 -16 3329 -2
rect 3295 -70 3329 -54
rect 3295 -88 3329 -70
rect -244 -138 -210 -126
rect -244 -160 -210 -138
rect 3295 -138 3329 -126
rect -37 -180 -35 -146
rect -35 -180 -3 -146
rect 35 -180 67 -146
rect 67 -180 69 -146
rect 468 -180 470 -146
rect 470 -180 502 -146
rect 540 -180 572 -146
rect 572 -180 574 -146
rect 726 -180 728 -146
rect 728 -180 760 -146
rect 798 -180 830 -146
rect 830 -180 832 -146
rect 1231 -180 1233 -146
rect 1233 -180 1265 -146
rect 1303 -180 1335 -146
rect 1335 -180 1337 -146
rect 1489 -180 1491 -146
rect 1491 -180 1523 -146
rect 1561 -180 1593 -146
rect 1593 -180 1595 -146
rect 1747 -180 1749 -146
rect 1749 -180 1781 -146
rect 1819 -180 1851 -146
rect 1851 -180 1853 -146
rect 2252 -180 2254 -146
rect 2254 -180 2286 -146
rect 2324 -180 2356 -146
rect 2356 -180 2358 -146
rect 2510 -180 2512 -146
rect 2512 -180 2544 -146
rect 2582 -180 2614 -146
rect 2614 -180 2616 -146
rect 3016 -180 3018 -146
rect 3018 -180 3050 -146
rect 3088 -180 3120 -146
rect 3120 -180 3122 -146
rect 3295 -160 3329 -138
rect -244 -206 -210 -198
rect -244 -232 -210 -206
rect -244 -274 -210 -270
rect -244 -304 -210 -274
rect -244 -376 -210 -342
rect -244 -444 -210 -414
rect -244 -448 -210 -444
rect -244 -512 -210 -486
rect 3295 -206 3329 -198
rect 3295 -232 3329 -206
rect 3295 -274 3329 -270
rect 3295 -304 3329 -274
rect 3295 -376 3329 -342
rect 3295 -444 3329 -414
rect 3295 -448 3329 -444
rect -244 -520 -210 -512
rect -37 -543 -35 -509
rect -35 -543 -3 -509
rect 35 -543 67 -509
rect 67 -543 69 -509
rect 468 -543 470 -509
rect 470 -543 502 -509
rect 540 -543 572 -509
rect 572 -543 574 -509
rect 726 -543 728 -509
rect 728 -543 760 -509
rect 798 -543 830 -509
rect 830 -543 832 -509
rect 1231 -543 1233 -509
rect 1233 -543 1265 -509
rect 1303 -543 1335 -509
rect 1335 -543 1337 -509
rect 1489 -543 1491 -509
rect 1491 -543 1523 -509
rect 1561 -543 1593 -509
rect 1593 -543 1595 -509
rect 1747 -543 1749 -509
rect 1749 -543 1781 -509
rect 1819 -543 1851 -509
rect 1851 -543 1853 -509
rect 2252 -543 2254 -509
rect 2254 -543 2286 -509
rect 2324 -543 2356 -509
rect 2356 -543 2358 -509
rect 2510 -543 2512 -509
rect 2512 -543 2544 -509
rect 2582 -543 2614 -509
rect 2614 -543 2616 -509
rect 3016 -543 3018 -509
rect 3018 -543 3050 -509
rect 3088 -543 3120 -509
rect 3120 -543 3122 -509
rect 3295 -512 3329 -486
rect 3295 -520 3329 -512
rect -244 -580 -210 -558
rect -244 -592 -210 -580
rect -244 -648 -210 -630
rect -244 -664 -210 -648
rect -244 -716 -210 -702
rect -244 -736 -210 -716
rect -244 -784 -210 -774
rect -244 -808 -210 -784
rect -130 -630 -96 -628
rect -130 -662 -96 -630
rect -130 -732 -96 -700
rect -130 -734 -96 -732
rect 128 -630 162 -628
rect 128 -662 162 -630
rect 128 -732 162 -700
rect 128 -734 162 -732
rect 375 -630 409 -628
rect 375 -662 409 -630
rect 375 -732 409 -700
rect 375 -734 409 -732
rect 633 -630 667 -628
rect 633 -662 667 -630
rect 633 -732 667 -700
rect 633 -734 667 -732
rect 891 -630 925 -628
rect 891 -662 925 -630
rect 891 -732 925 -700
rect 891 -734 925 -732
rect 1138 -630 1172 -628
rect 1138 -662 1172 -630
rect 1138 -732 1172 -700
rect 1138 -734 1172 -732
rect 1396 -630 1430 -628
rect 1396 -662 1430 -630
rect 1396 -732 1430 -700
rect 1396 -734 1430 -732
rect 1654 -630 1688 -628
rect 1654 -662 1688 -630
rect 1654 -732 1688 -700
rect 1654 -734 1688 -732
rect 1912 -630 1946 -628
rect 1912 -662 1946 -630
rect 1912 -732 1946 -700
rect 1912 -734 1946 -732
rect 2159 -630 2193 -628
rect 2159 -662 2193 -630
rect 2159 -732 2193 -700
rect 2159 -734 2193 -732
rect 2417 -630 2451 -628
rect 2417 -662 2451 -630
rect 2417 -732 2451 -700
rect 2417 -734 2451 -732
rect 2675 -630 2709 -628
rect 2675 -662 2709 -630
rect 2675 -732 2709 -700
rect 2675 -734 2709 -732
rect 2923 -630 2957 -628
rect 2923 -662 2957 -630
rect 2923 -732 2957 -700
rect 2923 -734 2957 -732
rect 3181 -630 3215 -628
rect 3181 -662 3215 -630
rect 3181 -732 3215 -700
rect 3181 -734 3215 -732
rect 3295 -580 3329 -558
rect 3295 -592 3329 -580
rect 3295 -648 3329 -630
rect 3295 -664 3329 -648
rect 3295 -716 3329 -702
rect 3295 -736 3329 -716
rect 3295 -784 3329 -774
rect -244 -852 -210 -846
rect -244 -880 -210 -852
rect -244 -952 -210 -918
rect -244 -1024 -210 -990
rect 3295 -808 3329 -784
rect 3295 -852 3329 -846
rect 3295 -880 3329 -852
rect 3295 -952 3329 -918
rect 3295 -1024 3329 -990
rect -244 -1096 -210 -1062
rect -244 -1168 -210 -1134
rect -244 -1234 -210 -1206
rect -244 -1240 -210 -1234
rect -244 -1302 -210 -1278
rect 3295 -1096 3329 -1062
rect 3295 -1168 3329 -1134
rect 3295 -1234 3329 -1206
rect 3295 -1240 3329 -1234
rect -244 -1312 -210 -1302
rect -244 -1370 -210 -1350
rect -244 -1384 -210 -1370
rect -244 -1438 -210 -1422
rect -244 -1456 -210 -1438
rect -244 -1506 -210 -1494
rect -244 -1528 -210 -1506
rect -130 -1354 -96 -1352
rect -130 -1386 -96 -1354
rect -130 -1456 -96 -1424
rect -130 -1458 -96 -1456
rect 128 -1354 162 -1352
rect 128 -1386 162 -1354
rect 128 -1456 162 -1424
rect 128 -1458 162 -1456
rect 375 -1354 409 -1352
rect 375 -1386 409 -1354
rect 375 -1456 409 -1424
rect 375 -1458 409 -1456
rect 633 -1354 667 -1352
rect 633 -1386 667 -1354
rect 633 -1456 667 -1424
rect 633 -1458 667 -1456
rect 891 -1354 925 -1352
rect 891 -1386 925 -1354
rect 891 -1456 925 -1424
rect 891 -1458 925 -1456
rect 1138 -1354 1172 -1352
rect 1138 -1386 1172 -1354
rect 1138 -1456 1172 -1424
rect 1138 -1458 1172 -1456
rect 1396 -1354 1430 -1352
rect 1396 -1386 1430 -1354
rect 1396 -1456 1430 -1424
rect 1396 -1458 1430 -1456
rect 1654 -1354 1688 -1352
rect 1654 -1386 1688 -1354
rect 1654 -1456 1688 -1424
rect 1654 -1458 1688 -1456
rect 1912 -1354 1946 -1352
rect 1912 -1386 1946 -1354
rect 1912 -1456 1946 -1424
rect 1912 -1458 1946 -1456
rect 2159 -1354 2193 -1352
rect 2159 -1386 2193 -1354
rect 2159 -1456 2193 -1424
rect 2159 -1458 2193 -1456
rect 2417 -1354 2451 -1352
rect 2417 -1386 2451 -1354
rect 2417 -1456 2451 -1424
rect 2417 -1458 2451 -1456
rect 2675 -1354 2709 -1352
rect 2675 -1386 2709 -1354
rect 2675 -1456 2709 -1424
rect 2675 -1458 2709 -1456
rect 2923 -1354 2957 -1352
rect 2923 -1386 2957 -1354
rect 2923 -1456 2957 -1424
rect 2923 -1458 2957 -1456
rect 3181 -1354 3215 -1352
rect 3181 -1386 3215 -1354
rect 3181 -1456 3215 -1424
rect 3181 -1458 3215 -1456
rect 3295 -1302 3329 -1278
rect 3295 -1312 3329 -1302
rect 3295 -1370 3329 -1350
rect 3295 -1384 3329 -1370
rect 3295 -1438 3329 -1422
rect 3295 -1456 3329 -1438
rect 3295 -1506 3329 -1494
rect 3295 -1528 3329 -1506
rect -244 -1574 -210 -1566
rect -244 -1600 -210 -1574
rect -37 -1577 -35 -1543
rect -35 -1577 -3 -1543
rect 35 -1577 67 -1543
rect 67 -1577 69 -1543
rect 468 -1577 470 -1543
rect 470 -1577 502 -1543
rect 540 -1577 572 -1543
rect 572 -1577 574 -1543
rect 726 -1577 728 -1543
rect 728 -1577 760 -1543
rect 798 -1577 830 -1543
rect 830 -1577 832 -1543
rect 1231 -1577 1233 -1543
rect 1233 -1577 1265 -1543
rect 1303 -1577 1335 -1543
rect 1335 -1577 1337 -1543
rect 1489 -1577 1491 -1543
rect 1491 -1577 1523 -1543
rect 1561 -1577 1593 -1543
rect 1593 -1577 1595 -1543
rect 1747 -1577 1749 -1543
rect 1749 -1577 1781 -1543
rect 1819 -1577 1851 -1543
rect 1851 -1577 1853 -1543
rect 2252 -1577 2254 -1543
rect 2254 -1577 2286 -1543
rect 2324 -1577 2356 -1543
rect 2356 -1577 2358 -1543
rect 2510 -1577 2512 -1543
rect 2512 -1577 2544 -1543
rect 2582 -1577 2614 -1543
rect 2614 -1577 2616 -1543
rect 3016 -1577 3018 -1543
rect 3018 -1577 3050 -1543
rect 3088 -1577 3120 -1543
rect 3120 -1577 3122 -1543
rect 3295 -1574 3329 -1566
rect -244 -1642 -210 -1638
rect -244 -1672 -210 -1642
rect -244 -1744 -210 -1710
rect -244 -1812 -210 -1782
rect -244 -1816 -210 -1812
rect -244 -1880 -210 -1854
rect -244 -1888 -210 -1880
rect 3295 -1600 3329 -1574
rect 3295 -1642 3329 -1638
rect 3295 -1672 3329 -1642
rect 3295 -1744 3329 -1710
rect 3295 -1812 3329 -1782
rect 3295 -1816 3329 -1812
rect 3295 -1880 3329 -1854
rect 3295 -1888 3329 -1880
rect -244 -1948 -210 -1926
rect -37 -1940 -35 -1906
rect -35 -1940 -3 -1906
rect 35 -1940 67 -1906
rect 67 -1940 69 -1906
rect 468 -1940 470 -1906
rect 470 -1940 502 -1906
rect 540 -1940 572 -1906
rect 572 -1940 574 -1906
rect 726 -1940 728 -1906
rect 728 -1940 760 -1906
rect 798 -1940 830 -1906
rect 830 -1940 832 -1906
rect 1231 -1940 1233 -1906
rect 1233 -1940 1265 -1906
rect 1303 -1940 1335 -1906
rect 1335 -1940 1337 -1906
rect 1489 -1940 1491 -1906
rect 1491 -1940 1523 -1906
rect 1561 -1940 1593 -1906
rect 1593 -1940 1595 -1906
rect 1747 -1940 1749 -1906
rect 1749 -1940 1781 -1906
rect 1819 -1940 1851 -1906
rect 1851 -1940 1853 -1906
rect 2252 -1940 2254 -1906
rect 2254 -1940 2286 -1906
rect 2324 -1940 2356 -1906
rect 2356 -1940 2358 -1906
rect 2510 -1940 2512 -1906
rect 2512 -1940 2544 -1906
rect 2582 -1940 2614 -1906
rect 2614 -1940 2616 -1906
rect 3016 -1940 3018 -1906
rect 3018 -1940 3050 -1906
rect 3088 -1940 3120 -1906
rect 3120 -1940 3122 -1906
rect -244 -1960 -210 -1948
rect 3295 -1948 3329 -1926
rect 3295 -1960 3329 -1948
rect -244 -2016 -210 -1998
rect -244 -2032 -210 -2016
rect -244 -2084 -210 -2070
rect -244 -2104 -210 -2084
rect -244 -2152 -210 -2142
rect -244 -2176 -210 -2152
rect -130 -2027 -96 -2025
rect -130 -2059 -96 -2027
rect -130 -2129 -96 -2097
rect -130 -2131 -96 -2129
rect 128 -2027 162 -2025
rect 128 -2059 162 -2027
rect 128 -2129 162 -2097
rect 128 -2131 162 -2129
rect 375 -2027 409 -2025
rect 375 -2059 409 -2027
rect 375 -2129 409 -2097
rect 375 -2131 409 -2129
rect 633 -2027 667 -2025
rect 633 -2059 667 -2027
rect 633 -2129 667 -2097
rect 633 -2131 667 -2129
rect 891 -2027 925 -2025
rect 891 -2059 925 -2027
rect 891 -2129 925 -2097
rect 891 -2131 925 -2129
rect 1138 -2027 1172 -2025
rect 1138 -2059 1172 -2027
rect 1138 -2129 1172 -2097
rect 1138 -2131 1172 -2129
rect 1396 -2027 1430 -2025
rect 1396 -2059 1430 -2027
rect 1396 -2129 1430 -2097
rect 1396 -2131 1430 -2129
rect 1654 -2027 1688 -2025
rect 1654 -2059 1688 -2027
rect 1654 -2129 1688 -2097
rect 1654 -2131 1688 -2129
rect 1912 -2027 1946 -2025
rect 1912 -2059 1946 -2027
rect 1912 -2129 1946 -2097
rect 1912 -2131 1946 -2129
rect 2159 -2027 2193 -2025
rect 2159 -2059 2193 -2027
rect 2159 -2129 2193 -2097
rect 2159 -2131 2193 -2129
rect 2417 -2027 2451 -2025
rect 2417 -2059 2451 -2027
rect 2417 -2129 2451 -2097
rect 2417 -2131 2451 -2129
rect 2675 -2027 2709 -2025
rect 2675 -2059 2709 -2027
rect 2675 -2129 2709 -2097
rect 2675 -2131 2709 -2129
rect 2923 -2027 2957 -2025
rect 2923 -2059 2957 -2027
rect 2923 -2129 2957 -2097
rect 2923 -2131 2957 -2129
rect 3181 -2027 3215 -2025
rect 3181 -2059 3215 -2027
rect 3181 -2129 3215 -2097
rect 3181 -2131 3215 -2129
rect 3295 -2016 3329 -1998
rect 3295 -2032 3329 -2016
rect 3295 -2084 3329 -2070
rect 3295 -2104 3329 -2084
rect 3295 -2152 3329 -2142
rect 3295 -2176 3329 -2152
rect -244 -2220 -210 -2214
rect -244 -2248 -210 -2220
rect -244 -2288 -210 -2286
rect -244 -2320 -210 -2288
rect -244 -2390 -210 -2358
rect -244 -2392 -210 -2390
rect 3295 -2220 3329 -2214
rect 3295 -2248 3329 -2220
rect 3295 -2288 3329 -2286
rect 3295 -2320 3329 -2288
rect 3295 -2390 3329 -2358
rect 3295 -2392 3329 -2390
rect -244 -2458 -210 -2430
rect 3295 -2458 3329 -2430
rect -244 -2464 -210 -2458
rect -244 -2526 -210 -2502
rect -244 -2536 -210 -2526
rect -244 -2594 -210 -2574
rect -244 -2608 -210 -2594
rect -244 -2662 -210 -2646
rect -244 -2680 -210 -2662
rect 3295 -2464 3329 -2458
rect 3295 -2526 3329 -2502
rect 3295 -2536 3329 -2526
rect 3295 -2594 3329 -2574
rect 3295 -2608 3329 -2594
rect 3295 -2662 3329 -2646
rect 3295 -2680 3329 -2662
rect -244 -2730 -210 -2718
rect -244 -2752 -210 -2730
rect -244 -2798 -210 -2790
rect -244 -2824 -210 -2798
rect -244 -2866 -210 -2862
rect -244 -2896 -210 -2866
rect -130 -2753 -96 -2751
rect -130 -2785 -96 -2753
rect -130 -2855 -96 -2823
rect -130 -2857 -96 -2855
rect 128 -2753 162 -2751
rect 128 -2785 162 -2753
rect 128 -2855 162 -2823
rect 128 -2857 162 -2855
rect 375 -2753 409 -2751
rect 375 -2785 409 -2753
rect 375 -2855 409 -2823
rect 375 -2857 409 -2855
rect 633 -2753 667 -2751
rect 633 -2785 667 -2753
rect 633 -2855 667 -2823
rect 633 -2857 667 -2855
rect 891 -2753 925 -2751
rect 891 -2785 925 -2753
rect 891 -2855 925 -2823
rect 891 -2857 925 -2855
rect 1138 -2753 1172 -2751
rect 1138 -2785 1172 -2753
rect 1138 -2855 1172 -2823
rect 1138 -2857 1172 -2855
rect 1396 -2753 1430 -2751
rect 1396 -2785 1430 -2753
rect 1396 -2855 1430 -2823
rect 1396 -2857 1430 -2855
rect 1654 -2753 1688 -2751
rect 1654 -2785 1688 -2753
rect 1654 -2855 1688 -2823
rect 1654 -2857 1688 -2855
rect 1912 -2753 1946 -2751
rect 1912 -2785 1946 -2753
rect 1912 -2855 1946 -2823
rect 1912 -2857 1946 -2855
rect 2159 -2753 2193 -2751
rect 2159 -2785 2193 -2753
rect 2159 -2855 2193 -2823
rect 2159 -2857 2193 -2855
rect 2417 -2753 2451 -2751
rect 2417 -2785 2451 -2753
rect 2417 -2855 2451 -2823
rect 2417 -2857 2451 -2855
rect 2675 -2753 2709 -2751
rect 2675 -2785 2709 -2753
rect 2675 -2855 2709 -2823
rect 2675 -2857 2709 -2855
rect 2923 -2753 2957 -2751
rect 2923 -2785 2957 -2753
rect 2923 -2855 2957 -2823
rect 2923 -2857 2957 -2855
rect 3181 -2753 3215 -2751
rect 3181 -2785 3215 -2753
rect 3181 -2855 3215 -2823
rect 3181 -2857 3215 -2855
rect 3295 -2730 3329 -2718
rect 3295 -2752 3329 -2730
rect 3295 -2798 3329 -2790
rect 3295 -2824 3329 -2798
rect 3295 -2866 3329 -2862
rect 3295 -2896 3329 -2866
rect -244 -2968 -210 -2934
rect -37 -2976 -35 -2942
rect -35 -2976 -3 -2942
rect 35 -2976 67 -2942
rect 67 -2976 69 -2942
rect 468 -2976 470 -2942
rect 470 -2976 502 -2942
rect 540 -2976 572 -2942
rect 572 -2976 574 -2942
rect 726 -2976 728 -2942
rect 728 -2976 760 -2942
rect 798 -2976 830 -2942
rect 830 -2976 832 -2942
rect 1231 -2976 1233 -2942
rect 1233 -2976 1265 -2942
rect 1303 -2976 1335 -2942
rect 1335 -2976 1337 -2942
rect 1489 -2976 1491 -2942
rect 1491 -2976 1523 -2942
rect 1561 -2976 1593 -2942
rect 1593 -2976 1595 -2942
rect 1747 -2976 1749 -2942
rect 1749 -2976 1781 -2942
rect 1819 -2976 1851 -2942
rect 1851 -2976 1853 -2942
rect 2252 -2976 2254 -2942
rect 2254 -2976 2286 -2942
rect 2324 -2976 2356 -2942
rect 2356 -2976 2358 -2942
rect 2510 -2976 2512 -2942
rect 2512 -2976 2544 -2942
rect 2582 -2976 2614 -2942
rect 2614 -2976 2616 -2942
rect 3016 -2976 3018 -2942
rect 3018 -2976 3050 -2942
rect 3088 -2976 3120 -2942
rect 3120 -2976 3122 -2942
rect 3295 -2968 3329 -2934
rect -80 -3075 -59 -3041
rect -59 -3075 -46 -3041
rect -8 -3075 9 -3041
rect 9 -3075 26 -3041
rect 64 -3075 77 -3041
rect 77 -3075 98 -3041
rect 136 -3075 145 -3041
rect 145 -3075 170 -3041
rect 208 -3075 213 -3041
rect 213 -3075 242 -3041
rect 280 -3075 281 -3041
rect 281 -3075 314 -3041
rect 352 -3075 383 -3041
rect 383 -3075 386 -3041
rect 424 -3075 451 -3041
rect 451 -3075 458 -3041
rect 496 -3075 519 -3041
rect 519 -3075 530 -3041
rect 568 -3075 587 -3041
rect 587 -3075 602 -3041
rect 640 -3075 655 -3041
rect 655 -3075 674 -3041
rect 712 -3075 723 -3041
rect 723 -3075 746 -3041
rect 784 -3075 791 -3041
rect 791 -3075 818 -3041
rect 856 -3075 859 -3041
rect 859 -3075 890 -3041
rect 928 -3075 961 -3041
rect 961 -3075 962 -3041
rect 1000 -3075 1029 -3041
rect 1029 -3075 1034 -3041
rect 1072 -3075 1097 -3041
rect 1097 -3075 1106 -3041
rect 1144 -3075 1165 -3041
rect 1165 -3075 1178 -3041
rect 1216 -3075 1233 -3041
rect 1233 -3075 1250 -3041
rect 1288 -3075 1301 -3041
rect 1301 -3075 1322 -3041
rect 1360 -3075 1369 -3041
rect 1369 -3075 1394 -3041
rect 1432 -3075 1437 -3041
rect 1437 -3075 1466 -3041
rect 1504 -3075 1505 -3041
rect 1505 -3075 1538 -3041
rect 1576 -3075 1607 -3041
rect 1607 -3075 1610 -3041
rect 1648 -3075 1675 -3041
rect 1675 -3075 1682 -3041
rect 1720 -3075 1743 -3041
rect 1743 -3075 1754 -3041
rect 1792 -3075 1811 -3041
rect 1811 -3075 1826 -3041
rect 1864 -3075 1879 -3041
rect 1879 -3075 1898 -3041
rect 1936 -3075 1947 -3041
rect 1947 -3075 1970 -3041
rect 2008 -3075 2015 -3041
rect 2015 -3075 2042 -3041
rect 2080 -3075 2083 -3041
rect 2083 -3075 2114 -3041
rect 2152 -3075 2185 -3041
rect 2185 -3075 2186 -3041
rect 2224 -3075 2253 -3041
rect 2253 -3075 2258 -3041
rect 2296 -3075 2321 -3041
rect 2321 -3075 2330 -3041
rect 2368 -3075 2389 -3041
rect 2389 -3075 2402 -3041
rect 2440 -3075 2457 -3041
rect 2457 -3075 2474 -3041
rect 2512 -3075 2525 -3041
rect 2525 -3075 2546 -3041
rect 2584 -3075 2593 -3041
rect 2593 -3075 2618 -3041
rect 2656 -3075 2661 -3041
rect 2661 -3075 2690 -3041
rect 2728 -3075 2729 -3041
rect 2729 -3075 2762 -3041
rect 2800 -3075 2831 -3041
rect 2831 -3075 2834 -3041
rect 2872 -3075 2899 -3041
rect 2899 -3075 2906 -3041
rect 2944 -3075 2967 -3041
rect 2967 -3075 2978 -3041
rect 3016 -3075 3035 -3041
rect 3035 -3075 3050 -3041
rect 3088 -3075 3103 -3041
rect 3103 -3075 3122 -3041
rect 3160 -3075 3171 -3041
rect 3171 -3075 3194 -3041
<< metal1 >>
rect -269 989 3354 1014
rect -269 955 -80 989
rect -46 955 -8 989
rect 26 955 64 989
rect 98 955 136 989
rect 170 955 208 989
rect 242 955 280 989
rect 314 955 352 989
rect 386 955 424 989
rect 458 955 496 989
rect 530 955 568 989
rect 602 955 640 989
rect 674 955 712 989
rect 746 955 784 989
rect 818 955 856 989
rect 890 955 928 989
rect 962 955 1000 989
rect 1034 955 1072 989
rect 1106 955 1144 989
rect 1178 955 1216 989
rect 1250 955 1288 989
rect 1322 955 1360 989
rect 1394 955 1432 989
rect 1466 955 1504 989
rect 1538 955 1576 989
rect 1610 955 1648 989
rect 1682 955 1720 989
rect 1754 955 1792 989
rect 1826 955 1864 989
rect 1898 955 1936 989
rect 1970 955 2008 989
rect 2042 955 2080 989
rect 2114 955 2152 989
rect 2186 955 2224 989
rect 2258 955 2296 989
rect 2330 955 2368 989
rect 2402 955 2440 989
rect 2474 955 2512 989
rect 2546 955 2584 989
rect 2618 955 2656 989
rect 2690 955 2728 989
rect 2762 955 2800 989
rect 2834 955 2872 989
rect 2906 955 2944 989
rect 2978 955 3016 989
rect 3050 955 3088 989
rect 3122 955 3160 989
rect 3194 955 3354 989
rect -269 890 3354 955
rect -269 882 -37 890
rect -269 848 -244 882
rect -210 856 -37 882
rect -3 856 35 890
rect 69 856 468 890
rect 502 856 540 890
rect 574 856 726 890
rect 760 856 798 890
rect 832 856 1231 890
rect 1265 856 1303 890
rect 1337 856 1489 890
rect 1523 856 1561 890
rect 1595 856 1747 890
rect 1781 856 1819 890
rect 1853 856 2252 890
rect 2286 856 2324 890
rect 2358 856 2510 890
rect 2544 856 2582 890
rect 2616 856 3016 890
rect 3050 856 3088 890
rect 3122 882 3354 890
rect 3122 856 3295 882
rect -210 850 3295 856
rect -210 848 168 850
rect -269 810 168 848
rect -269 776 -244 810
rect -210 776 168 810
rect -269 771 168 776
rect -269 738 -130 771
rect -269 704 -244 738
rect -210 737 -130 738
rect -96 737 128 771
rect 162 737 168 771
rect -210 704 168 737
rect -269 699 168 704
rect -269 666 -130 699
rect -269 632 -244 666
rect -210 665 -130 666
rect -96 665 128 699
rect 162 665 168 699
rect -210 632 168 665
rect -269 594 168 632
rect 369 771 415 850
rect 369 737 375 771
rect 409 737 415 771
rect 369 699 415 737
rect 369 665 375 699
rect 409 665 415 699
rect 369 618 415 665
rect 627 771 673 850
rect 627 737 633 771
rect 667 737 673 771
rect 627 699 673 737
rect 627 665 633 699
rect 667 665 673 699
rect 627 618 673 665
rect 885 771 931 850
rect 885 737 891 771
rect 925 737 931 771
rect 885 699 931 737
rect 885 665 891 699
rect 925 665 931 699
rect 885 618 931 665
rect 1132 771 1178 850
rect 1132 737 1138 771
rect 1172 737 1178 771
rect 1132 699 1178 737
rect 1132 665 1138 699
rect 1172 665 1178 699
rect 1132 618 1178 665
rect 1390 771 1436 850
rect 1390 737 1396 771
rect 1430 737 1436 771
rect 1390 699 1436 737
rect 1390 665 1396 699
rect 1430 665 1436 699
rect 1390 618 1436 665
rect 1648 771 1694 850
rect 1648 737 1654 771
rect 1688 737 1694 771
rect 1648 699 1694 737
rect 1648 665 1654 699
rect 1688 665 1694 699
rect 1648 618 1694 665
rect 1906 771 1952 850
rect 1906 737 1912 771
rect 1946 737 1952 771
rect 1906 699 1952 737
rect 1906 665 1912 699
rect 1946 665 1952 699
rect 1906 618 1952 665
rect 2153 771 2199 850
rect 2153 737 2159 771
rect 2193 737 2199 771
rect 2153 699 2199 737
rect 2153 665 2159 699
rect 2193 665 2199 699
rect 2153 618 2199 665
rect 2411 771 2457 850
rect 2411 737 2417 771
rect 2451 737 2457 771
rect 2411 699 2457 737
rect 2411 665 2417 699
rect 2451 665 2457 699
rect 2411 618 2457 665
rect 2669 771 2715 850
rect 2669 737 2675 771
rect 2709 737 2715 771
rect 2669 699 2715 737
rect 2669 665 2675 699
rect 2709 665 2715 699
rect 2669 618 2715 665
rect 2917 848 3295 850
rect 3329 848 3354 882
rect 2917 810 3354 848
rect 2917 776 3295 810
rect 3329 776 3354 810
rect 2917 771 3354 776
rect 2917 737 2923 771
rect 2957 737 3181 771
rect 3215 738 3354 771
rect 3215 737 3295 738
rect 2917 704 3295 737
rect 3329 704 3354 738
rect 2917 699 3354 704
rect 2917 665 2923 699
rect 2957 665 3181 699
rect 3215 666 3354 699
rect 3215 665 3295 666
rect 2917 632 3295 665
rect 3329 632 3354 666
rect -269 560 -244 594
rect -210 560 168 594
rect -269 522 168 560
rect 2917 594 3354 632
rect 2917 560 3295 594
rect 3329 560 3354 594
rect -269 488 -244 522
rect -210 488 168 522
rect -269 450 168 488
rect 1058 521 1254 529
rect 1058 469 1067 521
rect 1119 469 1131 521
rect 1183 469 1195 521
rect 1247 469 1254 521
rect 1058 459 1254 469
rect 1575 521 1771 529
rect 1575 469 1584 521
rect 1636 469 1648 521
rect 1700 469 1712 521
rect 1764 469 1771 521
rect 1575 459 1771 469
rect 2917 522 3354 560
rect 2917 488 3295 522
rect 3329 488 3354 522
rect -269 416 -244 450
rect -210 416 168 450
rect -269 378 168 416
rect -269 344 -244 378
rect -210 344 168 378
rect -269 306 168 344
rect -269 272 -244 306
rect -210 272 168 306
rect -269 234 168 272
rect -269 200 -244 234
rect -210 200 168 234
rect -269 162 168 200
rect -269 128 -244 162
rect -210 128 168 162
rect -269 90 168 128
rect -269 56 -244 90
rect -210 56 168 90
rect -269 45 168 56
rect -269 18 -130 45
rect -269 -16 -244 18
rect -210 11 -130 18
rect -96 11 128 45
rect 162 11 168 45
rect -210 -16 168 11
rect -269 -27 168 -16
rect -269 -54 -130 -27
rect -269 -88 -244 -54
rect -210 -61 -130 -54
rect -96 -61 128 -27
rect 162 -61 168 -27
rect -210 -88 168 -61
rect -269 -126 168 -88
rect 369 422 931 430
rect 369 370 378 422
rect 430 370 442 422
rect 494 370 506 422
rect 558 370 744 422
rect 796 370 808 422
rect 860 370 872 422
rect 924 370 931 422
rect 369 360 931 370
rect 369 45 415 360
rect 551 211 747 219
rect 551 159 560 211
rect 612 159 624 211
rect 676 159 688 211
rect 740 159 747 211
rect 551 149 747 159
rect 369 11 375 45
rect 409 11 415 45
rect 369 -27 415 11
rect 369 -61 375 -27
rect 409 -61 415 -27
rect 369 -108 415 -61
rect 627 45 673 149
rect 627 11 633 45
rect 667 11 673 45
rect 627 -27 673 11
rect 627 -61 633 -27
rect 667 -61 673 -27
rect 627 -108 673 -61
rect 885 45 931 360
rect 885 11 891 45
rect 925 11 931 45
rect 885 -27 931 11
rect 885 -61 891 -27
rect 925 -61 931 -27
rect 885 -108 931 -61
rect 1132 45 1178 459
rect 1315 310 1511 318
rect 1315 258 1324 310
rect 1376 258 1388 310
rect 1440 258 1452 310
rect 1504 258 1511 310
rect 1315 248 1511 258
rect 1132 11 1138 45
rect 1172 11 1178 45
rect 1132 -27 1178 11
rect 1132 -61 1138 -27
rect 1172 -61 1178 -27
rect 1132 -108 1178 -61
rect 1390 45 1436 248
rect 1390 11 1396 45
rect 1430 11 1436 45
rect 1390 -27 1436 11
rect 1390 -61 1396 -27
rect 1430 -61 1436 -27
rect 1390 -108 1436 -61
rect 1648 45 1694 459
rect 2917 450 3354 488
rect 2153 422 2715 430
rect 2153 370 2162 422
rect 2214 370 2226 422
rect 2278 370 2290 422
rect 2342 370 2528 422
rect 2580 370 2592 422
rect 2644 370 2656 422
rect 2708 370 2715 422
rect 2153 360 2715 370
rect 1832 310 2028 318
rect 1832 258 1841 310
rect 1893 258 1905 310
rect 1957 258 1969 310
rect 2021 258 2028 310
rect 1832 248 2028 258
rect 1648 11 1654 45
rect 1688 11 1694 45
rect 1648 -27 1694 11
rect 1648 -61 1654 -27
rect 1688 -61 1694 -27
rect 1648 -108 1694 -61
rect 1906 45 1952 248
rect 1906 11 1912 45
rect 1946 11 1952 45
rect 1906 -27 1952 11
rect 1906 -61 1912 -27
rect 1946 -61 1952 -27
rect 1906 -108 1952 -61
rect 2153 45 2199 360
rect 2336 211 2532 219
rect 2336 159 2345 211
rect 2397 159 2409 211
rect 2461 159 2473 211
rect 2525 159 2532 211
rect 2336 149 2532 159
rect 2153 11 2159 45
rect 2193 11 2199 45
rect 2153 -27 2199 11
rect 2153 -61 2159 -27
rect 2193 -61 2199 -27
rect 2153 -108 2199 -61
rect 2411 45 2457 149
rect 2411 11 2417 45
rect 2451 11 2457 45
rect 2411 -27 2457 11
rect 2411 -61 2417 -27
rect 2451 -61 2457 -27
rect 2411 -108 2457 -61
rect 2669 45 2715 360
rect 2669 11 2675 45
rect 2709 11 2715 45
rect 2669 -27 2715 11
rect 2669 -61 2675 -27
rect 2709 -61 2715 -27
rect 2669 -108 2715 -61
rect 2917 416 3295 450
rect 3329 416 3354 450
rect 2917 378 3354 416
rect 2917 344 3295 378
rect 3329 344 3354 378
rect 2917 306 3354 344
rect 2917 272 3295 306
rect 3329 272 3354 306
rect 2917 234 3354 272
rect 2917 200 3295 234
rect 3329 200 3354 234
rect 2917 162 3354 200
rect 2917 128 3295 162
rect 3329 128 3354 162
rect 2917 90 3354 128
rect 2917 56 3295 90
rect 3329 56 3354 90
rect 2917 45 3354 56
rect 2917 11 2923 45
rect 2957 11 3181 45
rect 3215 18 3354 45
rect 3215 11 3295 18
rect 2917 -16 3295 11
rect 3329 -16 3354 18
rect 2917 -27 3354 -16
rect 2917 -61 2923 -27
rect 2957 -61 3181 -27
rect 3215 -54 3354 -27
rect 3215 -61 3295 -54
rect 2917 -88 3295 -61
rect 3329 -88 3354 -54
rect -269 -160 -244 -126
rect -210 -146 168 -126
rect 2917 -126 3354 -88
rect -210 -160 -37 -146
rect -269 -180 -37 -160
rect -3 -180 35 -146
rect 69 -180 168 -146
rect -269 -198 168 -180
rect -269 -232 -244 -198
rect -210 -232 168 -198
rect -269 -270 168 -232
rect -269 -304 -244 -270
rect -210 -304 168 -270
rect -269 -342 168 -304
rect -269 -376 -244 -342
rect -210 -376 168 -342
rect -269 -414 168 -376
rect 425 -146 875 -140
rect 425 -180 468 -146
rect 502 -180 540 -146
rect 574 -164 726 -146
rect 425 -216 551 -180
rect 603 -216 615 -164
rect 667 -216 679 -164
rect 760 -180 798 -146
rect 832 -180 875 -146
rect 731 -216 875 -180
rect 425 -315 875 -216
rect 425 -367 551 -315
rect 603 -367 615 -315
rect 667 -367 679 -315
rect 731 -367 875 -315
rect 425 -380 875 -367
rect 964 -146 2121 -140
rect 964 -180 1231 -146
rect 1265 -180 1303 -146
rect 1337 -180 1489 -146
rect 1523 -180 1561 -146
rect 1595 -180 1747 -146
rect 1781 -180 1819 -146
rect 1853 -180 2121 -146
rect 964 -236 2121 -180
rect -269 -448 -244 -414
rect -210 -448 168 -414
rect -269 -486 168 -448
rect 964 -453 1099 -236
rect -269 -520 -244 -486
rect -210 -509 168 -486
rect -210 -520 -37 -509
rect -269 -543 -37 -520
rect -3 -543 35 -509
rect 69 -543 168 -509
rect -269 -558 168 -543
rect 425 -473 1099 -453
rect 425 -509 551 -473
rect 425 -543 468 -509
rect 502 -543 540 -509
rect 603 -525 615 -473
rect 667 -525 679 -473
rect 731 -509 1099 -473
rect 574 -543 726 -525
rect 760 -543 798 -509
rect 832 -543 1099 -509
rect 425 -549 1099 -543
rect 1188 -315 1896 -299
rect 1188 -367 1217 -315
rect 1269 -367 1281 -315
rect 1333 -367 1345 -315
rect 1397 -367 1446 -315
rect 1498 -367 1510 -315
rect 1562 -367 1574 -315
rect 1626 -367 1684 -315
rect 1736 -367 1748 -315
rect 1800 -367 1812 -315
rect 1864 -367 1896 -315
rect 1188 -509 1896 -367
rect 1188 -543 1231 -509
rect 1265 -543 1303 -509
rect 1337 -543 1489 -509
rect 1523 -543 1561 -509
rect 1595 -543 1747 -509
rect 1781 -543 1819 -509
rect 1853 -543 1896 -509
rect 1188 -549 1896 -543
rect 1988 -453 2121 -236
rect 2209 -146 2659 -140
rect 2209 -180 2252 -146
rect 2286 -180 2324 -146
rect 2358 -164 2510 -146
rect 2209 -216 2335 -180
rect 2387 -216 2399 -164
rect 2451 -216 2463 -164
rect 2544 -180 2582 -146
rect 2616 -180 2659 -146
rect 2515 -216 2659 -180
rect 2209 -315 2659 -216
rect 2209 -367 2335 -315
rect 2387 -367 2399 -315
rect 2451 -367 2463 -315
rect 2515 -367 2659 -315
rect 2209 -380 2659 -367
rect 2917 -146 3295 -126
rect 2917 -180 3016 -146
rect 3050 -180 3088 -146
rect 3122 -160 3295 -146
rect 3329 -160 3354 -126
rect 3122 -180 3354 -160
rect 2917 -198 3354 -180
rect 2917 -232 3295 -198
rect 3329 -232 3354 -198
rect 2917 -270 3354 -232
rect 2917 -304 3295 -270
rect 3329 -304 3354 -270
rect 2917 -342 3354 -304
rect 2917 -376 3295 -342
rect 3329 -376 3354 -342
rect 2917 -414 3354 -376
rect 2917 -448 3295 -414
rect 3329 -448 3354 -414
rect 1988 -473 2659 -453
rect 1988 -509 2335 -473
rect 1988 -543 2252 -509
rect 2286 -543 2324 -509
rect 2387 -525 2399 -473
rect 2451 -525 2463 -473
rect 2515 -509 2659 -473
rect 2358 -543 2510 -525
rect 2544 -543 2582 -509
rect 2616 -543 2659 -509
rect 1988 -549 2659 -543
rect 2917 -486 3354 -448
rect 2917 -509 3295 -486
rect 2917 -543 3016 -509
rect 3050 -543 3088 -509
rect 3122 -520 3295 -509
rect 3329 -520 3354 -486
rect 3122 -543 3354 -520
rect -269 -592 -244 -558
rect -210 -592 168 -558
rect 2917 -558 3354 -543
rect -269 -628 168 -592
rect -269 -630 -130 -628
rect -269 -664 -244 -630
rect -210 -662 -130 -630
rect -96 -662 128 -628
rect 162 -662 168 -628
rect -210 -664 168 -662
rect -269 -700 168 -664
rect -269 -702 -130 -700
rect -269 -736 -244 -702
rect -210 -734 -130 -702
rect -96 -734 128 -700
rect 162 -734 168 -700
rect -210 -736 168 -734
rect -269 -774 168 -736
rect -269 -808 -244 -774
rect -210 -808 168 -774
rect -269 -846 168 -808
rect -269 -880 -244 -846
rect -210 -880 168 -846
rect -269 -918 168 -880
rect -269 -952 -244 -918
rect -210 -952 168 -918
rect -269 -990 168 -952
rect -269 -1024 -244 -990
rect -210 -1024 168 -990
rect -269 -1062 168 -1024
rect -269 -1096 -244 -1062
rect -210 -1096 168 -1062
rect 369 -628 415 -581
rect 369 -662 375 -628
rect 409 -662 415 -628
rect 369 -700 415 -662
rect 369 -734 375 -700
rect 409 -734 415 -700
rect 369 -1063 415 -734
rect 627 -628 673 -581
rect 627 -662 633 -628
rect 667 -662 673 -628
rect 627 -700 673 -662
rect 627 -734 633 -700
rect 667 -734 673 -700
rect 627 -853 673 -734
rect 885 -628 931 -581
rect 885 -662 891 -628
rect 925 -662 931 -628
rect 885 -700 931 -662
rect 885 -734 891 -700
rect 925 -734 931 -700
rect 553 -863 749 -853
rect 553 -915 560 -863
rect 612 -915 624 -863
rect 676 -915 688 -863
rect 740 -915 749 -863
rect 553 -923 749 -915
rect -269 -1134 168 -1096
rect 294 -1073 490 -1063
rect 294 -1125 301 -1073
rect 353 -1125 365 -1073
rect 417 -1125 429 -1073
rect 481 -1125 490 -1073
rect 294 -1133 490 -1125
rect -269 -1168 -244 -1134
rect -210 -1168 168 -1134
rect -269 -1206 168 -1168
rect -269 -1240 -244 -1206
rect -210 -1240 168 -1206
rect -269 -1278 168 -1240
rect -269 -1312 -244 -1278
rect -210 -1312 168 -1278
rect -269 -1350 168 -1312
rect -269 -1384 -244 -1350
rect -210 -1352 168 -1350
rect -210 -1384 -130 -1352
rect -269 -1386 -130 -1384
rect -96 -1386 128 -1352
rect 162 -1386 168 -1352
rect -269 -1422 168 -1386
rect -269 -1456 -244 -1422
rect -210 -1424 168 -1422
rect -210 -1456 -130 -1424
rect -269 -1458 -130 -1456
rect -96 -1458 128 -1424
rect 162 -1458 168 -1424
rect -269 -1494 168 -1458
rect -269 -1528 -244 -1494
rect -210 -1528 168 -1494
rect 369 -1352 415 -1133
rect 369 -1386 375 -1352
rect 409 -1386 415 -1352
rect 369 -1424 415 -1386
rect 369 -1458 375 -1424
rect 409 -1458 415 -1424
rect 369 -1505 415 -1458
rect 627 -1352 673 -923
rect 885 -1063 931 -734
rect 1132 -628 1178 -581
rect 1132 -662 1138 -628
rect 1172 -662 1178 -628
rect 1132 -700 1178 -662
rect 1132 -734 1138 -700
rect 1172 -734 1178 -700
rect 1132 -952 1178 -734
rect 1390 -628 1436 -581
rect 1390 -662 1396 -628
rect 1430 -662 1436 -628
rect 1390 -700 1436 -662
rect 1390 -734 1396 -700
rect 1430 -734 1436 -700
rect 1057 -962 1253 -952
rect 1057 -1014 1064 -962
rect 1116 -1014 1128 -962
rect 1180 -1014 1192 -962
rect 1244 -1014 1253 -962
rect 1057 -1022 1253 -1014
rect 813 -1073 1009 -1063
rect 813 -1125 820 -1073
rect 872 -1125 884 -1073
rect 936 -1125 948 -1073
rect 1000 -1125 1009 -1073
rect 813 -1133 1009 -1125
rect 627 -1386 633 -1352
rect 667 -1386 673 -1352
rect 627 -1424 673 -1386
rect 627 -1458 633 -1424
rect 667 -1458 673 -1424
rect 627 -1505 673 -1458
rect 885 -1352 931 -1133
rect 885 -1386 891 -1352
rect 925 -1386 931 -1352
rect 885 -1424 931 -1386
rect 885 -1458 891 -1424
rect 925 -1458 931 -1424
rect 885 -1505 931 -1458
rect 1132 -1352 1178 -1022
rect 1390 -1163 1436 -734
rect 1648 -628 1694 -581
rect 1648 -662 1654 -628
rect 1688 -662 1694 -628
rect 1648 -700 1694 -662
rect 1648 -734 1654 -700
rect 1688 -734 1694 -700
rect 1648 -952 1694 -734
rect 1906 -628 1952 -581
rect 1906 -662 1912 -628
rect 1946 -662 1952 -628
rect 1906 -700 1952 -662
rect 1906 -734 1912 -700
rect 1946 -734 1952 -700
rect 1574 -962 1770 -952
rect 1574 -1014 1581 -962
rect 1633 -1014 1645 -962
rect 1697 -1014 1709 -962
rect 1761 -1014 1770 -962
rect 1574 -1022 1770 -1014
rect 1314 -1173 1510 -1163
rect 1314 -1225 1321 -1173
rect 1373 -1225 1385 -1173
rect 1437 -1225 1449 -1173
rect 1501 -1225 1510 -1173
rect 1314 -1233 1510 -1225
rect 1132 -1386 1138 -1352
rect 1172 -1386 1178 -1352
rect 1132 -1424 1178 -1386
rect 1132 -1458 1138 -1424
rect 1172 -1458 1178 -1424
rect 1132 -1505 1178 -1458
rect 1390 -1352 1436 -1233
rect 1390 -1386 1396 -1352
rect 1430 -1386 1436 -1352
rect 1390 -1424 1436 -1386
rect 1390 -1458 1396 -1424
rect 1430 -1458 1436 -1424
rect 1390 -1505 1436 -1458
rect 1648 -1352 1694 -1022
rect 1906 -1163 1952 -734
rect 2153 -628 2199 -581
rect 2153 -662 2159 -628
rect 2193 -662 2199 -628
rect 2153 -700 2199 -662
rect 2153 -734 2159 -700
rect 2193 -734 2199 -700
rect 2153 -1063 2199 -734
rect 2411 -628 2457 -581
rect 2411 -662 2417 -628
rect 2451 -662 2457 -628
rect 2411 -700 2457 -662
rect 2411 -734 2417 -700
rect 2451 -734 2457 -700
rect 2411 -853 2457 -734
rect 2669 -628 2715 -581
rect 2669 -662 2675 -628
rect 2709 -662 2715 -628
rect 2669 -700 2715 -662
rect 2669 -734 2675 -700
rect 2709 -734 2715 -700
rect 2337 -863 2533 -853
rect 2337 -915 2344 -863
rect 2396 -915 2408 -863
rect 2460 -915 2472 -863
rect 2524 -915 2533 -863
rect 2337 -923 2533 -915
rect 2080 -1073 2276 -1063
rect 2080 -1125 2087 -1073
rect 2139 -1125 2151 -1073
rect 2203 -1125 2215 -1073
rect 2267 -1125 2276 -1073
rect 2080 -1133 2276 -1125
rect 1831 -1173 2027 -1163
rect 1831 -1225 1838 -1173
rect 1890 -1225 1902 -1173
rect 1954 -1225 1966 -1173
rect 2018 -1225 2027 -1173
rect 1831 -1233 2027 -1225
rect 1648 -1386 1654 -1352
rect 1688 -1386 1694 -1352
rect 1648 -1424 1694 -1386
rect 1648 -1458 1654 -1424
rect 1688 -1458 1694 -1424
rect 1648 -1505 1694 -1458
rect 1906 -1352 1952 -1233
rect 1906 -1386 1912 -1352
rect 1946 -1386 1952 -1352
rect 1906 -1424 1952 -1386
rect 1906 -1458 1912 -1424
rect 1946 -1458 1952 -1424
rect 1906 -1505 1952 -1458
rect 2153 -1352 2199 -1133
rect 2153 -1386 2159 -1352
rect 2193 -1386 2199 -1352
rect 2153 -1424 2199 -1386
rect 2153 -1458 2159 -1424
rect 2193 -1458 2199 -1424
rect 2153 -1505 2199 -1458
rect 2411 -1352 2457 -923
rect 2669 -1063 2715 -734
rect 2917 -592 3295 -558
rect 3329 -592 3354 -558
rect 2917 -628 3354 -592
rect 2917 -662 2923 -628
rect 2957 -662 3181 -628
rect 3215 -630 3354 -628
rect 3215 -662 3295 -630
rect 2917 -664 3295 -662
rect 3329 -664 3354 -630
rect 2917 -700 3354 -664
rect 2917 -734 2923 -700
rect 2957 -734 3181 -700
rect 3215 -702 3354 -700
rect 3215 -734 3295 -702
rect 2917 -736 3295 -734
rect 3329 -736 3354 -702
rect 2917 -774 3354 -736
rect 2917 -808 3295 -774
rect 3329 -808 3354 -774
rect 2917 -846 3354 -808
rect 2917 -880 3295 -846
rect 3329 -880 3354 -846
rect 2917 -918 3354 -880
rect 2917 -952 3295 -918
rect 3329 -952 3354 -918
rect 2917 -990 3354 -952
rect 2917 -1024 3295 -990
rect 3329 -1024 3354 -990
rect 2917 -1062 3354 -1024
rect 2597 -1073 2793 -1063
rect 2597 -1125 2604 -1073
rect 2656 -1125 2668 -1073
rect 2720 -1125 2732 -1073
rect 2784 -1125 2793 -1073
rect 2597 -1133 2793 -1125
rect 2917 -1096 3295 -1062
rect 3329 -1096 3354 -1062
rect 2411 -1386 2417 -1352
rect 2451 -1386 2457 -1352
rect 2411 -1424 2457 -1386
rect 2411 -1458 2417 -1424
rect 2451 -1458 2457 -1424
rect 2411 -1505 2457 -1458
rect 2669 -1352 2715 -1133
rect 2669 -1386 2675 -1352
rect 2709 -1386 2715 -1352
rect 2669 -1424 2715 -1386
rect 2669 -1458 2675 -1424
rect 2709 -1458 2715 -1424
rect 2669 -1505 2715 -1458
rect 2917 -1134 3354 -1096
rect 2917 -1168 3295 -1134
rect 3329 -1168 3354 -1134
rect 2917 -1206 3354 -1168
rect 2917 -1240 3295 -1206
rect 3329 -1240 3354 -1206
rect 2917 -1278 3354 -1240
rect 2917 -1312 3295 -1278
rect 3329 -1312 3354 -1278
rect 2917 -1350 3354 -1312
rect 2917 -1352 3295 -1350
rect 2917 -1386 2923 -1352
rect 2957 -1386 3181 -1352
rect 3215 -1384 3295 -1352
rect 3329 -1384 3354 -1350
rect 3215 -1386 3354 -1384
rect 2917 -1422 3354 -1386
rect 2917 -1424 3295 -1422
rect 2917 -1458 2923 -1424
rect 2957 -1458 3181 -1424
rect 3215 -1456 3295 -1424
rect 3329 -1456 3354 -1422
rect 3215 -1458 3354 -1456
rect 2917 -1494 3354 -1458
rect -269 -1543 168 -1528
rect 2917 -1528 3295 -1494
rect 3329 -1528 3354 -1494
rect -269 -1566 -37 -1543
rect -269 -1600 -244 -1566
rect -210 -1577 -37 -1566
rect -3 -1577 35 -1543
rect 69 -1577 168 -1543
rect -210 -1600 168 -1577
rect -269 -1638 168 -1600
rect 425 -1543 1099 -1537
rect 425 -1577 468 -1543
rect 502 -1577 540 -1543
rect 574 -1561 726 -1543
rect 425 -1613 551 -1577
rect 603 -1613 615 -1561
rect 667 -1613 679 -1561
rect 760 -1577 798 -1543
rect 832 -1577 1099 -1543
rect 731 -1613 1099 -1577
rect 425 -1633 1099 -1613
rect -269 -1672 -244 -1638
rect -210 -1672 168 -1638
rect -269 -1710 168 -1672
rect -269 -1744 -244 -1710
rect -210 -1744 168 -1710
rect -269 -1782 168 -1744
rect -269 -1816 -244 -1782
rect -210 -1816 168 -1782
rect -269 -1854 168 -1816
rect -269 -1888 -244 -1854
rect -210 -1888 168 -1854
rect -269 -1906 168 -1888
rect -269 -1926 -37 -1906
rect -269 -1960 -244 -1926
rect -210 -1940 -37 -1926
rect -3 -1940 35 -1906
rect 69 -1940 168 -1906
rect -210 -1960 168 -1940
rect 425 -1718 875 -1706
rect 425 -1770 551 -1718
rect 603 -1770 615 -1718
rect 667 -1770 679 -1718
rect 731 -1770 875 -1718
rect 425 -1870 875 -1770
rect 425 -1906 551 -1870
rect 425 -1940 468 -1906
rect 502 -1940 540 -1906
rect 603 -1922 615 -1870
rect 667 -1922 679 -1870
rect 731 -1906 875 -1870
rect 574 -1940 726 -1922
rect 760 -1940 798 -1906
rect 832 -1940 875 -1906
rect 425 -1946 875 -1940
rect 964 -1850 1099 -1633
rect 1188 -1543 1896 -1537
rect 1188 -1577 1231 -1543
rect 1265 -1577 1303 -1543
rect 1337 -1577 1489 -1543
rect 1523 -1577 1561 -1543
rect 1595 -1577 1747 -1543
rect 1781 -1577 1819 -1543
rect 1853 -1577 1896 -1543
rect 1188 -1718 1896 -1577
rect 1188 -1770 1217 -1718
rect 1269 -1770 1281 -1718
rect 1333 -1770 1345 -1718
rect 1397 -1770 1446 -1718
rect 1498 -1770 1510 -1718
rect 1562 -1770 1574 -1718
rect 1626 -1770 1684 -1718
rect 1736 -1770 1748 -1718
rect 1800 -1770 1812 -1718
rect 1864 -1770 1896 -1718
rect 1188 -1787 1896 -1770
rect 1988 -1543 2659 -1537
rect 1988 -1577 2252 -1543
rect 2286 -1577 2324 -1543
rect 2358 -1561 2510 -1543
rect 1988 -1613 2335 -1577
rect 2387 -1613 2399 -1561
rect 2451 -1613 2463 -1561
rect 2544 -1577 2582 -1543
rect 2616 -1577 2659 -1543
rect 2515 -1613 2659 -1577
rect 1988 -1633 2659 -1613
rect 2917 -1543 3354 -1528
rect 2917 -1577 3016 -1543
rect 3050 -1577 3088 -1543
rect 3122 -1566 3354 -1543
rect 3122 -1577 3295 -1566
rect 2917 -1600 3295 -1577
rect 3329 -1600 3354 -1566
rect 1988 -1850 2121 -1633
rect 2917 -1638 3354 -1600
rect 2917 -1672 3295 -1638
rect 3329 -1672 3354 -1638
rect 964 -1906 2121 -1850
rect 964 -1940 1231 -1906
rect 1265 -1940 1303 -1906
rect 1337 -1940 1489 -1906
rect 1523 -1940 1561 -1906
rect 1595 -1940 1747 -1906
rect 1781 -1940 1819 -1906
rect 1853 -1940 2121 -1906
rect 964 -1946 2121 -1940
rect 2209 -1718 2659 -1706
rect 2209 -1770 2335 -1718
rect 2387 -1770 2399 -1718
rect 2451 -1770 2463 -1718
rect 2515 -1770 2659 -1718
rect 2209 -1870 2659 -1770
rect 2209 -1906 2335 -1870
rect 2209 -1940 2252 -1906
rect 2286 -1940 2324 -1906
rect 2387 -1922 2399 -1870
rect 2451 -1922 2463 -1870
rect 2515 -1906 2659 -1870
rect 2358 -1940 2510 -1922
rect 2544 -1940 2582 -1906
rect 2616 -1940 2659 -1906
rect 2209 -1946 2659 -1940
rect 2917 -1710 3354 -1672
rect 2917 -1744 3295 -1710
rect 3329 -1744 3354 -1710
rect 2917 -1782 3354 -1744
rect 2917 -1816 3295 -1782
rect 3329 -1816 3354 -1782
rect 2917 -1854 3354 -1816
rect 2917 -1888 3295 -1854
rect 3329 -1888 3354 -1854
rect 2917 -1906 3354 -1888
rect 2917 -1940 3016 -1906
rect 3050 -1940 3088 -1906
rect 3122 -1926 3354 -1906
rect 3122 -1940 3295 -1926
rect -269 -1998 168 -1960
rect 2917 -1960 3295 -1940
rect 3329 -1960 3354 -1926
rect -269 -2032 -244 -1998
rect -210 -2025 168 -1998
rect -210 -2032 -130 -2025
rect -269 -2059 -130 -2032
rect -96 -2059 128 -2025
rect 162 -2059 168 -2025
rect -269 -2070 168 -2059
rect -269 -2104 -244 -2070
rect -210 -2097 168 -2070
rect -210 -2104 -130 -2097
rect -269 -2131 -130 -2104
rect -96 -2131 128 -2097
rect 162 -2131 168 -2097
rect -269 -2142 168 -2131
rect -269 -2176 -244 -2142
rect -210 -2176 168 -2142
rect -269 -2214 168 -2176
rect -269 -2248 -244 -2214
rect -210 -2248 168 -2214
rect -269 -2286 168 -2248
rect -269 -2320 -244 -2286
rect -210 -2320 168 -2286
rect -269 -2358 168 -2320
rect -269 -2392 -244 -2358
rect -210 -2392 168 -2358
rect -269 -2430 168 -2392
rect -269 -2464 -244 -2430
rect -210 -2464 168 -2430
rect -269 -2502 168 -2464
rect -269 -2536 -244 -2502
rect -210 -2536 168 -2502
rect 369 -2025 415 -1978
rect 369 -2059 375 -2025
rect 409 -2059 415 -2025
rect 369 -2097 415 -2059
rect 369 -2131 375 -2097
rect 409 -2131 415 -2097
rect 369 -2446 415 -2131
rect 627 -2025 673 -1978
rect 627 -2059 633 -2025
rect 667 -2059 673 -2025
rect 627 -2097 673 -2059
rect 627 -2131 633 -2097
rect 667 -2131 673 -2097
rect 627 -2235 673 -2131
rect 885 -2025 931 -1978
rect 885 -2059 891 -2025
rect 925 -2059 931 -2025
rect 885 -2097 931 -2059
rect 885 -2131 891 -2097
rect 925 -2131 931 -2097
rect 553 -2245 749 -2235
rect 553 -2297 560 -2245
rect 612 -2297 624 -2245
rect 676 -2297 688 -2245
rect 740 -2297 749 -2245
rect 553 -2305 749 -2297
rect 885 -2446 931 -2131
rect 1132 -2025 1178 -1978
rect 1132 -2059 1138 -2025
rect 1172 -2059 1178 -2025
rect 1132 -2097 1178 -2059
rect 1132 -2131 1138 -2097
rect 1172 -2131 1178 -2097
rect 1132 -2334 1178 -2131
rect 1390 -2025 1436 -1978
rect 1390 -2059 1396 -2025
rect 1430 -2059 1436 -2025
rect 1390 -2097 1436 -2059
rect 1390 -2131 1396 -2097
rect 1430 -2131 1436 -2097
rect 1057 -2344 1253 -2334
rect 1057 -2396 1064 -2344
rect 1116 -2396 1128 -2344
rect 1180 -2396 1192 -2344
rect 1244 -2396 1253 -2344
rect 1057 -2404 1253 -2396
rect 369 -2456 931 -2446
rect 369 -2508 376 -2456
rect 428 -2508 440 -2456
rect 492 -2508 504 -2456
rect 556 -2508 742 -2456
rect 794 -2508 806 -2456
rect 858 -2508 870 -2456
rect 922 -2508 931 -2456
rect 369 -2516 931 -2508
rect -269 -2574 168 -2536
rect 1390 -2545 1436 -2131
rect 1648 -2025 1694 -1978
rect 1648 -2059 1654 -2025
rect 1688 -2059 1694 -2025
rect 1648 -2097 1694 -2059
rect 1648 -2131 1654 -2097
rect 1688 -2131 1694 -2097
rect 1648 -2334 1694 -2131
rect 1906 -2025 1952 -1978
rect 1906 -2059 1912 -2025
rect 1946 -2059 1952 -2025
rect 1906 -2097 1952 -2059
rect 1906 -2131 1912 -2097
rect 1946 -2131 1952 -2097
rect 1574 -2344 1770 -2334
rect 1574 -2396 1581 -2344
rect 1633 -2396 1645 -2344
rect 1697 -2396 1709 -2344
rect 1761 -2396 1770 -2344
rect 1574 -2404 1770 -2396
rect 1906 -2545 1952 -2131
rect 2153 -2025 2199 -1978
rect 2153 -2059 2159 -2025
rect 2193 -2059 2199 -2025
rect 2153 -2097 2199 -2059
rect 2153 -2131 2159 -2097
rect 2193 -2131 2199 -2097
rect 2153 -2446 2199 -2131
rect 2411 -2025 2457 -1978
rect 2411 -2059 2417 -2025
rect 2451 -2059 2457 -2025
rect 2411 -2097 2457 -2059
rect 2411 -2131 2417 -2097
rect 2451 -2131 2457 -2097
rect 2411 -2235 2457 -2131
rect 2669 -2025 2715 -1978
rect 2669 -2059 2675 -2025
rect 2709 -2059 2715 -2025
rect 2669 -2097 2715 -2059
rect 2669 -2131 2675 -2097
rect 2709 -2131 2715 -2097
rect 2337 -2245 2533 -2235
rect 2337 -2297 2344 -2245
rect 2396 -2297 2408 -2245
rect 2460 -2297 2472 -2245
rect 2524 -2297 2533 -2245
rect 2337 -2305 2533 -2297
rect 2669 -2446 2715 -2131
rect 2153 -2456 2715 -2446
rect 2153 -2508 2160 -2456
rect 2212 -2508 2224 -2456
rect 2276 -2508 2288 -2456
rect 2340 -2508 2526 -2456
rect 2578 -2508 2590 -2456
rect 2642 -2508 2654 -2456
rect 2706 -2508 2715 -2456
rect 2153 -2516 2715 -2508
rect 2917 -1998 3354 -1960
rect 2917 -2025 3295 -1998
rect 2917 -2059 2923 -2025
rect 2957 -2059 3181 -2025
rect 3215 -2032 3295 -2025
rect 3329 -2032 3354 -1998
rect 3215 -2059 3354 -2032
rect 2917 -2070 3354 -2059
rect 2917 -2097 3295 -2070
rect 2917 -2131 2923 -2097
rect 2957 -2131 3181 -2097
rect 3215 -2104 3295 -2097
rect 3329 -2104 3354 -2070
rect 3215 -2131 3354 -2104
rect 2917 -2142 3354 -2131
rect 2917 -2176 3295 -2142
rect 3329 -2176 3354 -2142
rect 2917 -2214 3354 -2176
rect 2917 -2248 3295 -2214
rect 3329 -2248 3354 -2214
rect 2917 -2286 3354 -2248
rect 2917 -2320 3295 -2286
rect 3329 -2320 3354 -2286
rect 2917 -2358 3354 -2320
rect 2917 -2392 3295 -2358
rect 3329 -2392 3354 -2358
rect 2917 -2430 3354 -2392
rect 2917 -2464 3295 -2430
rect 3329 -2464 3354 -2430
rect 2917 -2502 3354 -2464
rect 2917 -2536 3295 -2502
rect 3329 -2536 3354 -2502
rect -269 -2608 -244 -2574
rect -210 -2608 168 -2574
rect -269 -2646 168 -2608
rect 1314 -2555 1510 -2545
rect 1314 -2607 1321 -2555
rect 1373 -2607 1385 -2555
rect 1437 -2607 1449 -2555
rect 1501 -2607 1510 -2555
rect 1314 -2615 1510 -2607
rect 1831 -2555 2027 -2545
rect 1831 -2607 1838 -2555
rect 1890 -2607 1902 -2555
rect 1954 -2607 1966 -2555
rect 2018 -2607 2027 -2555
rect 1831 -2615 2027 -2607
rect 2917 -2574 3354 -2536
rect 2917 -2608 3295 -2574
rect 3329 -2608 3354 -2574
rect -269 -2680 -244 -2646
rect -210 -2680 168 -2646
rect -269 -2718 168 -2680
rect 2917 -2646 3354 -2608
rect 2917 -2680 3295 -2646
rect 3329 -2680 3354 -2646
rect -269 -2752 -244 -2718
rect -210 -2751 168 -2718
rect -210 -2752 -130 -2751
rect -269 -2785 -130 -2752
rect -96 -2785 128 -2751
rect 162 -2785 168 -2751
rect -269 -2790 168 -2785
rect -269 -2824 -244 -2790
rect -210 -2823 168 -2790
rect -210 -2824 -130 -2823
rect -269 -2857 -130 -2824
rect -96 -2857 128 -2823
rect 162 -2857 168 -2823
rect -269 -2862 168 -2857
rect -269 -2896 -244 -2862
rect -210 -2896 168 -2862
rect -269 -2934 168 -2896
rect -269 -2968 -244 -2934
rect -210 -2936 168 -2934
rect 369 -2751 415 -2704
rect 369 -2785 375 -2751
rect 409 -2785 415 -2751
rect 369 -2823 415 -2785
rect 369 -2857 375 -2823
rect 409 -2857 415 -2823
rect 369 -2936 415 -2857
rect 627 -2751 673 -2704
rect 627 -2785 633 -2751
rect 667 -2785 673 -2751
rect 627 -2823 673 -2785
rect 627 -2857 633 -2823
rect 667 -2857 673 -2823
rect 627 -2936 673 -2857
rect 885 -2751 931 -2704
rect 885 -2785 891 -2751
rect 925 -2785 931 -2751
rect 885 -2823 931 -2785
rect 885 -2857 891 -2823
rect 925 -2857 931 -2823
rect 885 -2936 931 -2857
rect 1132 -2751 1178 -2704
rect 1132 -2785 1138 -2751
rect 1172 -2785 1178 -2751
rect 1132 -2823 1178 -2785
rect 1132 -2857 1138 -2823
rect 1172 -2857 1178 -2823
rect 1132 -2936 1178 -2857
rect 1390 -2751 1436 -2704
rect 1390 -2785 1396 -2751
rect 1430 -2785 1436 -2751
rect 1390 -2823 1436 -2785
rect 1390 -2857 1396 -2823
rect 1430 -2857 1436 -2823
rect 1390 -2936 1436 -2857
rect 1648 -2751 1694 -2704
rect 1648 -2785 1654 -2751
rect 1688 -2785 1694 -2751
rect 1648 -2823 1694 -2785
rect 1648 -2857 1654 -2823
rect 1688 -2857 1694 -2823
rect 1648 -2936 1694 -2857
rect 1906 -2751 1952 -2704
rect 1906 -2785 1912 -2751
rect 1946 -2785 1952 -2751
rect 1906 -2823 1952 -2785
rect 1906 -2857 1912 -2823
rect 1946 -2857 1952 -2823
rect 1906 -2936 1952 -2857
rect 2153 -2751 2199 -2704
rect 2153 -2785 2159 -2751
rect 2193 -2785 2199 -2751
rect 2153 -2823 2199 -2785
rect 2153 -2857 2159 -2823
rect 2193 -2857 2199 -2823
rect 2153 -2936 2199 -2857
rect 2411 -2751 2457 -2704
rect 2411 -2785 2417 -2751
rect 2451 -2785 2457 -2751
rect 2411 -2823 2457 -2785
rect 2411 -2857 2417 -2823
rect 2451 -2857 2457 -2823
rect 2411 -2936 2457 -2857
rect 2669 -2751 2715 -2704
rect 2669 -2785 2675 -2751
rect 2709 -2785 2715 -2751
rect 2669 -2823 2715 -2785
rect 2669 -2857 2675 -2823
rect 2709 -2857 2715 -2823
rect 2669 -2936 2715 -2857
rect 2917 -2718 3354 -2680
rect 2917 -2751 3295 -2718
rect 2917 -2785 2923 -2751
rect 2957 -2785 3181 -2751
rect 3215 -2752 3295 -2751
rect 3329 -2752 3354 -2718
rect 3215 -2785 3354 -2752
rect 2917 -2790 3354 -2785
rect 2917 -2823 3295 -2790
rect 2917 -2857 2923 -2823
rect 2957 -2857 3181 -2823
rect 3215 -2824 3295 -2823
rect 3329 -2824 3354 -2790
rect 3215 -2857 3354 -2824
rect 2917 -2862 3354 -2857
rect 2917 -2896 3295 -2862
rect 3329 -2896 3354 -2862
rect 2917 -2934 3354 -2896
rect 2917 -2936 3295 -2934
rect -210 -2942 3295 -2936
rect -210 -2968 -37 -2942
rect -269 -2976 -37 -2968
rect -3 -2976 35 -2942
rect 69 -2976 468 -2942
rect 502 -2976 540 -2942
rect 574 -2976 726 -2942
rect 760 -2976 798 -2942
rect 832 -2976 1231 -2942
rect 1265 -2976 1303 -2942
rect 1337 -2976 1489 -2942
rect 1523 -2976 1561 -2942
rect 1595 -2976 1747 -2942
rect 1781 -2976 1819 -2942
rect 1853 -2976 2252 -2942
rect 2286 -2976 2324 -2942
rect 2358 -2976 2510 -2942
rect 2544 -2976 2582 -2942
rect 2616 -2976 3016 -2942
rect 3050 -2976 3088 -2942
rect 3122 -2968 3295 -2942
rect 3329 -2968 3354 -2934
rect 3122 -2976 3354 -2968
rect -269 -3041 3354 -2976
rect -269 -3075 -80 -3041
rect -46 -3075 -8 -3041
rect 26 -3075 64 -3041
rect 98 -3075 136 -3041
rect 170 -3075 208 -3041
rect 242 -3075 280 -3041
rect 314 -3075 352 -3041
rect 386 -3075 424 -3041
rect 458 -3075 496 -3041
rect 530 -3075 568 -3041
rect 602 -3075 640 -3041
rect 674 -3075 712 -3041
rect 746 -3075 784 -3041
rect 818 -3075 856 -3041
rect 890 -3075 928 -3041
rect 962 -3075 1000 -3041
rect 1034 -3075 1072 -3041
rect 1106 -3075 1144 -3041
rect 1178 -3075 1216 -3041
rect 1250 -3075 1288 -3041
rect 1322 -3075 1360 -3041
rect 1394 -3075 1432 -3041
rect 1466 -3075 1504 -3041
rect 1538 -3075 1576 -3041
rect 1610 -3075 1648 -3041
rect 1682 -3075 1720 -3041
rect 1754 -3075 1792 -3041
rect 1826 -3075 1864 -3041
rect 1898 -3075 1936 -3041
rect 1970 -3075 2008 -3041
rect 2042 -3075 2080 -3041
rect 2114 -3075 2152 -3041
rect 2186 -3075 2224 -3041
rect 2258 -3075 2296 -3041
rect 2330 -3075 2368 -3041
rect 2402 -3075 2440 -3041
rect 2474 -3075 2512 -3041
rect 2546 -3075 2584 -3041
rect 2618 -3075 2656 -3041
rect 2690 -3075 2728 -3041
rect 2762 -3075 2800 -3041
rect 2834 -3075 2872 -3041
rect 2906 -3075 2944 -3041
rect 2978 -3075 3016 -3041
rect 3050 -3075 3088 -3041
rect 3122 -3075 3160 -3041
rect 3194 -3075 3354 -3041
rect -269 -3100 3354 -3075
<< via1 >>
rect 1067 469 1119 521
rect 1131 469 1183 521
rect 1195 469 1247 521
rect 1584 469 1636 521
rect 1648 469 1700 521
rect 1712 469 1764 521
rect 378 370 430 422
rect 442 370 494 422
rect 506 370 558 422
rect 744 370 796 422
rect 808 370 860 422
rect 872 370 924 422
rect 560 159 612 211
rect 624 159 676 211
rect 688 159 740 211
rect 1324 258 1376 310
rect 1388 258 1440 310
rect 1452 258 1504 310
rect 2162 370 2214 422
rect 2226 370 2278 422
rect 2290 370 2342 422
rect 2528 370 2580 422
rect 2592 370 2644 422
rect 2656 370 2708 422
rect 1841 258 1893 310
rect 1905 258 1957 310
rect 1969 258 2021 310
rect 2345 159 2397 211
rect 2409 159 2461 211
rect 2473 159 2525 211
rect 551 -180 574 -164
rect 574 -180 603 -164
rect 551 -216 603 -180
rect 615 -216 667 -164
rect 679 -180 726 -164
rect 726 -180 731 -164
rect 679 -216 731 -180
rect 551 -367 603 -315
rect 615 -367 667 -315
rect 679 -367 731 -315
rect 551 -509 603 -473
rect 551 -525 574 -509
rect 574 -525 603 -509
rect 615 -525 667 -473
rect 679 -509 731 -473
rect 679 -525 726 -509
rect 726 -525 731 -509
rect 1217 -367 1269 -315
rect 1281 -367 1333 -315
rect 1345 -367 1397 -315
rect 1446 -367 1498 -315
rect 1510 -367 1562 -315
rect 1574 -367 1626 -315
rect 1684 -367 1736 -315
rect 1748 -367 1800 -315
rect 1812 -367 1864 -315
rect 2335 -180 2358 -164
rect 2358 -180 2387 -164
rect 2335 -216 2387 -180
rect 2399 -216 2451 -164
rect 2463 -180 2510 -164
rect 2510 -180 2515 -164
rect 2463 -216 2515 -180
rect 2335 -367 2387 -315
rect 2399 -367 2451 -315
rect 2463 -367 2515 -315
rect 2335 -509 2387 -473
rect 2335 -525 2358 -509
rect 2358 -525 2387 -509
rect 2399 -525 2451 -473
rect 2463 -509 2515 -473
rect 2463 -525 2510 -509
rect 2510 -525 2515 -509
rect 560 -915 612 -863
rect 624 -915 676 -863
rect 688 -915 740 -863
rect 301 -1125 353 -1073
rect 365 -1125 417 -1073
rect 429 -1125 481 -1073
rect 1064 -1014 1116 -962
rect 1128 -1014 1180 -962
rect 1192 -1014 1244 -962
rect 820 -1125 872 -1073
rect 884 -1125 936 -1073
rect 948 -1125 1000 -1073
rect 1581 -1014 1633 -962
rect 1645 -1014 1697 -962
rect 1709 -1014 1761 -962
rect 1321 -1225 1373 -1173
rect 1385 -1225 1437 -1173
rect 1449 -1225 1501 -1173
rect 2344 -915 2396 -863
rect 2408 -915 2460 -863
rect 2472 -915 2524 -863
rect 2087 -1125 2139 -1073
rect 2151 -1125 2203 -1073
rect 2215 -1125 2267 -1073
rect 1838 -1225 1890 -1173
rect 1902 -1225 1954 -1173
rect 1966 -1225 2018 -1173
rect 2604 -1125 2656 -1073
rect 2668 -1125 2720 -1073
rect 2732 -1125 2784 -1073
rect 551 -1577 574 -1561
rect 574 -1577 603 -1561
rect 551 -1613 603 -1577
rect 615 -1613 667 -1561
rect 679 -1577 726 -1561
rect 726 -1577 731 -1561
rect 679 -1613 731 -1577
rect 551 -1770 603 -1718
rect 615 -1770 667 -1718
rect 679 -1770 731 -1718
rect 551 -1906 603 -1870
rect 551 -1922 574 -1906
rect 574 -1922 603 -1906
rect 615 -1922 667 -1870
rect 679 -1906 731 -1870
rect 679 -1922 726 -1906
rect 726 -1922 731 -1906
rect 1217 -1770 1269 -1718
rect 1281 -1770 1333 -1718
rect 1345 -1770 1397 -1718
rect 1446 -1770 1498 -1718
rect 1510 -1770 1562 -1718
rect 1574 -1770 1626 -1718
rect 1684 -1770 1736 -1718
rect 1748 -1770 1800 -1718
rect 1812 -1770 1864 -1718
rect 2335 -1577 2358 -1561
rect 2358 -1577 2387 -1561
rect 2335 -1613 2387 -1577
rect 2399 -1613 2451 -1561
rect 2463 -1577 2510 -1561
rect 2510 -1577 2515 -1561
rect 2463 -1613 2515 -1577
rect 2335 -1770 2387 -1718
rect 2399 -1770 2451 -1718
rect 2463 -1770 2515 -1718
rect 2335 -1906 2387 -1870
rect 2335 -1922 2358 -1906
rect 2358 -1922 2387 -1906
rect 2399 -1922 2451 -1870
rect 2463 -1906 2515 -1870
rect 2463 -1922 2510 -1906
rect 2510 -1922 2515 -1906
rect 560 -2297 612 -2245
rect 624 -2297 676 -2245
rect 688 -2297 740 -2245
rect 1064 -2396 1116 -2344
rect 1128 -2396 1180 -2344
rect 1192 -2396 1244 -2344
rect 376 -2508 428 -2456
rect 440 -2508 492 -2456
rect 504 -2508 556 -2456
rect 742 -2508 794 -2456
rect 806 -2508 858 -2456
rect 870 -2508 922 -2456
rect 1581 -2396 1633 -2344
rect 1645 -2396 1697 -2344
rect 1709 -2396 1761 -2344
rect 2344 -2297 2396 -2245
rect 2408 -2297 2460 -2245
rect 2472 -2297 2524 -2245
rect 2160 -2508 2212 -2456
rect 2224 -2508 2276 -2456
rect 2288 -2508 2340 -2456
rect 2526 -2508 2578 -2456
rect 2590 -2508 2642 -2456
rect 2654 -2508 2706 -2456
rect 1321 -2607 1373 -2555
rect 1385 -2607 1437 -2555
rect 1449 -2607 1501 -2555
rect 1838 -2607 1890 -2555
rect 1902 -2607 1954 -2555
rect 1966 -2607 2018 -2555
<< metal2 >>
rect -269 521 1861 529
rect -269 507 1067 521
rect -269 451 -229 507
rect -173 451 -149 507
rect -93 451 -69 507
rect -13 469 1067 507
rect 1119 469 1131 521
rect 1183 469 1195 521
rect 1247 469 1584 521
rect 1636 469 1648 521
rect 1700 469 1712 521
rect 1764 469 1861 521
rect -13 459 1861 469
rect -13 451 31 459
rect -269 429 31 451
rect 369 422 3354 430
rect 369 370 378 422
rect 430 370 442 422
rect 494 370 506 422
rect 558 370 744 422
rect 796 370 808 422
rect 860 370 872 422
rect 924 370 2162 422
rect 2214 370 2226 422
rect 2278 370 2290 422
rect 2342 370 2528 422
rect 2580 370 2592 422
rect 2644 370 2656 422
rect 2708 408 3354 422
rect 2708 370 3094 408
rect 369 360 3094 370
rect 3054 352 3094 360
rect 3150 352 3174 408
rect 3230 352 3254 408
rect 3310 352 3354 408
rect 3054 330 3354 352
rect 163 310 2028 318
rect 163 296 1324 310
rect 163 240 203 296
rect 259 240 283 296
rect 339 240 363 296
rect 419 258 1324 296
rect 1376 258 1388 310
rect 1440 258 1452 310
rect 1504 258 1841 310
rect 1893 258 1905 310
rect 1957 258 1969 310
rect 2021 258 2028 310
rect 419 248 2028 258
rect 419 240 463 248
rect 163 218 463 240
rect 551 211 2922 219
rect 551 159 560 211
rect 612 159 624 211
rect 676 159 688 211
rect 740 159 2345 211
rect 2397 159 2409 211
rect 2461 159 2473 211
rect 2525 197 2922 211
rect 2525 159 2662 197
rect 551 149 2662 159
rect 2622 141 2662 149
rect 2718 141 2742 197
rect 2798 141 2822 197
rect 2878 141 2922 197
rect 2622 119 2922 141
rect 1906 -140 2206 -136
rect 425 -158 2662 -140
rect 425 -164 1946 -158
rect 425 -216 551 -164
rect 603 -216 615 -164
rect 667 -216 679 -164
rect 731 -214 1946 -164
rect 2002 -214 2026 -158
rect 2082 -214 2106 -158
rect 2162 -164 2662 -158
rect 2162 -214 2335 -164
rect 731 -216 2335 -214
rect 2387 -216 2399 -164
rect 2451 -216 2463 -164
rect 2515 -216 2662 -164
rect 425 -236 2662 -216
rect 425 -315 2662 -299
rect 425 -367 551 -315
rect 603 -367 615 -315
rect 667 -367 679 -315
rect 731 -367 1217 -315
rect 1269 -367 1281 -315
rect 1333 -367 1345 -315
rect 1397 -367 1446 -315
rect 1498 -367 1510 -315
rect 1562 -367 1574 -315
rect 1626 -367 1684 -315
rect 1736 -367 1748 -315
rect 1800 -367 1812 -315
rect 1864 -321 2335 -315
rect 1864 -367 1946 -321
rect 425 -377 1946 -367
rect 2002 -377 2026 -321
rect 2082 -377 2106 -321
rect 2162 -367 2335 -321
rect 2387 -367 2399 -315
rect 2451 -367 2463 -315
rect 2515 -367 2662 -315
rect 2162 -377 2662 -367
rect 425 -380 2662 -377
rect 1906 -399 2206 -380
rect 425 -473 2662 -453
rect 425 -525 551 -473
rect 603 -525 615 -473
rect 667 -525 679 -473
rect 731 -475 2335 -473
rect 731 -525 919 -475
rect 425 -531 919 -525
rect 975 -531 999 -475
rect 1055 -531 1079 -475
rect 1135 -525 2335 -475
rect 2387 -525 2399 -473
rect 2451 -525 2463 -473
rect 2515 -525 2662 -473
rect 1135 -531 2662 -525
rect 425 -549 2662 -531
rect 879 -553 1179 -549
rect 163 -845 463 -823
rect 163 -901 203 -845
rect 259 -901 283 -845
rect 339 -901 363 -845
rect 419 -853 463 -845
rect 419 -863 2533 -853
rect 419 -901 560 -863
rect 163 -915 560 -901
rect 612 -915 624 -863
rect 676 -915 688 -863
rect 740 -915 2344 -863
rect 2396 -915 2408 -863
rect 2460 -915 2472 -863
rect 2524 -915 2533 -863
rect 163 -923 2533 -915
rect 2622 -944 2922 -922
rect 2622 -952 2662 -944
rect 1057 -962 2662 -952
rect 1057 -1014 1064 -962
rect 1116 -1014 1128 -962
rect 1180 -1014 1192 -962
rect 1244 -1014 1581 -962
rect 1633 -1014 1645 -962
rect 1697 -1014 1709 -962
rect 1761 -1000 2662 -962
rect 2718 -1000 2742 -944
rect 2798 -1000 2822 -944
rect 2878 -1000 2922 -944
rect 1761 -1014 2922 -1000
rect 1057 -1022 2922 -1014
rect -269 -1055 31 -1033
rect -269 -1111 -229 -1055
rect -173 -1111 -149 -1055
rect -93 -1111 -69 -1055
rect -13 -1063 31 -1055
rect -13 -1073 2793 -1063
rect -13 -1111 301 -1073
rect -269 -1125 301 -1111
rect 353 -1125 365 -1073
rect 417 -1125 429 -1073
rect 481 -1125 820 -1073
rect 872 -1125 884 -1073
rect 936 -1125 948 -1073
rect 1000 -1125 2087 -1073
rect 2139 -1125 2151 -1073
rect 2203 -1125 2215 -1073
rect 2267 -1125 2604 -1073
rect 2656 -1125 2668 -1073
rect 2720 -1125 2732 -1073
rect 2784 -1125 2793 -1073
rect -269 -1133 2793 -1125
rect 1314 -1173 3354 -1163
rect 1314 -1225 1321 -1173
rect 1373 -1225 1385 -1173
rect 1437 -1225 1449 -1173
rect 1501 -1225 1838 -1173
rect 1890 -1225 1902 -1173
rect 1954 -1225 1966 -1173
rect 2018 -1185 3354 -1173
rect 2018 -1225 3094 -1185
rect 1314 -1233 3094 -1225
rect 3054 -1241 3094 -1233
rect 3150 -1241 3174 -1185
rect 3230 -1241 3254 -1185
rect 3310 -1241 3354 -1185
rect 3054 -1263 3354 -1241
rect 879 -1537 1179 -1533
rect 425 -1555 2662 -1537
rect 425 -1561 919 -1555
rect 425 -1613 551 -1561
rect 603 -1613 615 -1561
rect 667 -1613 679 -1561
rect 731 -1611 919 -1561
rect 975 -1611 999 -1555
rect 1055 -1611 1079 -1555
rect 1135 -1561 2662 -1555
rect 1135 -1611 2335 -1561
rect 731 -1613 2335 -1611
rect 2387 -1613 2399 -1561
rect 2451 -1613 2463 -1561
rect 2515 -1613 2662 -1561
rect 425 -1633 2662 -1613
rect 1906 -1706 2206 -1687
rect 425 -1709 2662 -1706
rect 425 -1718 1946 -1709
rect 425 -1770 551 -1718
rect 603 -1770 615 -1718
rect 667 -1770 679 -1718
rect 731 -1770 1217 -1718
rect 1269 -1770 1281 -1718
rect 1333 -1770 1345 -1718
rect 1397 -1770 1446 -1718
rect 1498 -1770 1510 -1718
rect 1562 -1770 1574 -1718
rect 1626 -1770 1684 -1718
rect 1736 -1770 1748 -1718
rect 1800 -1770 1812 -1718
rect 1864 -1765 1946 -1718
rect 2002 -1765 2026 -1709
rect 2082 -1765 2106 -1709
rect 2162 -1718 2662 -1709
rect 2162 -1765 2335 -1718
rect 1864 -1770 2335 -1765
rect 2387 -1770 2399 -1718
rect 2451 -1770 2463 -1718
rect 2515 -1770 2662 -1718
rect 425 -1787 2662 -1770
rect 425 -1870 2662 -1850
rect 425 -1922 551 -1870
rect 603 -1922 615 -1870
rect 667 -1922 679 -1870
rect 731 -1872 2335 -1870
rect 731 -1922 1946 -1872
rect 425 -1928 1946 -1922
rect 2002 -1928 2026 -1872
rect 2082 -1928 2106 -1872
rect 2162 -1922 2335 -1872
rect 2387 -1922 2399 -1870
rect 2451 -1922 2463 -1870
rect 2515 -1922 2662 -1870
rect 2162 -1928 2662 -1922
rect 425 -1946 2662 -1928
rect 1906 -1950 2206 -1946
rect 2622 -2227 2922 -2205
rect 2622 -2235 2662 -2227
rect 550 -2245 2662 -2235
rect 550 -2297 560 -2245
rect 612 -2297 624 -2245
rect 676 -2297 688 -2245
rect 740 -2297 2344 -2245
rect 2396 -2297 2408 -2245
rect 2460 -2297 2472 -2245
rect 2524 -2283 2662 -2245
rect 2718 -2283 2742 -2227
rect 2798 -2283 2822 -2227
rect 2878 -2283 2922 -2227
rect 2524 -2297 2922 -2283
rect 550 -2305 2922 -2297
rect 163 -2327 463 -2305
rect 163 -2383 203 -2327
rect 259 -2383 283 -2327
rect 339 -2383 363 -2327
rect 419 -2334 463 -2327
rect 419 -2344 1770 -2334
rect 419 -2383 1064 -2344
rect 163 -2396 1064 -2383
rect 1116 -2396 1128 -2344
rect 1180 -2396 1192 -2344
rect 1244 -2396 1581 -2344
rect 1633 -2396 1645 -2344
rect 1697 -2396 1709 -2344
rect 1761 -2396 1770 -2344
rect 163 -2405 1770 -2396
rect 3054 -2438 3354 -2416
rect 3054 -2446 3094 -2438
rect 369 -2456 3094 -2446
rect 369 -2508 376 -2456
rect 428 -2508 440 -2456
rect 492 -2508 504 -2456
rect 556 -2508 742 -2456
rect 794 -2508 806 -2456
rect 858 -2508 870 -2456
rect 922 -2508 2160 -2456
rect 2212 -2508 2224 -2456
rect 2276 -2508 2288 -2456
rect 2340 -2508 2526 -2456
rect 2578 -2508 2590 -2456
rect 2642 -2508 2654 -2456
rect 2706 -2494 3094 -2456
rect 3150 -2494 3174 -2438
rect 3230 -2494 3254 -2438
rect 3310 -2494 3354 -2438
rect 2706 -2508 3354 -2494
rect -269 -2537 31 -2515
rect 369 -2516 3354 -2508
rect -269 -2593 -229 -2537
rect -173 -2593 -149 -2537
rect -93 -2593 -69 -2537
rect -13 -2545 31 -2537
rect -13 -2555 2027 -2545
rect -13 -2593 1321 -2555
rect -269 -2607 1321 -2593
rect 1373 -2607 1385 -2555
rect 1437 -2607 1449 -2555
rect 1501 -2607 1838 -2555
rect 1890 -2607 1902 -2555
rect 1954 -2607 1966 -2555
rect 2018 -2607 2027 -2555
rect -269 -2615 2027 -2607
<< via2 >>
rect -229 451 -173 507
rect -149 451 -93 507
rect -69 451 -13 507
rect 3094 352 3150 408
rect 3174 352 3230 408
rect 3254 352 3310 408
rect 203 240 259 296
rect 283 240 339 296
rect 363 240 419 296
rect 2662 141 2718 197
rect 2742 141 2798 197
rect 2822 141 2878 197
rect 1946 -214 2002 -158
rect 2026 -214 2082 -158
rect 2106 -214 2162 -158
rect 1946 -377 2002 -321
rect 2026 -377 2082 -321
rect 2106 -377 2162 -321
rect 919 -531 975 -475
rect 999 -531 1055 -475
rect 1079 -531 1135 -475
rect 203 -901 259 -845
rect 283 -901 339 -845
rect 363 -901 419 -845
rect 2662 -1000 2718 -944
rect 2742 -1000 2798 -944
rect 2822 -1000 2878 -944
rect -229 -1111 -173 -1055
rect -149 -1111 -93 -1055
rect -69 -1111 -13 -1055
rect 3094 -1241 3150 -1185
rect 3174 -1241 3230 -1185
rect 3254 -1241 3310 -1185
rect 919 -1611 975 -1555
rect 999 -1611 1055 -1555
rect 1079 -1611 1135 -1555
rect 1946 -1765 2002 -1709
rect 2026 -1765 2082 -1709
rect 2106 -1765 2162 -1709
rect 1946 -1928 2002 -1872
rect 2026 -1928 2082 -1872
rect 2106 -1928 2162 -1872
rect 2662 -2283 2718 -2227
rect 2742 -2283 2798 -2227
rect 2822 -2283 2878 -2227
rect 203 -2383 259 -2327
rect 283 -2383 339 -2327
rect 363 -2383 419 -2327
rect 3094 -2494 3150 -2438
rect 3174 -2494 3230 -2438
rect 3254 -2494 3310 -2438
rect -229 -2593 -173 -2537
rect -149 -2593 -93 -2537
rect -69 -2593 -13 -2537
<< metal3 >>
rect -269 507 31 529
rect -269 451 -229 507
rect -173 451 -149 507
rect -93 451 -69 507
rect -13 451 31 507
rect -269 -1055 31 451
rect 3054 408 3354 430
rect 3054 352 3094 408
rect 3150 352 3174 408
rect 3230 352 3254 408
rect 3310 352 3354 408
rect -269 -1111 -229 -1055
rect -173 -1111 -149 -1055
rect -93 -1111 -69 -1055
rect -13 -1111 31 -1055
rect -269 -2537 31 -1111
rect 163 296 463 318
rect 163 240 203 296
rect 259 240 283 296
rect 339 240 363 296
rect 419 240 463 296
rect 163 -845 463 240
rect 2622 197 2922 219
rect 2622 141 2662 197
rect 2718 141 2742 197
rect 2798 141 2822 197
rect 2878 141 2922 197
rect 1906 -158 2206 -136
rect 1906 -214 1946 -158
rect 2002 -214 2026 -158
rect 2082 -214 2106 -158
rect 2162 -214 2206 -158
rect 1906 -321 2206 -214
rect 1906 -377 1946 -321
rect 2002 -377 2026 -321
rect 2082 -377 2106 -321
rect 2162 -377 2206 -321
rect 163 -901 203 -845
rect 259 -901 283 -845
rect 339 -901 363 -845
rect 419 -901 463 -845
rect 163 -2327 463 -901
rect 879 -475 1180 -453
rect 879 -531 919 -475
rect 975 -531 999 -475
rect 1055 -531 1079 -475
rect 1135 -531 1180 -475
rect 879 -1555 1180 -531
rect 879 -1611 919 -1555
rect 975 -1611 999 -1555
rect 1055 -1611 1079 -1555
rect 1135 -1611 1180 -1555
rect 879 -1633 1180 -1611
rect 1906 -1709 2206 -377
rect 1906 -1765 1946 -1709
rect 2002 -1765 2026 -1709
rect 2082 -1765 2106 -1709
rect 2162 -1765 2206 -1709
rect 1906 -1872 2206 -1765
rect 1906 -1928 1946 -1872
rect 2002 -1928 2026 -1872
rect 2082 -1928 2106 -1872
rect 2162 -1928 2206 -1872
rect 1906 -1950 2206 -1928
rect 2622 -944 2922 141
rect 2622 -1000 2662 -944
rect 2718 -1000 2742 -944
rect 2798 -1000 2822 -944
rect 2878 -1000 2922 -944
rect 2622 -2227 2922 -1000
rect 2622 -2283 2662 -2227
rect 2718 -2283 2742 -2227
rect 2798 -2283 2822 -2227
rect 2878 -2283 2922 -2227
rect 2622 -2305 2922 -2283
rect 3054 -1185 3354 352
rect 3054 -1241 3094 -1185
rect 3150 -1241 3174 -1185
rect 3230 -1241 3254 -1185
rect 3310 -1241 3354 -1185
rect 163 -2383 203 -2327
rect 259 -2383 283 -2327
rect 339 -2383 363 -2327
rect 419 -2383 463 -2327
rect 163 -2405 463 -2383
rect 3054 -2438 3354 -1241
rect 3054 -2494 3094 -2438
rect 3150 -2494 3174 -2438
rect 3230 -2494 3254 -2438
rect 3310 -2494 3354 -2438
rect 3054 -2516 3354 -2494
rect -269 -2593 -229 -2537
rect -173 -2593 -149 -2537
rect -93 -2593 -69 -2537
rect -13 -2593 31 -2537
rect -269 -2615 31 -2593
<< end >>
