magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< metal1 >>
rect -25399 11832 17024 11904
rect -25399 11810 -24568 11832
rect -7560 11810 -3505 11832
rect 4759 11810 8311 11832
rect 16824 11810 17024 11832
rect -25399 11483 17024 11810
rect -25399 11243 -24568 11483
rect -20686 11404 -20490 11412
rect -20686 11352 -20679 11404
rect -20627 11352 -20615 11404
rect -20563 11352 -20551 11404
rect -20499 11352 -20490 11404
rect -20686 11342 -20490 11352
rect -20364 11404 -20168 11412
rect -20364 11352 -20357 11404
rect -20305 11352 -20293 11404
rect -20241 11352 -20229 11404
rect -20177 11352 -20168 11404
rect -20364 11342 -20168 11352
rect -11979 11404 -11783 11412
rect -11979 11352 -11972 11404
rect -11920 11352 -11908 11404
rect -11856 11352 -11844 11404
rect -11792 11352 -11783 11404
rect -11979 11342 -11783 11352
rect -11640 11404 -11444 11412
rect -11640 11352 -11633 11404
rect -11581 11352 -11569 11404
rect -11517 11352 -11505 11404
rect -11453 11352 -11444 11404
rect -11640 11342 -11444 11352
rect -7560 11243 -3505 11483
rect 403 11404 599 11412
rect 403 11352 410 11404
rect 462 11352 474 11404
rect 526 11352 538 11404
rect 590 11352 599 11404
rect 403 11342 599 11352
rect 755 11404 951 11412
rect 755 11352 762 11404
rect 814 11352 826 11404
rect 878 11352 890 11404
rect 942 11352 951 11404
rect 755 11342 951 11352
rect 4759 11243 8311 11483
rect -25399 11235 -24560 11243
rect -25399 11183 -24747 11235
rect -24695 11183 -24683 11235
rect -24631 11183 -24619 11235
rect -24567 11183 -24560 11235
rect -25399 11173 -24560 11183
rect -16380 11235 -16184 11243
rect -16380 11183 -16371 11235
rect -16319 11183 -16307 11235
rect -16255 11183 -16243 11235
rect -16191 11183 -16184 11235
rect -16380 11173 -16184 11183
rect -15977 11235 -15781 11243
rect -15977 11183 -15968 11235
rect -15916 11183 -15904 11235
rect -15852 11183 -15840 11235
rect -15788 11183 -15781 11235
rect -15977 11173 -15781 11183
rect -7686 11235 -3401 11243
rect -7686 11183 -7677 11235
rect -7625 11183 -7613 11235
rect -7561 11183 -7549 11235
rect -7497 11183 -3588 11235
rect -3536 11183 -3524 11235
rect -3472 11183 -3460 11235
rect -3408 11183 -3401 11235
rect -7686 11173 -3401 11183
rect 4746 11235 8311 11243
rect 4746 11183 4755 11235
rect 4807 11183 4819 11235
rect 4871 11183 4883 11235
rect 4935 11183 8311 11235
rect 16824 11234 17024 11483
rect 4746 11173 8311 11183
rect 16861 11182 16873 11234
rect 16925 11182 17024 11234
rect -25399 9276 -24568 11173
rect -20685 9714 -20489 9722
rect -20685 9662 -20678 9714
rect -20626 9662 -20614 9714
rect -20562 9662 -20550 9714
rect -20498 9662 -20489 9714
rect -20685 9652 -20489 9662
rect -20363 9714 -20167 9722
rect -20363 9662 -20356 9714
rect -20304 9662 -20292 9714
rect -20240 9662 -20228 9714
rect -20176 9662 -20167 9714
rect -20363 9652 -20167 9662
rect -11978 9714 -11782 9722
rect -11978 9662 -11971 9714
rect -11919 9662 -11907 9714
rect -11855 9662 -11843 9714
rect -11791 9662 -11782 9714
rect -11978 9652 -11782 9662
rect -11640 9714 -11444 9722
rect -11640 9662 -11633 9714
rect -11581 9662 -11569 9714
rect -11517 9662 -11505 9714
rect -11453 9662 -11444 9714
rect -11640 9652 -11444 9662
rect -7560 9276 -3505 11173
rect 404 9714 600 9722
rect 404 9662 411 9714
rect 463 9662 475 9714
rect 527 9662 539 9714
rect 591 9662 600 9714
rect 404 9652 600 9662
rect 756 9714 952 9722
rect 756 9662 763 9714
rect 815 9662 827 9714
rect 879 9662 891 9714
rect 943 9662 952 9714
rect 756 9652 952 9662
rect 4759 9276 8311 11173
rect -25399 9268 -24558 9276
rect -25399 9216 -24745 9268
rect -24693 9216 -24681 9268
rect -24629 9216 -24617 9268
rect -24565 9216 -24558 9268
rect -25399 9206 -24558 9216
rect -16379 9268 -16183 9276
rect -16379 9216 -16370 9268
rect -16318 9216 -16306 9268
rect -16254 9216 -16242 9268
rect -16190 9216 -16183 9268
rect -16379 9206 -16183 9216
rect -15976 9268 -15780 9276
rect -15976 9216 -15967 9268
rect -15915 9216 -15903 9268
rect -15851 9216 -15839 9268
rect -15787 9216 -15780 9268
rect -15976 9206 -15780 9216
rect -7684 9268 -3399 9276
rect -7684 9216 -7675 9268
rect -7623 9216 -7611 9268
rect -7559 9216 -7547 9268
rect -7495 9216 -3586 9268
rect -3534 9216 -3522 9268
rect -3470 9216 -3458 9268
rect -3406 9216 -3399 9268
rect -7684 9206 -3399 9216
rect 4748 9268 8311 9276
rect 16824 9268 17024 11182
rect 4748 9216 4757 9268
rect 4809 9216 4821 9268
rect 4873 9216 4885 9268
rect 4937 9216 8311 9268
rect 16847 9216 16859 9268
rect 16911 9216 17024 9268
rect 4748 9206 8311 9216
rect -25399 7768 -24568 9206
rect -7560 7768 -3505 9206
rect 4759 7768 8311 9206
rect -25399 7758 -24562 7768
rect -25399 7706 -24749 7758
rect -24697 7706 -24685 7758
rect -24633 7706 -24621 7758
rect -24569 7706 -24562 7758
rect -25399 7698 -24562 7706
rect -16383 7758 -16187 7768
rect -16383 7706 -16374 7758
rect -16322 7706 -16310 7758
rect -16258 7706 -16246 7758
rect -16194 7706 -16187 7758
rect -16383 7698 -16187 7706
rect -15980 7758 -15784 7768
rect -15980 7706 -15971 7758
rect -15919 7706 -15907 7758
rect -15855 7706 -15843 7758
rect -15791 7706 -15784 7758
rect -15980 7698 -15784 7706
rect -7688 7758 -3403 7768
rect -7688 7706 -7679 7758
rect -7627 7706 -7615 7758
rect -7563 7706 -7551 7758
rect -7499 7706 -3590 7758
rect -3538 7706 -3526 7758
rect -3474 7706 -3462 7758
rect -3410 7706 -3403 7758
rect -7688 7698 -3403 7706
rect 4744 7758 8311 7768
rect 16824 7758 17024 9216
rect 4744 7706 4753 7758
rect 4805 7706 4817 7758
rect 4869 7706 4881 7758
rect 4933 7706 8311 7758
rect 16850 7706 16862 7758
rect 16914 7706 17024 7758
rect 4744 7698 8311 7706
rect -25399 6370 -24568 7698
rect -20709 7590 -20513 7600
rect -20709 7538 -20702 7590
rect -20650 7538 -20638 7590
rect -20586 7538 -20574 7590
rect -20522 7538 -20513 7590
rect -20709 7530 -20513 7538
rect -20387 7590 -20191 7600
rect -20387 7538 -20380 7590
rect -20328 7538 -20316 7590
rect -20264 7538 -20252 7590
rect -20200 7538 -20191 7590
rect -20387 7530 -20191 7538
rect -12002 7590 -11806 7600
rect -12002 7538 -11995 7590
rect -11943 7538 -11931 7590
rect -11879 7538 -11867 7590
rect -11815 7538 -11806 7590
rect -12002 7530 -11806 7538
rect -11663 7590 -11467 7600
rect -11663 7538 -11656 7590
rect -11604 7538 -11592 7590
rect -11540 7538 -11528 7590
rect -11476 7538 -11467 7590
rect -11663 7530 -11467 7538
rect -20688 6530 -20492 6538
rect -20688 6478 -20681 6530
rect -20629 6478 -20617 6530
rect -20565 6478 -20553 6530
rect -20501 6478 -20492 6530
rect -20688 6468 -20492 6478
rect -20367 6530 -20171 6538
rect -20367 6478 -20360 6530
rect -20308 6478 -20296 6530
rect -20244 6478 -20232 6530
rect -20180 6478 -20171 6530
rect -20367 6468 -20171 6478
rect -11981 6530 -11785 6538
rect -11981 6478 -11974 6530
rect -11922 6478 -11910 6530
rect -11858 6478 -11846 6530
rect -11794 6478 -11785 6530
rect -11981 6468 -11785 6478
rect -11643 6530 -11447 6538
rect -11643 6478 -11636 6530
rect -11584 6478 -11572 6530
rect -11520 6478 -11508 6530
rect -11456 6478 -11447 6530
rect -11643 6468 -11447 6478
rect -7560 6370 -3505 7698
rect 380 7590 576 7600
rect 380 7538 387 7590
rect 439 7538 451 7590
rect 503 7538 515 7590
rect 567 7538 576 7590
rect 380 7530 576 7538
rect 732 7590 928 7600
rect 732 7538 739 7590
rect 791 7538 803 7590
rect 855 7538 867 7590
rect 919 7538 928 7590
rect 732 7530 928 7538
rect 400 6530 596 6538
rect 400 6478 407 6530
rect 459 6478 471 6530
rect 523 6478 535 6530
rect 587 6478 596 6530
rect 400 6468 596 6478
rect 753 6530 949 6538
rect 753 6478 760 6530
rect 812 6478 824 6530
rect 876 6478 888 6530
rect 940 6478 949 6530
rect 753 6468 949 6478
rect 4759 6370 8311 7698
rect -25399 6362 -24551 6370
rect -25399 6310 -24738 6362
rect -24686 6310 -24674 6362
rect -24622 6310 -24610 6362
rect -24558 6310 -24551 6362
rect -25399 6300 -24551 6310
rect -16372 6362 -16176 6370
rect -16372 6310 -16363 6362
rect -16311 6310 -16299 6362
rect -16247 6310 -16235 6362
rect -16183 6310 -16176 6362
rect -16372 6300 -16176 6310
rect -15969 6362 -15773 6370
rect -15969 6310 -15960 6362
rect -15908 6310 -15896 6362
rect -15844 6310 -15832 6362
rect -15780 6310 -15773 6362
rect -15969 6300 -15773 6310
rect -7677 6362 -3392 6370
rect -7677 6310 -7668 6362
rect -7616 6310 -7604 6362
rect -7552 6310 -7540 6362
rect -7488 6310 -3579 6362
rect -3527 6310 -3515 6362
rect -3463 6310 -3451 6362
rect -3399 6310 -3392 6362
rect -7677 6300 -3392 6310
rect 4755 6362 8311 6370
rect 4755 6310 4764 6362
rect 4816 6310 4828 6362
rect 4880 6310 4892 6362
rect 4944 6310 8311 6362
rect 16824 6361 17024 7706
rect 4755 6300 8311 6310
rect 16846 6309 16858 6361
rect 16910 6309 17024 6361
rect -25399 4862 -24568 6300
rect -7560 4862 -3505 6300
rect 4759 4862 8311 6300
rect -25399 4852 -24551 4862
rect -25399 4800 -24738 4852
rect -24686 4800 -24674 4852
rect -24622 4800 -24610 4852
rect -24558 4800 -24551 4852
rect -25399 4792 -24551 4800
rect -16372 4852 -16176 4862
rect -16372 4800 -16363 4852
rect -16311 4800 -16299 4852
rect -16247 4800 -16235 4852
rect -16183 4800 -16176 4852
rect -16372 4792 -16176 4800
rect -15969 4852 -15773 4862
rect -15969 4800 -15960 4852
rect -15908 4800 -15896 4852
rect -15844 4800 -15832 4852
rect -15780 4800 -15773 4852
rect -15969 4792 -15773 4800
rect -7677 4852 -3392 4862
rect -7677 4800 -7668 4852
rect -7616 4800 -7604 4852
rect -7552 4800 -7540 4852
rect -7488 4800 -3579 4852
rect -3527 4800 -3515 4852
rect -3463 4800 -3451 4852
rect -3399 4800 -3392 4852
rect -7677 4792 -3392 4800
rect 4755 4852 8311 4862
rect 4755 4800 4764 4852
rect 4816 4800 4828 4852
rect 4880 4800 4892 4852
rect 4944 4851 8311 4852
rect 16824 4851 17024 6309
rect 4944 4800 8306 4851
rect 4755 4799 8306 4800
rect 16834 4799 16846 4851
rect 16898 4799 17024 4851
rect 4755 4792 8311 4799
rect -25399 2895 -24568 4792
rect -20704 4406 -20508 4416
rect -20704 4354 -20697 4406
rect -20645 4354 -20633 4406
rect -20581 4354 -20569 4406
rect -20517 4354 -20508 4406
rect -20704 4346 -20508 4354
rect -20383 4406 -20187 4416
rect -20383 4354 -20376 4406
rect -20324 4354 -20312 4406
rect -20260 4354 -20248 4406
rect -20196 4354 -20187 4406
rect -20383 4346 -20187 4354
rect -11998 4406 -11802 4416
rect -11998 4354 -11991 4406
rect -11939 4354 -11927 4406
rect -11875 4354 -11863 4406
rect -11811 4354 -11802 4406
rect -11998 4346 -11802 4354
rect -11659 4406 -11463 4416
rect -11659 4354 -11652 4406
rect -11600 4354 -11588 4406
rect -11536 4354 -11524 4406
rect -11472 4354 -11463 4406
rect -11659 4346 -11463 4354
rect -7560 2895 -3505 4792
rect 384 4406 580 4416
rect 384 4354 391 4406
rect 443 4354 455 4406
rect 507 4354 519 4406
rect 571 4354 580 4406
rect 384 4346 580 4354
rect 737 4406 933 4416
rect 737 4354 744 4406
rect 796 4354 808 4406
rect 860 4354 872 4406
rect 924 4354 933 4406
rect 737 4346 933 4354
rect 4759 2895 8311 4792
rect -25399 2885 -24560 2895
rect -25399 2833 -24747 2885
rect -24695 2833 -24683 2885
rect -24631 2833 -24619 2885
rect -24567 2833 -24560 2885
rect -25399 2825 -24560 2833
rect -16380 2885 -16184 2895
rect -16380 2833 -16371 2885
rect -16319 2833 -16307 2885
rect -16255 2833 -16243 2885
rect -16191 2833 -16184 2885
rect -16380 2825 -16184 2833
rect -15977 2885 -15781 2895
rect -15977 2833 -15968 2885
rect -15916 2833 -15904 2885
rect -15852 2833 -15840 2885
rect -15788 2833 -15781 2885
rect -15977 2825 -15781 2833
rect -7686 2885 -3401 2895
rect -7686 2833 -7677 2885
rect -7625 2833 -7613 2885
rect -7561 2833 -7549 2885
rect -7497 2833 -3588 2885
rect -3536 2833 -3524 2885
rect -3472 2833 -3460 2885
rect -3408 2833 -3401 2885
rect -7686 2825 -3401 2833
rect 4746 2885 8311 2895
rect 16824 2885 17024 4799
rect 4746 2833 4755 2885
rect 4807 2833 4819 2885
rect 4871 2833 4883 2885
rect 4935 2833 8311 2885
rect 16860 2833 16872 2885
rect 16924 2833 17024 2885
rect 4746 2825 8311 2833
rect -25399 2584 -24568 2825
rect -20686 2716 -20490 2726
rect -20686 2664 -20679 2716
rect -20627 2664 -20615 2716
rect -20563 2664 -20551 2716
rect -20499 2664 -20490 2716
rect -20686 2656 -20490 2664
rect -20365 2716 -20169 2726
rect -20365 2664 -20358 2716
rect -20306 2664 -20294 2716
rect -20242 2664 -20230 2716
rect -20178 2664 -20169 2716
rect -20365 2656 -20169 2664
rect -11980 2716 -11784 2726
rect -11980 2664 -11973 2716
rect -11921 2664 -11909 2716
rect -11857 2664 -11845 2716
rect -11793 2664 -11784 2716
rect -11980 2656 -11784 2664
rect -11641 2716 -11445 2726
rect -11641 2664 -11634 2716
rect -11582 2664 -11570 2716
rect -11518 2664 -11506 2716
rect -11454 2664 -11445 2716
rect -11641 2656 -11445 2664
rect -7560 2584 -3505 2825
rect 402 2716 598 2726
rect 402 2664 409 2716
rect 461 2664 473 2716
rect 525 2664 537 2716
rect 589 2664 598 2716
rect 402 2656 598 2664
rect 755 2716 951 2726
rect 755 2664 762 2716
rect 814 2664 826 2716
rect 878 2664 890 2716
rect 942 2664 951 2716
rect 755 2656 951 2664
rect 4759 2584 8311 2825
rect 16824 2584 17024 2833
rect -25399 1289 17024 2584
rect -25399 -7610 -24989 1289
rect -16981 -7610 -15305 1289
rect -7178 -7610 -3423 1289
rect 4759 -5343 8311 1289
rect 16824 1040 17024 1289
rect 16861 988 16873 1040
rect 16925 988 17024 1040
rect 16824 -926 17024 988
rect 16847 -978 16859 -926
rect 16911 -978 17024 -926
rect 16824 -2436 17024 -978
rect 16850 -2488 16862 -2436
rect 16914 -2488 17024 -2436
rect 16824 -3833 17024 -2488
rect 16846 -3885 16858 -3833
rect 16910 -3885 17024 -3833
rect 16824 -5343 17024 -3885
rect 4759 -5395 8306 -5343
rect 16834 -5395 16846 -5343
rect 16898 -5395 17024 -5343
rect 4759 -7610 8311 -5395
rect 16824 -7309 17024 -5395
rect 16860 -7361 16872 -7309
rect 16924 -7361 17024 -7309
rect 16824 -7610 17024 -7361
rect -25399 -8030 17024 -7610
rect -2711 -9828 16785 -9521
rect -2711 -9917 16722 -9828
rect -2711 -13240 -520 -9917
rect 2266 -13240 9108 -9917
rect 12290 -13240 13427 -9917
rect -2711 -13417 16651 -13240
rect -2711 -14407 16785 -13417
rect -2577 -14552 16785 -14407
rect 4126 -14611 9375 -14552
rect -2631 -14619 -2435 -14611
rect -2631 -14671 -2622 -14619
rect -2570 -14671 -2558 -14619
rect -2506 -14671 -2494 -14619
rect -2442 -14671 -2435 -14619
rect -2631 -14681 -2435 -14671
rect 4126 -14619 9428 -14611
rect 4126 -14671 4208 -14619
rect 4260 -14671 4272 -14619
rect 4324 -14671 4336 -14619
rect 4388 -14671 9241 -14619
rect 9293 -14671 9305 -14619
rect 9357 -14671 9369 -14619
rect 9421 -14671 9428 -14619
rect 4126 -14681 9428 -14671
rect 15975 -14619 16785 -14552
rect 15975 -14671 16107 -14619
rect 16159 -14671 16171 -14619
rect 16223 -14671 16235 -14619
rect 16287 -14671 16785 -14619
rect 649 -14734 845 -14726
rect 649 -14786 658 -14734
rect 710 -14786 722 -14734
rect 774 -14786 786 -14734
rect 838 -14786 845 -14734
rect 649 -14796 845 -14786
rect 1030 -14734 1226 -14726
rect 1030 -14786 1039 -14734
rect 1091 -14786 1103 -14734
rect 1155 -14786 1167 -14734
rect 1219 -14786 1226 -14734
rect 1030 -14796 1226 -14786
rect 4126 -16234 9375 -14681
rect 12495 -14734 12691 -14726
rect 12495 -14786 12504 -14734
rect 12556 -14786 12568 -14734
rect 12620 -14786 12632 -14734
rect 12684 -14786 12691 -14734
rect 12495 -14796 12691 -14786
rect 12909 -14734 13105 -14726
rect 12909 -14786 12918 -14734
rect 12970 -14786 12982 -14734
rect 13034 -14786 13046 -14734
rect 13098 -14786 13105 -14734
rect 12909 -14796 13105 -14786
rect -2640 -16244 -2444 -16234
rect -2640 -16296 -2633 -16244
rect -2581 -16296 -2569 -16244
rect -2517 -16296 -2505 -16244
rect -2453 -16296 -2444 -16244
rect -2640 -16304 -2444 -16296
rect 4126 -16244 9419 -16234
rect 4126 -16296 4197 -16244
rect 4249 -16296 4261 -16244
rect 4313 -16296 4325 -16244
rect 4377 -16296 9230 -16244
rect 9282 -16296 9294 -16244
rect 9346 -16296 9358 -16244
rect 9410 -16296 9419 -16244
rect 4126 -16304 9419 -16296
rect 15975 -16244 16785 -14671
rect 15975 -16296 16096 -16244
rect 16148 -16296 16160 -16244
rect 16212 -16296 16224 -16244
rect 16276 -16296 16785 -16244
rect 623 -16343 819 -16333
rect 623 -16395 630 -16343
rect 682 -16395 694 -16343
rect 746 -16395 758 -16343
rect 810 -16395 819 -16343
rect 623 -16403 819 -16395
rect 1004 -16343 1200 -16333
rect 1004 -16395 1011 -16343
rect 1063 -16395 1075 -16343
rect 1127 -16395 1139 -16343
rect 1191 -16395 1200 -16343
rect 1004 -16403 1200 -16395
rect 601 -17626 797 -17616
rect 601 -17678 608 -17626
rect 660 -17678 672 -17626
rect 724 -17678 736 -17626
rect 788 -17678 797 -17626
rect 601 -17686 797 -17678
rect 981 -17626 1177 -17616
rect 981 -17678 988 -17626
rect 1040 -17678 1052 -17626
rect 1104 -17678 1116 -17626
rect 1168 -17678 1177 -17626
rect 981 -17686 1177 -17678
rect 4126 -17715 9375 -16304
rect 12469 -16343 12665 -16333
rect 12469 -16395 12476 -16343
rect 12528 -16395 12540 -16343
rect 12592 -16395 12604 -16343
rect 12656 -16395 12665 -16343
rect 12469 -16403 12665 -16395
rect 12883 -16343 13079 -16333
rect 12883 -16395 12890 -16343
rect 12942 -16395 12954 -16343
rect 13006 -16395 13018 -16343
rect 13070 -16395 13079 -16343
rect 12883 -16403 13079 -16395
rect 12446 -17626 12642 -17616
rect 12446 -17678 12453 -17626
rect 12505 -17678 12517 -17626
rect 12569 -17678 12581 -17626
rect 12633 -17678 12642 -17626
rect 12446 -17686 12642 -17678
rect 12860 -17626 13056 -17616
rect 12860 -17678 12867 -17626
rect 12919 -17678 12931 -17626
rect 12983 -17678 12995 -17626
rect 13047 -17678 13056 -17626
rect 12860 -17686 13056 -17678
rect -2633 -17725 -2437 -17715
rect -2633 -17777 -2626 -17725
rect -2574 -17777 -2562 -17725
rect -2510 -17777 -2498 -17725
rect -2446 -17777 -2437 -17725
rect -2633 -17785 -2437 -17777
rect 4126 -17725 9426 -17715
rect 4126 -17777 4204 -17725
rect 4256 -17777 4268 -17725
rect 4320 -17777 4332 -17725
rect 4384 -17777 9237 -17725
rect 9289 -17777 9301 -17725
rect 9353 -17777 9365 -17725
rect 9417 -17777 9426 -17725
rect 4126 -17785 9426 -17777
rect 15975 -17725 16785 -16296
rect 15975 -17777 16103 -17725
rect 16155 -17777 16167 -17725
rect 16219 -17777 16231 -17725
rect 16283 -17777 16785 -17725
rect 4126 -17874 9375 -17785
rect 15975 -17874 16785 -17777
rect -2649 -17955 16785 -17874
rect -2711 -18271 16785 -17955
<< via1 >>
rect -20679 11352 -20627 11404
rect -20615 11352 -20563 11404
rect -20551 11352 -20499 11404
rect -20357 11352 -20305 11404
rect -20293 11352 -20241 11404
rect -20229 11352 -20177 11404
rect -11972 11352 -11920 11404
rect -11908 11352 -11856 11404
rect -11844 11352 -11792 11404
rect -11633 11352 -11581 11404
rect -11569 11352 -11517 11404
rect -11505 11352 -11453 11404
rect 410 11352 462 11404
rect 474 11352 526 11404
rect 538 11352 590 11404
rect 762 11352 814 11404
rect 826 11352 878 11404
rect 890 11352 942 11404
rect 12398 11351 12450 11403
rect 12462 11351 12514 11403
rect 12526 11351 12578 11403
rect 12689 11351 12741 11403
rect 12753 11351 12805 11403
rect 12817 11351 12869 11403
rect -24747 11183 -24695 11235
rect -24683 11183 -24631 11235
rect -24619 11183 -24567 11235
rect -16371 11183 -16319 11235
rect -16307 11183 -16255 11235
rect -16243 11183 -16191 11235
rect -15968 11183 -15916 11235
rect -15904 11183 -15852 11235
rect -15840 11183 -15788 11235
rect -7677 11183 -7625 11235
rect -7613 11183 -7561 11235
rect -7549 11183 -7497 11235
rect -3588 11183 -3536 11235
rect -3524 11183 -3472 11235
rect -3460 11183 -3408 11235
rect 4755 11183 4807 11235
rect 4819 11183 4871 11235
rect 4883 11183 4935 11235
rect 8333 11182 8385 11234
rect 8397 11182 8449 11234
rect 8461 11182 8513 11234
rect 16745 11182 16797 11234
rect 16809 11182 16861 11234
rect 16873 11182 16925 11234
rect -20678 9662 -20626 9714
rect -20614 9662 -20562 9714
rect -20550 9662 -20498 9714
rect -20356 9662 -20304 9714
rect -20292 9662 -20240 9714
rect -20228 9662 -20176 9714
rect -11971 9662 -11919 9714
rect -11907 9662 -11855 9714
rect -11843 9662 -11791 9714
rect -11633 9662 -11581 9714
rect -11569 9662 -11517 9714
rect -11505 9662 -11453 9714
rect 411 9662 463 9714
rect 475 9662 527 9714
rect 539 9662 591 9714
rect 763 9662 815 9714
rect 827 9662 879 9714
rect 891 9662 943 9714
rect 12385 9661 12437 9713
rect 12449 9661 12501 9713
rect 12513 9661 12565 9713
rect 12670 9661 12722 9713
rect 12734 9661 12786 9713
rect 12798 9661 12850 9713
rect -24745 9216 -24693 9268
rect -24681 9216 -24629 9268
rect -24617 9216 -24565 9268
rect -16370 9216 -16318 9268
rect -16306 9216 -16254 9268
rect -16242 9216 -16190 9268
rect -15967 9216 -15915 9268
rect -15903 9216 -15851 9268
rect -15839 9216 -15787 9268
rect -7675 9216 -7623 9268
rect -7611 9216 -7559 9268
rect -7547 9216 -7495 9268
rect -3586 9216 -3534 9268
rect -3522 9216 -3470 9268
rect -3458 9216 -3406 9268
rect 4757 9216 4809 9268
rect 4821 9216 4873 9268
rect 4885 9216 4937 9268
rect 8320 9216 8372 9268
rect 8384 9216 8436 9268
rect 8448 9216 8500 9268
rect 16731 9216 16783 9268
rect 16795 9216 16847 9268
rect 16859 9216 16911 9268
rect -24749 7706 -24697 7758
rect -24685 7706 -24633 7758
rect -24621 7706 -24569 7758
rect -16374 7706 -16322 7758
rect -16310 7706 -16258 7758
rect -16246 7706 -16194 7758
rect -15971 7706 -15919 7758
rect -15907 7706 -15855 7758
rect -15843 7706 -15791 7758
rect -7679 7706 -7627 7758
rect -7615 7706 -7563 7758
rect -7551 7706 -7499 7758
rect -3590 7706 -3538 7758
rect -3526 7706 -3474 7758
rect -3462 7706 -3410 7758
rect 4753 7706 4805 7758
rect 4817 7706 4869 7758
rect 4881 7706 4933 7758
rect 8323 7706 8375 7758
rect 8387 7706 8439 7758
rect 8451 7706 8503 7758
rect 16734 7706 16786 7758
rect 16798 7706 16850 7758
rect 16862 7706 16914 7758
rect -20702 7538 -20650 7590
rect -20638 7538 -20586 7590
rect -20574 7538 -20522 7590
rect -20380 7538 -20328 7590
rect -20316 7538 -20264 7590
rect -20252 7538 -20200 7590
rect -11995 7538 -11943 7590
rect -11931 7538 -11879 7590
rect -11867 7538 -11815 7590
rect -11656 7538 -11604 7590
rect -11592 7538 -11540 7590
rect -11528 7538 -11476 7590
rect -20681 6478 -20629 6530
rect -20617 6478 -20565 6530
rect -20553 6478 -20501 6530
rect -20360 6478 -20308 6530
rect -20296 6478 -20244 6530
rect -20232 6478 -20180 6530
rect -11974 6478 -11922 6530
rect -11910 6478 -11858 6530
rect -11846 6478 -11794 6530
rect -11636 6478 -11584 6530
rect -11572 6478 -11520 6530
rect -11508 6478 -11456 6530
rect 387 7538 439 7590
rect 451 7538 503 7590
rect 515 7538 567 7590
rect 739 7538 791 7590
rect 803 7538 855 7590
rect 867 7538 919 7590
rect 407 6478 459 6530
rect 471 6478 523 6530
rect 535 6478 587 6530
rect 760 6478 812 6530
rect 824 6478 876 6530
rect 888 6478 940 6530
rect 12384 7537 12436 7589
rect 12448 7537 12500 7589
rect 12512 7537 12564 7589
rect 12685 7537 12737 7589
rect 12749 7537 12801 7589
rect 12813 7537 12865 7589
rect 12363 6478 12415 6530
rect 12427 6478 12479 6530
rect 12491 6478 12543 6530
rect 12674 6478 12726 6530
rect 12738 6478 12790 6530
rect 12802 6478 12854 6530
rect -24738 6310 -24686 6362
rect -24674 6310 -24622 6362
rect -24610 6310 -24558 6362
rect -16363 6310 -16311 6362
rect -16299 6310 -16247 6362
rect -16235 6310 -16183 6362
rect -15960 6310 -15908 6362
rect -15896 6310 -15844 6362
rect -15832 6310 -15780 6362
rect -7668 6310 -7616 6362
rect -7604 6310 -7552 6362
rect -7540 6310 -7488 6362
rect -3579 6310 -3527 6362
rect -3515 6310 -3463 6362
rect -3451 6310 -3399 6362
rect 4764 6310 4816 6362
rect 4828 6310 4880 6362
rect 4892 6310 4944 6362
rect 8319 6309 8371 6361
rect 8383 6309 8435 6361
rect 8447 6309 8499 6361
rect 16730 6309 16782 6361
rect 16794 6309 16846 6361
rect 16858 6309 16910 6361
rect -24738 4800 -24686 4852
rect -24674 4800 -24622 4852
rect -24610 4800 -24558 4852
rect -16363 4800 -16311 4852
rect -16299 4800 -16247 4852
rect -16235 4800 -16183 4852
rect -15960 4800 -15908 4852
rect -15896 4800 -15844 4852
rect -15832 4800 -15780 4852
rect -7668 4800 -7616 4852
rect -7604 4800 -7552 4852
rect -7540 4800 -7488 4852
rect -3579 4800 -3527 4852
rect -3515 4800 -3463 4852
rect -3451 4800 -3399 4852
rect 4764 4800 4816 4852
rect 4828 4800 4880 4852
rect 4892 4800 4944 4852
rect 8306 4799 8358 4851
rect 8370 4799 8422 4851
rect 8434 4799 8486 4851
rect 16718 4799 16770 4851
rect 16782 4799 16834 4851
rect 16846 4799 16898 4851
rect -20697 4354 -20645 4406
rect -20633 4354 -20581 4406
rect -20569 4354 -20517 4406
rect -20376 4354 -20324 4406
rect -20312 4354 -20260 4406
rect -20248 4354 -20196 4406
rect -11991 4354 -11939 4406
rect -11927 4354 -11875 4406
rect -11863 4354 -11811 4406
rect -11652 4354 -11600 4406
rect -11588 4354 -11536 4406
rect -11524 4354 -11472 4406
rect 391 4354 443 4406
rect 455 4354 507 4406
rect 519 4354 571 4406
rect 744 4354 796 4406
rect 808 4354 860 4406
rect 872 4354 924 4406
rect 12392 4354 12444 4406
rect 12456 4354 12508 4406
rect 12520 4354 12572 4406
rect 12699 4354 12751 4406
rect 12763 4354 12815 4406
rect 12827 4354 12879 4406
rect -24747 2833 -24695 2885
rect -24683 2833 -24631 2885
rect -24619 2833 -24567 2885
rect -16371 2833 -16319 2885
rect -16307 2833 -16255 2885
rect -16243 2833 -16191 2885
rect -15968 2833 -15916 2885
rect -15904 2833 -15852 2885
rect -15840 2833 -15788 2885
rect -7677 2833 -7625 2885
rect -7613 2833 -7561 2885
rect -7549 2833 -7497 2885
rect -3588 2833 -3536 2885
rect -3524 2833 -3472 2885
rect -3460 2833 -3408 2885
rect 4755 2833 4807 2885
rect 4819 2833 4871 2885
rect 4883 2833 4935 2885
rect 8333 2833 8385 2885
rect 8397 2833 8449 2885
rect 8461 2833 8513 2885
rect 16744 2833 16796 2885
rect 16808 2833 16860 2885
rect 16872 2833 16924 2885
rect -20679 2664 -20627 2716
rect -20615 2664 -20563 2716
rect -20551 2664 -20499 2716
rect -20358 2664 -20306 2716
rect -20294 2664 -20242 2716
rect -20230 2664 -20178 2716
rect -11973 2664 -11921 2716
rect -11909 2664 -11857 2716
rect -11845 2664 -11793 2716
rect -11634 2664 -11582 2716
rect -11570 2664 -11518 2716
rect -11506 2664 -11454 2716
rect 409 2664 461 2716
rect 473 2664 525 2716
rect 537 2664 589 2716
rect 762 2664 814 2716
rect 826 2664 878 2716
rect 890 2664 942 2716
rect 12376 2664 12428 2716
rect 12440 2664 12492 2716
rect 12504 2664 12556 2716
rect 12673 2664 12725 2716
rect 12737 2664 12789 2716
rect 12801 2664 12853 2716
rect 12398 1157 12450 1209
rect 12462 1157 12514 1209
rect 12526 1157 12578 1209
rect 12689 1157 12741 1209
rect 12753 1157 12805 1209
rect 12817 1157 12869 1209
rect 8333 988 8385 1040
rect 8397 988 8449 1040
rect 8461 988 8513 1040
rect 16745 988 16797 1040
rect 16809 988 16861 1040
rect 16873 988 16925 1040
rect 12385 -533 12437 -481
rect 12449 -533 12501 -481
rect 12513 -533 12565 -481
rect 12670 -533 12722 -481
rect 12734 -533 12786 -481
rect 12798 -533 12850 -481
rect 8320 -978 8372 -926
rect 8384 -978 8436 -926
rect 8448 -978 8500 -926
rect 16731 -978 16783 -926
rect 16795 -978 16847 -926
rect 16859 -978 16911 -926
rect 8323 -2488 8375 -2436
rect 8387 -2488 8439 -2436
rect 8451 -2488 8503 -2436
rect 16734 -2488 16786 -2436
rect 16798 -2488 16850 -2436
rect 16862 -2488 16914 -2436
rect 12384 -2657 12436 -2605
rect 12448 -2657 12500 -2605
rect 12512 -2657 12564 -2605
rect 12685 -2657 12737 -2605
rect 12749 -2657 12801 -2605
rect 12813 -2657 12865 -2605
rect 12363 -3716 12415 -3664
rect 12427 -3716 12479 -3664
rect 12491 -3716 12543 -3664
rect 12674 -3716 12726 -3664
rect 12738 -3716 12790 -3664
rect 12802 -3716 12854 -3664
rect 8319 -3885 8371 -3833
rect 8383 -3885 8435 -3833
rect 8447 -3885 8499 -3833
rect 16730 -3885 16782 -3833
rect 16794 -3885 16846 -3833
rect 16858 -3885 16910 -3833
rect 8306 -5395 8358 -5343
rect 8370 -5395 8422 -5343
rect 8434 -5395 8486 -5343
rect 16718 -5395 16770 -5343
rect 16782 -5395 16834 -5343
rect 16846 -5395 16898 -5343
rect 12392 -5840 12444 -5788
rect 12456 -5840 12508 -5788
rect 12520 -5840 12572 -5788
rect 12699 -5840 12751 -5788
rect 12763 -5840 12815 -5788
rect 12827 -5840 12879 -5788
rect 8333 -7361 8385 -7309
rect 8397 -7361 8449 -7309
rect 8461 -7361 8513 -7309
rect 16744 -7361 16796 -7309
rect 16808 -7361 16860 -7309
rect 16872 -7361 16924 -7309
rect 12376 -7530 12428 -7478
rect 12440 -7530 12492 -7478
rect 12504 -7530 12556 -7478
rect 12673 -7530 12725 -7478
rect 12737 -7530 12789 -7478
rect 12801 -7530 12853 -7478
rect -2622 -14671 -2570 -14619
rect -2558 -14671 -2506 -14619
rect -2494 -14671 -2442 -14619
rect 4208 -14671 4260 -14619
rect 4272 -14671 4324 -14619
rect 4336 -14671 4388 -14619
rect 9241 -14671 9293 -14619
rect 9305 -14671 9357 -14619
rect 9369 -14671 9421 -14619
rect 16107 -14671 16159 -14619
rect 16171 -14671 16223 -14619
rect 16235 -14671 16287 -14619
rect 658 -14786 710 -14734
rect 722 -14786 774 -14734
rect 786 -14786 838 -14734
rect 1039 -14786 1091 -14734
rect 1103 -14786 1155 -14734
rect 1167 -14786 1219 -14734
rect 12504 -14786 12556 -14734
rect 12568 -14786 12620 -14734
rect 12632 -14786 12684 -14734
rect 12918 -14786 12970 -14734
rect 12982 -14786 13034 -14734
rect 13046 -14786 13098 -14734
rect -2633 -16296 -2581 -16244
rect -2569 -16296 -2517 -16244
rect -2505 -16296 -2453 -16244
rect 4197 -16296 4249 -16244
rect 4261 -16296 4313 -16244
rect 4325 -16296 4377 -16244
rect 9230 -16296 9282 -16244
rect 9294 -16296 9346 -16244
rect 9358 -16296 9410 -16244
rect 16096 -16296 16148 -16244
rect 16160 -16296 16212 -16244
rect 16224 -16296 16276 -16244
rect 630 -16395 682 -16343
rect 694 -16395 746 -16343
rect 758 -16395 810 -16343
rect 1011 -16395 1063 -16343
rect 1075 -16395 1127 -16343
rect 1139 -16395 1191 -16343
rect 608 -17678 660 -17626
rect 672 -17678 724 -17626
rect 736 -17678 788 -17626
rect 988 -17678 1040 -17626
rect 1052 -17678 1104 -17626
rect 1116 -17678 1168 -17626
rect 12476 -16395 12528 -16343
rect 12540 -16395 12592 -16343
rect 12604 -16395 12656 -16343
rect 12890 -16395 12942 -16343
rect 12954 -16395 13006 -16343
rect 13018 -16395 13070 -16343
rect 12453 -17678 12505 -17626
rect 12517 -17678 12569 -17626
rect 12581 -17678 12633 -17626
rect 12867 -17678 12919 -17626
rect 12931 -17678 12983 -17626
rect 12995 -17678 13047 -17626
rect -2626 -17777 -2574 -17725
rect -2562 -17777 -2510 -17725
rect -2498 -17777 -2446 -17725
rect 4204 -17777 4256 -17725
rect 4268 -17777 4320 -17725
rect 4332 -17777 4384 -17725
rect 9237 -17777 9289 -17725
rect 9301 -17777 9353 -17725
rect 9365 -17777 9417 -17725
rect 16103 -17777 16155 -17725
rect 16167 -17777 16219 -17725
rect 16231 -17777 16283 -17725
<< metal2 >>
rect -20686 11404 -20490 11412
rect -20686 11352 -20679 11404
rect -20627 11352 -20615 11404
rect -20563 11352 -20551 11404
rect -20499 11352 -20490 11404
rect -20686 11342 -20490 11352
rect -20364 11404 -20168 11412
rect -20364 11352 -20357 11404
rect -20305 11352 -20293 11404
rect -20241 11352 -20229 11404
rect -20177 11352 -20168 11404
rect -20364 11342 -20168 11352
rect -11979 11404 -11783 11412
rect -11979 11352 -11972 11404
rect -11920 11352 -11908 11404
rect -11856 11352 -11844 11404
rect -11792 11352 -11783 11404
rect -11979 11342 -11783 11352
rect -11640 11404 -11444 11412
rect -11640 11352 -11633 11404
rect -11581 11352 -11569 11404
rect -11517 11352 -11505 11404
rect -11453 11352 -11444 11404
rect -11640 11342 -11444 11352
rect 403 11404 599 11412
rect 403 11352 410 11404
rect 462 11352 474 11404
rect 526 11352 538 11404
rect 590 11352 599 11404
rect 403 11342 599 11352
rect 755 11404 951 11412
rect 755 11352 762 11404
rect 814 11352 826 11404
rect 878 11352 890 11404
rect 942 11352 951 11404
rect 755 11342 951 11352
rect 12389 11403 12585 11411
rect 12389 11351 12398 11403
rect 12450 11351 12462 11403
rect 12514 11351 12526 11403
rect 12578 11351 12585 11403
rect 12389 11341 12585 11351
rect 12680 11403 12876 11411
rect 12680 11351 12689 11403
rect 12741 11351 12753 11403
rect 12805 11351 12817 11403
rect 12869 11351 12876 11403
rect 12680 11341 12876 11351
rect -24756 11235 -24560 11243
rect -24756 11183 -24747 11235
rect -24695 11183 -24683 11235
rect -24631 11183 -24619 11235
rect -24567 11183 -24560 11235
rect -24756 11173 -24560 11183
rect -16380 11235 -16184 11243
rect -16380 11183 -16371 11235
rect -16319 11183 -16307 11235
rect -16255 11183 -16243 11235
rect -16191 11183 -16184 11235
rect -16380 11173 -16184 11183
rect -15977 11235 -15781 11243
rect -15977 11183 -15968 11235
rect -15916 11183 -15904 11235
rect -15852 11183 -15840 11235
rect -15788 11183 -15781 11235
rect -15977 11173 -15781 11183
rect -7686 11235 -7490 11243
rect -7686 11183 -7677 11235
rect -7625 11183 -7613 11235
rect -7561 11183 -7549 11235
rect -7497 11183 -7490 11235
rect -7686 11173 -7490 11183
rect -3597 11235 -3401 11243
rect -3597 11183 -3588 11235
rect -3536 11183 -3524 11235
rect -3472 11183 -3460 11235
rect -3408 11183 -3401 11235
rect -3597 11173 -3401 11183
rect 4746 11235 4942 11243
rect 4746 11183 4755 11235
rect 4807 11183 4819 11235
rect 4871 11183 4883 11235
rect 4935 11183 4942 11235
rect 4746 11173 4942 11183
rect 8324 11234 8520 11242
rect 8324 11182 8333 11234
rect 8385 11182 8397 11234
rect 8449 11182 8461 11234
rect 8513 11182 8520 11234
rect 8324 11172 8520 11182
rect 16736 11234 16932 11242
rect 16736 11182 16745 11234
rect 16797 11182 16809 11234
rect 16861 11182 16873 11234
rect 16925 11182 16932 11234
rect 16736 11172 16932 11182
rect -25759 10498 -25459 10510
rect -6617 10498 -6317 10510
rect -25759 10488 -22599 10498
rect -25759 10432 -25719 10488
rect -25663 10432 -25639 10488
rect -25583 10432 -25559 10488
rect -25503 10432 -22599 10488
rect -25759 10410 -22599 10432
rect -9476 10488 -6317 10498
rect -9476 10432 -6573 10488
rect -6517 10432 -6493 10488
rect -6437 10432 -6413 10488
rect -6357 10432 -6317 10488
rect -9476 10410 -6317 10432
rect -4750 10498 -4450 10510
rect 5753 10498 6053 10510
rect 6889 10498 7189 10510
rect 9816 10498 10116 10510
rect 15130 10498 15430 10510
rect 18395 10498 18695 10510
rect -4750 10488 -1553 10498
rect -4750 10432 -4706 10488
rect -4650 10432 -4626 10488
rect -4570 10432 -4546 10488
rect -4490 10432 -1553 10488
rect -4750 10410 -1553 10432
rect 2855 10488 8912 10498
rect 2855 10432 5793 10488
rect 5849 10432 5873 10488
rect 5929 10432 5953 10488
rect 6009 10432 6929 10488
rect 6985 10432 7009 10488
rect 7065 10432 7089 10488
rect 7145 10432 8912 10488
rect 2855 10410 8912 10432
rect 9816 10410 15430 10498
rect 15536 10488 18695 10498
rect 15536 10432 18435 10488
rect 18491 10432 18515 10488
rect 18571 10432 18595 10488
rect 18651 10432 18695 10488
rect 15536 10410 18695 10432
rect -25759 10178 -25459 10190
rect -6617 10178 -6317 10190
rect 5753 10178 6053 10189
rect 6889 10178 7189 10189
rect 10784 10178 11084 10189
rect 14162 10178 14462 10189
rect 18395 10178 18695 10189
rect -25759 10168 -22599 10178
rect -25759 10112 -25719 10168
rect -25663 10112 -25639 10168
rect -25583 10112 -25559 10168
rect -25503 10112 -22599 10168
rect -25759 10090 -22599 10112
rect -9476 10168 -6317 10178
rect -9476 10112 -6573 10168
rect -6517 10112 -6493 10168
rect -6437 10112 -6413 10168
rect -6357 10112 -6317 10168
rect -9476 10090 -6317 10112
rect -4712 10089 -1553 10178
rect 2855 10167 8912 10178
rect 2855 10111 5793 10167
rect 5849 10111 5873 10167
rect 5929 10111 5953 10167
rect 6009 10111 6929 10167
rect 6985 10111 7009 10167
rect 7065 10111 7089 10167
rect 7145 10111 8912 10167
rect 2855 10089 8912 10111
rect 10784 10089 14462 10178
rect 15536 10167 18695 10178
rect 15536 10111 18435 10167
rect 18491 10111 18515 10167
rect 18571 10111 18595 10167
rect 18651 10111 18695 10167
rect 15536 10089 18695 10111
rect -20685 9714 -20489 9722
rect -20685 9662 -20678 9714
rect -20626 9662 -20614 9714
rect -20562 9662 -20550 9714
rect -20498 9662 -20489 9714
rect -20685 9652 -20489 9662
rect -20363 9714 -20167 9722
rect -20363 9662 -20356 9714
rect -20304 9662 -20292 9714
rect -20240 9662 -20228 9714
rect -20176 9662 -20167 9714
rect -20363 9652 -20167 9662
rect -11978 9714 -11782 9722
rect -11978 9662 -11971 9714
rect -11919 9662 -11907 9714
rect -11855 9662 -11843 9714
rect -11791 9662 -11782 9714
rect -11978 9652 -11782 9662
rect -11640 9714 -11444 9722
rect -11640 9662 -11633 9714
rect -11581 9662 -11569 9714
rect -11517 9662 -11505 9714
rect -11453 9662 -11444 9714
rect -11640 9652 -11444 9662
rect 404 9714 600 9722
rect 404 9662 411 9714
rect 463 9662 475 9714
rect 527 9662 539 9714
rect 591 9662 600 9714
rect 404 9652 600 9662
rect 756 9714 952 9722
rect 756 9662 763 9714
rect 815 9662 827 9714
rect 879 9662 891 9714
rect 943 9662 952 9714
rect 756 9652 952 9662
rect 12376 9713 12572 9721
rect 12376 9661 12385 9713
rect 12437 9661 12449 9713
rect 12501 9661 12513 9713
rect 12565 9661 12572 9713
rect 12376 9651 12572 9661
rect 12661 9713 12857 9721
rect 12661 9661 12670 9713
rect 12722 9661 12734 9713
rect 12786 9661 12798 9713
rect 12850 9661 12857 9713
rect 12661 9651 12857 9661
rect 9816 9590 12150 9612
rect 9816 9534 9856 9590
rect 9912 9534 9936 9590
rect 9992 9534 10016 9590
rect 10072 9534 12150 9590
rect 9816 9512 12150 9534
rect 13101 9590 15430 9612
rect 13101 9534 15170 9590
rect 15226 9534 15250 9590
rect 15306 9534 15330 9590
rect 15386 9534 15430 9590
rect 13101 9512 15430 9534
rect 10784 9429 14468 9451
rect 10784 9373 10828 9429
rect 10884 9373 10908 9429
rect 10964 9373 10988 9429
rect 11044 9373 14206 9429
rect 14262 9373 14286 9429
rect 14342 9373 14366 9429
rect 14422 9373 14468 9429
rect 10784 9351 14468 9373
rect -24754 9268 -24558 9276
rect -24754 9216 -24745 9268
rect -24693 9216 -24681 9268
rect -24629 9216 -24617 9268
rect -24565 9216 -24558 9268
rect -24754 9206 -24558 9216
rect -16379 9268 -16183 9276
rect -16379 9216 -16370 9268
rect -16318 9216 -16306 9268
rect -16254 9216 -16242 9268
rect -16190 9216 -16183 9268
rect -16379 9206 -16183 9216
rect -15976 9268 -15780 9276
rect -15976 9216 -15967 9268
rect -15915 9216 -15903 9268
rect -15851 9216 -15839 9268
rect -15787 9216 -15780 9268
rect -15976 9206 -15780 9216
rect -7684 9268 -7488 9276
rect -7684 9216 -7675 9268
rect -7623 9216 -7611 9268
rect -7559 9216 -7547 9268
rect -7495 9216 -7488 9268
rect -7684 9206 -7488 9216
rect -3595 9268 -3399 9276
rect -3595 9216 -3586 9268
rect -3534 9216 -3522 9268
rect -3470 9216 -3458 9268
rect -3406 9216 -3399 9268
rect -3595 9206 -3399 9216
rect 4748 9268 4944 9276
rect 4748 9216 4757 9268
rect 4809 9216 4821 9268
rect 4873 9216 4885 9268
rect 4937 9216 4944 9268
rect 4748 9206 4944 9216
rect 8311 9268 8507 9276
rect 8311 9216 8320 9268
rect 8372 9216 8384 9268
rect 8436 9216 8448 9268
rect 8500 9216 8507 9268
rect 8311 9206 8507 9216
rect 16722 9268 16918 9276
rect 16722 9216 16731 9268
rect 16783 9216 16795 9268
rect 16847 9216 16859 9268
rect 16911 9216 16918 9268
rect 16722 9206 16918 9216
rect -25759 8851 -25459 8863
rect -6617 8851 -6317 8863
rect 5753 8851 6053 8863
rect 6889 8851 7189 8863
rect 18395 8851 18695 8863
rect -25759 8841 -22599 8851
rect -25759 8785 -25719 8841
rect -25663 8785 -25639 8841
rect -25583 8785 -25559 8841
rect -25503 8785 -22599 8841
rect -25759 8763 -22599 8785
rect -9476 8841 -6317 8851
rect -9476 8785 -6573 8841
rect -6517 8785 -6493 8841
rect -6437 8785 -6413 8841
rect -6357 8785 -6317 8841
rect -9476 8763 -6317 8785
rect -4712 8763 -1553 8851
rect 2855 8841 8912 8851
rect 2855 8785 5793 8841
rect 5849 8785 5873 8841
rect 5929 8785 5953 8841
rect 6009 8785 6929 8841
rect 6985 8785 7009 8841
rect 7065 8785 7089 8841
rect 7145 8785 8912 8841
rect 2855 8763 8912 8785
rect 10784 8763 14462 8851
rect 15536 8841 18695 8851
rect 15536 8785 18435 8841
rect 18491 8785 18515 8841
rect 18571 8785 18595 8841
rect 18651 8785 18695 8841
rect 15536 8763 18695 8785
rect 10784 8751 11084 8763
rect 14162 8751 14462 8763
rect -25759 8509 -22599 8531
rect -25759 8453 -25719 8509
rect -25663 8453 -25639 8509
rect -25583 8453 -25559 8509
rect -25503 8453 -22599 8509
rect -25759 8443 -22599 8453
rect -9476 8509 -6317 8531
rect -9476 8453 -6573 8509
rect -6517 8453 -6493 8509
rect -6437 8453 -6413 8509
rect -6357 8453 -6317 8509
rect -9476 8443 -6317 8453
rect -25759 8431 -25459 8443
rect -6617 8431 -6317 8443
rect -4750 8509 -1553 8531
rect -4750 8453 -4706 8509
rect -4650 8453 -4626 8509
rect -4570 8453 -4546 8509
rect -4490 8453 -1553 8509
rect -4750 8442 -1553 8453
rect 2855 8509 8912 8531
rect 2855 8453 5793 8509
rect 5849 8453 5873 8509
rect 5929 8453 5953 8509
rect 6009 8453 6929 8509
rect 6985 8453 7009 8509
rect 7065 8453 7089 8509
rect 7145 8453 8912 8509
rect 2855 8442 8912 8453
rect 9816 8442 15430 8531
rect 15536 8509 18695 8531
rect 15536 8453 18435 8509
rect 18491 8453 18515 8509
rect 18571 8453 18595 8509
rect 18651 8453 18695 8509
rect 15536 8442 18695 8453
rect -4750 8431 -4450 8442
rect 5753 8431 6053 8442
rect 6889 8431 7189 8442
rect 9816 8431 10116 8442
rect 15130 8431 15430 8442
rect 18395 8431 18695 8442
rect 9816 8077 12150 8099
rect 9816 8021 9856 8077
rect 9912 8021 9936 8077
rect 9992 8021 10016 8077
rect 10072 8021 12150 8077
rect 9816 7999 12150 8021
rect 13101 8077 15430 8099
rect 13101 8021 15170 8077
rect 15226 8021 15250 8077
rect 15306 8021 15330 8077
rect 15386 8021 15430 8077
rect 13101 7999 15430 8021
rect 10784 7909 14462 7931
rect 10784 7853 10828 7909
rect 10884 7853 10908 7909
rect 10964 7853 10988 7909
rect 11044 7853 14206 7909
rect 14262 7853 14286 7909
rect 14342 7853 14366 7909
rect 14422 7853 14462 7909
rect 10784 7831 14462 7853
rect -24758 7758 -24562 7768
rect -24758 7706 -24749 7758
rect -24697 7706 -24685 7758
rect -24633 7706 -24621 7758
rect -24569 7706 -24562 7758
rect -24758 7698 -24562 7706
rect -16383 7758 -16187 7768
rect -16383 7706 -16374 7758
rect -16322 7706 -16310 7758
rect -16258 7706 -16246 7758
rect -16194 7706 -16187 7758
rect -16383 7698 -16187 7706
rect -15980 7758 -15784 7768
rect -15980 7706 -15971 7758
rect -15919 7706 -15907 7758
rect -15855 7706 -15843 7758
rect -15791 7706 -15784 7758
rect -15980 7698 -15784 7706
rect -7688 7758 -7492 7768
rect -7688 7706 -7679 7758
rect -7627 7706 -7615 7758
rect -7563 7706 -7551 7758
rect -7499 7706 -7492 7758
rect -7688 7698 -7492 7706
rect -3599 7758 -3403 7768
rect -3599 7706 -3590 7758
rect -3538 7706 -3526 7758
rect -3474 7706 -3462 7758
rect -3410 7706 -3403 7758
rect -3599 7698 -3403 7706
rect 4744 7758 4940 7768
rect 4744 7706 4753 7758
rect 4805 7706 4817 7758
rect 4869 7706 4881 7758
rect 4933 7706 4940 7758
rect 4744 7698 4940 7706
rect 8314 7758 8510 7768
rect 8314 7706 8323 7758
rect 8375 7706 8387 7758
rect 8439 7706 8451 7758
rect 8503 7706 8510 7758
rect 8314 7698 8510 7706
rect 16725 7758 16921 7768
rect 16725 7706 16734 7758
rect 16786 7706 16798 7758
rect 16850 7706 16862 7758
rect 16914 7706 16921 7758
rect 16725 7698 16921 7706
rect -20709 7590 -20513 7600
rect -20709 7538 -20702 7590
rect -20650 7538 -20638 7590
rect -20586 7538 -20574 7590
rect -20522 7538 -20513 7590
rect -20709 7530 -20513 7538
rect -20387 7590 -20191 7600
rect -20387 7538 -20380 7590
rect -20328 7538 -20316 7590
rect -20264 7538 -20252 7590
rect -20200 7538 -20191 7590
rect -20387 7530 -20191 7538
rect -12002 7590 -11806 7600
rect -12002 7538 -11995 7590
rect -11943 7538 -11931 7590
rect -11879 7538 -11867 7590
rect -11815 7538 -11806 7590
rect -12002 7530 -11806 7538
rect -11663 7590 -11467 7600
rect -11663 7538 -11656 7590
rect -11604 7538 -11592 7590
rect -11540 7538 -11528 7590
rect -11476 7538 -11467 7590
rect -11663 7530 -11467 7538
rect 380 7590 576 7600
rect 380 7538 387 7590
rect 439 7538 451 7590
rect 503 7538 515 7590
rect 567 7538 576 7590
rect 380 7530 576 7538
rect 732 7590 928 7600
rect 732 7538 739 7590
rect 791 7538 803 7590
rect 855 7538 867 7590
rect 919 7538 928 7590
rect 732 7530 928 7538
rect 12375 7589 12571 7599
rect 12375 7537 12384 7589
rect 12436 7537 12448 7589
rect 12500 7537 12512 7589
rect 12564 7537 12571 7589
rect 12375 7529 12571 7537
rect 12676 7589 12872 7599
rect 12676 7537 12685 7589
rect 12737 7537 12749 7589
rect 12801 7537 12813 7589
rect 12865 7537 12872 7589
rect 12676 7529 12872 7537
rect -20688 6530 -20492 6538
rect -20688 6478 -20681 6530
rect -20629 6478 -20617 6530
rect -20565 6478 -20553 6530
rect -20501 6478 -20492 6530
rect -20688 6468 -20492 6478
rect -20367 6530 -20171 6538
rect -20367 6478 -20360 6530
rect -20308 6478 -20296 6530
rect -20244 6478 -20232 6530
rect -20180 6478 -20171 6530
rect -20367 6468 -20171 6478
rect -11981 6530 -11785 6538
rect -11981 6478 -11974 6530
rect -11922 6478 -11910 6530
rect -11858 6478 -11846 6530
rect -11794 6478 -11785 6530
rect -11981 6468 -11785 6478
rect -11643 6530 -11447 6538
rect -11643 6478 -11636 6530
rect -11584 6478 -11572 6530
rect -11520 6478 -11508 6530
rect -11456 6478 -11447 6530
rect -11643 6468 -11447 6478
rect 400 6530 596 6538
rect 400 6478 407 6530
rect 459 6478 471 6530
rect 523 6478 535 6530
rect 587 6478 596 6530
rect 400 6468 596 6478
rect 753 6530 949 6538
rect 753 6478 760 6530
rect 812 6478 824 6530
rect 876 6478 888 6530
rect 940 6478 949 6530
rect 753 6468 949 6478
rect 12354 6530 12550 6538
rect 12354 6478 12363 6530
rect 12415 6478 12427 6530
rect 12479 6478 12491 6530
rect 12543 6478 12550 6530
rect 12354 6468 12550 6478
rect 12665 6530 12861 6538
rect 12665 6478 12674 6530
rect 12726 6478 12738 6530
rect 12790 6478 12802 6530
rect 12854 6478 12861 6530
rect 12665 6468 12861 6478
rect -24747 6362 -24551 6370
rect -24747 6310 -24738 6362
rect -24686 6310 -24674 6362
rect -24622 6310 -24610 6362
rect -24558 6310 -24551 6362
rect -24747 6300 -24551 6310
rect -16372 6362 -16176 6370
rect -16372 6310 -16363 6362
rect -16311 6310 -16299 6362
rect -16247 6310 -16235 6362
rect -16183 6310 -16176 6362
rect -16372 6300 -16176 6310
rect -15969 6362 -15773 6370
rect -15969 6310 -15960 6362
rect -15908 6310 -15896 6362
rect -15844 6310 -15832 6362
rect -15780 6310 -15773 6362
rect -15969 6300 -15773 6310
rect -7677 6362 -7481 6370
rect -7677 6310 -7668 6362
rect -7616 6310 -7604 6362
rect -7552 6310 -7540 6362
rect -7488 6310 -7481 6362
rect -7677 6300 -7481 6310
rect -3588 6362 -3392 6370
rect -3588 6310 -3579 6362
rect -3527 6310 -3515 6362
rect -3463 6310 -3451 6362
rect -3399 6310 -3392 6362
rect -3588 6300 -3392 6310
rect 4755 6362 4951 6370
rect 4755 6310 4764 6362
rect 4816 6310 4828 6362
rect 4880 6310 4892 6362
rect 4944 6310 4951 6362
rect 4755 6300 4951 6310
rect 8310 6361 8506 6369
rect 8310 6309 8319 6361
rect 8371 6309 8383 6361
rect 8435 6309 8447 6361
rect 8499 6309 8506 6361
rect 8310 6299 8506 6309
rect 16721 6361 16917 6369
rect 16721 6309 16730 6361
rect 16782 6309 16794 6361
rect 16846 6309 16858 6361
rect 16910 6309 16917 6361
rect 16721 6299 16917 6309
rect 10784 6215 14462 6237
rect 10784 6159 10828 6215
rect 10884 6159 10908 6215
rect 10964 6159 10988 6215
rect 11044 6159 14206 6215
rect 14262 6159 14286 6215
rect 14342 6159 14366 6215
rect 14422 6159 14462 6215
rect 10784 6137 14462 6159
rect 9816 6046 12150 6068
rect 9816 5990 9856 6046
rect 9912 5990 9936 6046
rect 9992 5990 10016 6046
rect 10072 5990 12150 6046
rect 9816 5968 12150 5990
rect 13101 6046 15430 6068
rect 13101 5990 15170 6046
rect 15226 5990 15250 6046
rect 15306 5990 15330 6046
rect 15386 5990 15430 6046
rect 13101 5968 15430 5990
rect -25759 5625 -25459 5637
rect -6617 5625 -6317 5637
rect -25759 5615 -22599 5625
rect -25759 5559 -25719 5615
rect -25663 5559 -25639 5615
rect -25583 5559 -25559 5615
rect -25503 5559 -22599 5615
rect -25759 5537 -22599 5559
rect -9476 5615 -6317 5625
rect -9476 5559 -6573 5615
rect -6517 5559 -6493 5615
rect -6437 5559 -6413 5615
rect -6357 5559 -6317 5615
rect -9476 5537 -6317 5559
rect -4750 5625 -4450 5636
rect 5753 5625 6053 5636
rect 6889 5625 7189 5636
rect 9816 5625 10116 5636
rect 15130 5625 15430 5636
rect 18395 5625 18695 5636
rect -4750 5614 -1553 5625
rect -4750 5558 -4706 5614
rect -4650 5558 -4626 5614
rect -4570 5558 -4546 5614
rect -4490 5558 -1553 5614
rect -4750 5536 -1553 5558
rect 2855 5614 8912 5625
rect 2855 5558 5793 5614
rect 5849 5558 5873 5614
rect 5929 5558 5953 5614
rect 6009 5558 6929 5614
rect 6985 5558 7009 5614
rect 7065 5558 7089 5614
rect 7145 5558 8912 5614
rect 2855 5536 8912 5558
rect 9816 5536 15430 5625
rect 15536 5614 18695 5625
rect 15536 5558 18435 5614
rect 18491 5558 18515 5614
rect 18571 5558 18595 5614
rect 18651 5558 18695 5614
rect 15536 5536 18695 5558
rect -4750 5305 -4450 5316
rect 5753 5305 6053 5316
rect 6889 5305 7189 5316
rect 10784 5305 11084 5316
rect 14162 5305 14462 5316
rect 18395 5305 18695 5316
rect -25759 5283 -22599 5305
rect -25759 5227 -25719 5283
rect -25663 5227 -25639 5283
rect -25583 5227 -25559 5283
rect -25503 5227 -22599 5283
rect -25759 5217 -22599 5227
rect -9476 5283 -6317 5305
rect -9476 5227 -6573 5283
rect -6517 5227 -6493 5283
rect -6437 5227 -6413 5283
rect -6357 5227 -6317 5283
rect -9476 5217 -6317 5227
rect -25759 5205 -25459 5217
rect -6617 5205 -6317 5217
rect -4750 5294 -1553 5305
rect -4750 5238 -4706 5294
rect -4650 5238 -4626 5294
rect -4570 5238 -4546 5294
rect -4490 5238 -1553 5294
rect -4750 5216 -1553 5238
rect 2855 5288 8912 5305
rect 2855 5232 5793 5288
rect 5849 5232 5873 5288
rect 5929 5232 5953 5288
rect 6009 5232 6929 5288
rect 6985 5232 7009 5288
rect 7065 5232 7089 5288
rect 7145 5232 8912 5288
rect 2855 5216 8912 5232
rect 10784 5216 14462 5305
rect 15536 5288 18695 5305
rect 15536 5232 18435 5288
rect 18491 5232 18515 5288
rect 18571 5232 18595 5288
rect 18651 5232 18695 5288
rect 15536 5216 18695 5232
rect 5753 5205 6053 5216
rect 6889 5205 7189 5216
rect 18395 5205 18695 5216
rect -24747 4852 -24551 4862
rect -24747 4800 -24738 4852
rect -24686 4800 -24674 4852
rect -24622 4800 -24610 4852
rect -24558 4800 -24551 4852
rect -24747 4792 -24551 4800
rect -16372 4852 -16176 4862
rect -16372 4800 -16363 4852
rect -16311 4800 -16299 4852
rect -16247 4800 -16235 4852
rect -16183 4800 -16176 4852
rect -16372 4792 -16176 4800
rect -15969 4852 -15773 4862
rect -15969 4800 -15960 4852
rect -15908 4800 -15896 4852
rect -15844 4800 -15832 4852
rect -15780 4800 -15773 4852
rect -15969 4792 -15773 4800
rect -7677 4852 -7481 4862
rect -7677 4800 -7668 4852
rect -7616 4800 -7604 4852
rect -7552 4800 -7540 4852
rect -7488 4800 -7481 4852
rect -7677 4792 -7481 4800
rect -3588 4852 -3392 4862
rect -3588 4800 -3579 4852
rect -3527 4800 -3515 4852
rect -3463 4800 -3451 4852
rect -3399 4800 -3392 4852
rect -3588 4792 -3392 4800
rect 4755 4852 4951 4862
rect 4755 4800 4764 4852
rect 4816 4800 4828 4852
rect 4880 4800 4892 4852
rect 4944 4800 4951 4852
rect 4755 4792 4951 4800
rect 8297 4851 8493 4861
rect 8297 4799 8306 4851
rect 8358 4799 8370 4851
rect 8422 4799 8434 4851
rect 8486 4799 8493 4851
rect 8297 4791 8493 4799
rect 16709 4851 16905 4861
rect 16709 4799 16718 4851
rect 16770 4799 16782 4851
rect 16834 4799 16846 4851
rect 16898 4799 16905 4851
rect 16709 4791 16905 4799
rect 10784 4695 14462 4717
rect 10784 4639 10828 4695
rect 10884 4639 10908 4695
rect 10964 4639 10988 4695
rect 11044 4639 14206 4695
rect 14262 4639 14286 4695
rect 14342 4639 14366 4695
rect 14422 4639 14462 4695
rect 10784 4617 14462 4639
rect 9816 4534 12150 4556
rect 9816 4478 9856 4534
rect 9912 4478 9936 4534
rect 9992 4478 10016 4534
rect 10072 4478 12150 4534
rect 9816 4456 12150 4478
rect 13101 4534 15430 4556
rect 13101 4478 15170 4534
rect 15226 4478 15250 4534
rect 15306 4478 15330 4534
rect 15386 4478 15430 4534
rect 13101 4456 15430 4478
rect -20704 4406 -20508 4416
rect -20704 4354 -20697 4406
rect -20645 4354 -20633 4406
rect -20581 4354 -20569 4406
rect -20517 4354 -20508 4406
rect -20704 4346 -20508 4354
rect -20383 4406 -20187 4416
rect -20383 4354 -20376 4406
rect -20324 4354 -20312 4406
rect -20260 4354 -20248 4406
rect -20196 4354 -20187 4406
rect -20383 4346 -20187 4354
rect -11998 4406 -11802 4416
rect -11998 4354 -11991 4406
rect -11939 4354 -11927 4406
rect -11875 4354 -11863 4406
rect -11811 4354 -11802 4406
rect -11998 4346 -11802 4354
rect -11659 4406 -11463 4416
rect -11659 4354 -11652 4406
rect -11600 4354 -11588 4406
rect -11536 4354 -11524 4406
rect -11472 4354 -11463 4406
rect -11659 4346 -11463 4354
rect 384 4406 580 4416
rect 384 4354 391 4406
rect 443 4354 455 4406
rect 507 4354 519 4406
rect 571 4354 580 4406
rect 384 4346 580 4354
rect 737 4406 933 4416
rect 737 4354 744 4406
rect 796 4354 808 4406
rect 860 4354 872 4406
rect 924 4354 933 4406
rect 737 4346 933 4354
rect 12383 4406 12579 4416
rect 12383 4354 12392 4406
rect 12444 4354 12456 4406
rect 12508 4354 12520 4406
rect 12572 4354 12579 4406
rect 12383 4346 12579 4354
rect 12690 4406 12886 4416
rect 12690 4354 12699 4406
rect 12751 4354 12763 4406
rect 12815 4354 12827 4406
rect 12879 4354 12886 4406
rect 12690 4346 12886 4354
rect -25759 3956 -22599 3978
rect -25759 3900 -25719 3956
rect -25663 3900 -25639 3956
rect -25583 3900 -25559 3956
rect -25503 3900 -22599 3956
rect -25759 3890 -22599 3900
rect -9476 3956 -6317 3978
rect -9476 3900 -6573 3956
rect -6517 3900 -6493 3956
rect -6437 3900 -6413 3956
rect -6357 3900 -6317 3956
rect -9476 3890 -6317 3900
rect -25759 3878 -25459 3890
rect -6617 3878 -6317 3890
rect -4750 3956 -1553 3978
rect -4750 3900 -4706 3956
rect -4650 3900 -4626 3956
rect -4570 3900 -4546 3956
rect -4490 3900 -1553 3956
rect -4750 3889 -1553 3900
rect 2855 3956 8912 3978
rect 2855 3900 5793 3956
rect 5849 3900 5873 3956
rect 5929 3900 5953 3956
rect 6009 3900 6929 3956
rect 6985 3900 7009 3956
rect 7065 3900 7089 3956
rect 7145 3900 8912 3956
rect 2855 3889 8912 3900
rect 10784 3889 14462 3978
rect 15536 3956 18695 3978
rect 15536 3900 18435 3956
rect 18491 3900 18515 3956
rect 18571 3900 18595 3956
rect 18651 3900 18695 3956
rect 15536 3889 18695 3900
rect -4750 3878 -4450 3889
rect 5753 3878 6053 3889
rect 6889 3878 7189 3889
rect 10784 3878 11084 3889
rect 14162 3878 14462 3889
rect 18395 3878 18695 3889
rect -25759 3636 -22599 3658
rect -25759 3580 -25719 3636
rect -25663 3580 -25639 3636
rect -25583 3580 -25559 3636
rect -25503 3580 -22599 3636
rect -25759 3570 -22599 3580
rect -9476 3636 -6317 3658
rect -9476 3580 -6573 3636
rect -6517 3580 -6493 3636
rect -6437 3580 -6413 3636
rect -6357 3580 -6317 3636
rect -9476 3570 -6317 3580
rect -25759 3558 -25459 3570
rect -6617 3558 -6317 3570
rect -4750 3636 -1553 3658
rect -4750 3580 -4706 3636
rect -4650 3580 -4626 3636
rect -4570 3580 -4546 3636
rect -4490 3580 -1553 3636
rect -4750 3569 -1553 3580
rect 2855 3636 8912 3658
rect 2855 3580 5793 3636
rect 5849 3580 5873 3636
rect 5929 3580 5953 3636
rect 6009 3580 6929 3636
rect 6985 3580 7009 3636
rect 7065 3580 7089 3636
rect 7145 3580 8912 3636
rect 2855 3569 8912 3580
rect 9816 3569 15430 3658
rect 15536 3636 18695 3658
rect 15536 3580 18435 3636
rect 18491 3580 18515 3636
rect 18571 3580 18595 3636
rect 18651 3580 18695 3636
rect 15536 3569 18695 3580
rect -4750 3558 -4450 3569
rect 5753 3558 6053 3569
rect 6889 3558 7189 3569
rect 9816 3558 10116 3569
rect 15130 3558 15430 3569
rect 18395 3558 18695 3569
rect -24756 2885 -24560 2895
rect -24756 2833 -24747 2885
rect -24695 2833 -24683 2885
rect -24631 2833 -24619 2885
rect -24567 2833 -24560 2885
rect -24756 2825 -24560 2833
rect -16380 2885 -16184 2895
rect -16380 2833 -16371 2885
rect -16319 2833 -16307 2885
rect -16255 2833 -16243 2885
rect -16191 2833 -16184 2885
rect -16380 2825 -16184 2833
rect -15977 2885 -15781 2895
rect -15977 2833 -15968 2885
rect -15916 2833 -15904 2885
rect -15852 2833 -15840 2885
rect -15788 2833 -15781 2885
rect -15977 2825 -15781 2833
rect -7686 2885 -7490 2895
rect -7686 2833 -7677 2885
rect -7625 2833 -7613 2885
rect -7561 2833 -7549 2885
rect -7497 2833 -7490 2885
rect -7686 2825 -7490 2833
rect -3597 2885 -3401 2895
rect -3597 2833 -3588 2885
rect -3536 2833 -3524 2885
rect -3472 2833 -3460 2885
rect -3408 2833 -3401 2885
rect -3597 2825 -3401 2833
rect 4746 2885 4942 2895
rect 4746 2833 4755 2885
rect 4807 2833 4819 2885
rect 4871 2833 4883 2885
rect 4935 2833 4942 2885
rect 4746 2825 4942 2833
rect 8324 2885 8520 2895
rect 8324 2833 8333 2885
rect 8385 2833 8397 2885
rect 8449 2833 8461 2885
rect 8513 2833 8520 2885
rect 8324 2825 8520 2833
rect 16679 2885 16979 2895
rect 16679 2833 16744 2885
rect 16796 2833 16808 2885
rect 16860 2833 16872 2885
rect 16924 2833 16979 2885
rect 16679 2795 16979 2833
rect -20686 2716 -20490 2726
rect -20686 2664 -20679 2716
rect -20627 2664 -20615 2716
rect -20563 2664 -20551 2716
rect -20499 2664 -20490 2716
rect -20686 2656 -20490 2664
rect -20365 2716 -20169 2726
rect -20365 2664 -20358 2716
rect -20306 2664 -20294 2716
rect -20242 2664 -20230 2716
rect -20178 2664 -20169 2716
rect -20365 2656 -20169 2664
rect -11980 2716 -11784 2726
rect -11980 2664 -11973 2716
rect -11921 2664 -11909 2716
rect -11857 2664 -11845 2716
rect -11793 2664 -11784 2716
rect -11980 2656 -11784 2664
rect -11641 2716 -11445 2726
rect -11641 2664 -11634 2716
rect -11582 2664 -11570 2716
rect -11518 2664 -11506 2716
rect -11454 2664 -11445 2716
rect -11641 2656 -11445 2664
rect 402 2716 598 2726
rect 402 2664 409 2716
rect 461 2664 473 2716
rect 525 2664 537 2716
rect 589 2664 598 2716
rect 402 2656 598 2664
rect 755 2716 951 2726
rect 755 2664 762 2716
rect 814 2664 826 2716
rect 878 2664 890 2716
rect 942 2664 951 2716
rect 755 2656 951 2664
rect 12367 2716 12563 2726
rect 12367 2664 12376 2716
rect 12428 2664 12440 2716
rect 12492 2664 12504 2716
rect 12556 2664 12563 2716
rect 12367 2656 12563 2664
rect 12664 2716 12860 2726
rect 12664 2664 12673 2716
rect 12725 2664 12737 2716
rect 12789 2664 12801 2716
rect 12853 2664 12860 2716
rect 12664 2656 12860 2664
rect -11284 2497 -10275 2519
rect -11284 2441 -11240 2497
rect -11184 2441 -11160 2497
rect -11104 2441 -11080 2497
rect -11024 2441 -10531 2497
rect -10475 2441 -10451 2497
rect -10395 2441 -10371 2497
rect -10315 2441 -10275 2497
rect -11284 2397 -10275 2441
rect -11284 2341 -11240 2397
rect -11184 2341 -11160 2397
rect -11104 2341 -11080 2397
rect -11024 2341 -10531 2397
rect -10475 2341 -10451 2397
rect -10395 2341 -10371 2397
rect -10315 2341 -10275 2397
rect -11284 2319 -10275 2341
rect -46 2414 1404 2436
rect -46 2358 -6 2414
rect 50 2358 74 2414
rect 130 2358 154 2414
rect 210 2358 562 2414
rect 618 2358 642 2414
rect 698 2358 722 2414
rect 778 2358 1144 2414
rect 1200 2358 1224 2414
rect 1280 2358 1304 2414
rect 1360 2358 1404 2414
rect -46 2314 1404 2358
rect -46 2258 -6 2314
rect 50 2258 74 2314
rect 130 2258 154 2314
rect 210 2258 562 2314
rect 618 2258 642 2314
rect 698 2258 722 2314
rect 778 2258 1144 2314
rect 1200 2258 1224 2314
rect 1280 2258 1304 2314
rect 1360 2258 1404 2314
rect -46 2214 1404 2258
rect -24359 2140 -6931 2162
rect -24359 2084 -24315 2140
rect -24259 2084 -24235 2140
rect -24179 2084 -24155 2140
rect -24099 2084 -16749 2140
rect -16693 2084 -16669 2140
rect -16613 2084 -16589 2140
rect -16533 2084 -15598 2140
rect -15542 2084 -15518 2140
rect -15462 2084 -15438 2140
rect -15382 2084 -11400 2140
rect -11344 2084 -11320 2140
rect -11264 2084 -11240 2140
rect -11184 2084 -8032 2140
rect -7976 2084 -7952 2140
rect -7896 2084 -7872 2140
rect -7816 2084 -7187 2140
rect -7131 2084 -7107 2140
rect -7051 2084 -7027 2140
rect -6971 2084 -6931 2140
rect -24359 2040 -6931 2084
rect -24359 1984 -24315 2040
rect -24259 1984 -24235 2040
rect -24179 1984 -24155 2040
rect -24099 1984 -16749 2040
rect -16693 1984 -16669 2040
rect -16613 1984 -16589 2040
rect -16533 1984 -15598 2040
rect -15542 1984 -15518 2040
rect -15462 1984 -15438 2040
rect -15382 1984 -11400 2040
rect -11344 1984 -11320 2040
rect -11264 1984 -11240 2040
rect -11184 1984 -8032 2040
rect -7976 1984 -7952 2040
rect -7896 1984 -7872 2040
rect -7816 1984 -7187 2040
rect -7131 1984 -7107 2040
rect -7051 1984 -7027 2040
rect -6971 1984 -6931 2040
rect -46 2158 -6 2214
rect 50 2158 74 2214
rect 130 2158 154 2214
rect 210 2158 562 2214
rect 618 2158 642 2214
rect 698 2158 722 2214
rect 778 2158 1144 2214
rect 1200 2158 1224 2214
rect 1280 2158 1304 2214
rect 1360 2158 1404 2214
rect -46 2114 1404 2158
rect -46 2058 -6 2114
rect 50 2058 74 2114
rect 130 2058 154 2114
rect 210 2058 562 2114
rect 618 2058 642 2114
rect 698 2058 722 2114
rect 778 2058 1144 2114
rect 1200 2058 1224 2114
rect 1280 2058 1304 2114
rect 1360 2058 1404 2114
rect -46 2036 1404 2058
rect -24359 1962 -6931 1984
rect -25356 1791 -10275 1813
rect -25356 1735 -25310 1791
rect -25254 1735 -25230 1791
rect -25174 1735 -25150 1791
rect -25094 1735 -21107 1791
rect -21051 1735 -21027 1791
rect -20971 1735 -20947 1791
rect -20891 1735 -19957 1791
rect -19901 1735 -19877 1791
rect -19821 1735 -19797 1791
rect -19741 1735 -16899 1791
rect -16843 1735 -16819 1791
rect -16763 1735 -16739 1791
rect -16683 1735 -12390 1791
rect -12334 1735 -12310 1791
rect -12254 1735 -12230 1791
rect -12174 1735 -10531 1791
rect -10475 1735 -10451 1791
rect -10395 1735 -10371 1791
rect -10315 1735 -10275 1791
rect -25356 1691 -10275 1735
rect -25356 1635 -25310 1691
rect -25254 1635 -25230 1691
rect -25174 1635 -25150 1691
rect -25094 1635 -21107 1691
rect -21051 1635 -21027 1691
rect -20971 1635 -20947 1691
rect -20891 1635 -19957 1691
rect -19901 1635 -19877 1691
rect -19821 1635 -19797 1691
rect -19741 1635 -16899 1691
rect -16843 1635 -16819 1691
rect -16763 1635 -16739 1691
rect -16683 1635 -12390 1691
rect -12334 1635 -12310 1691
rect -12254 1635 -12230 1691
rect -12174 1635 -10531 1691
rect -10475 1635 -10451 1691
rect -10395 1635 -10371 1691
rect -10315 1635 -10275 1691
rect -25356 1613 -10275 1635
rect -3676 1808 5035 1830
rect -3676 1752 -3636 1808
rect -3580 1752 -3556 1808
rect -3500 1752 -3476 1808
rect -3420 1752 -3214 1808
rect -3158 1752 -3134 1808
rect -3078 1752 -3054 1808
rect -2998 1752 4352 1808
rect 4408 1752 4432 1808
rect 4488 1752 4512 1808
rect 4568 1752 4775 1808
rect 4831 1752 4855 1808
rect 4911 1752 4935 1808
rect 4991 1752 5035 1808
rect -3676 1708 5035 1752
rect -3676 1652 -3636 1708
rect -3580 1652 -3556 1708
rect -3500 1652 -3476 1708
rect -3420 1652 -3214 1708
rect -3158 1652 -3134 1708
rect -3078 1652 -3054 1708
rect -2998 1652 4352 1708
rect 4408 1652 4432 1708
rect 4488 1652 4512 1708
rect 4568 1652 4775 1708
rect 4831 1652 4855 1708
rect 4911 1652 4935 1708
rect 4991 1652 5035 1708
rect -3676 1608 5035 1652
rect -3676 1552 -3636 1608
rect -3580 1552 -3556 1608
rect -3500 1552 -3476 1608
rect -3420 1552 -3214 1608
rect -3158 1552 -3134 1608
rect -3078 1552 -3054 1608
rect -2998 1552 4352 1608
rect 4408 1552 4432 1608
rect 4488 1552 4512 1608
rect 4568 1552 4775 1608
rect 4831 1552 4855 1608
rect 4911 1552 4935 1608
rect 4991 1552 5035 1608
rect -3676 1508 5035 1552
rect -3676 1452 -3636 1508
rect -3580 1452 -3556 1508
rect -3500 1452 -3476 1508
rect -3420 1452 -3214 1508
rect -3158 1452 -3134 1508
rect -3078 1452 -3054 1508
rect -2998 1452 4352 1508
rect 4408 1452 4432 1508
rect 4488 1452 4512 1508
rect 4568 1452 4775 1508
rect 4831 1452 4855 1508
rect 4911 1452 4935 1508
rect 4991 1452 5035 1508
rect -3676 1430 5035 1452
rect 5753 1331 7189 1353
rect 5753 1275 5793 1331
rect 5849 1275 5873 1331
rect 5929 1275 5953 1331
rect 6009 1275 6929 1331
rect 6985 1275 7009 1331
rect 7065 1275 7089 1331
rect 7145 1275 7189 1331
rect 5753 1231 7189 1275
rect 5753 1175 5793 1231
rect 5849 1175 5873 1231
rect 5929 1175 5953 1231
rect 6009 1175 6929 1231
rect 6985 1175 7009 1231
rect 7065 1175 7089 1231
rect 7145 1175 7189 1231
rect 5753 1131 7189 1175
rect 12389 1209 12585 1217
rect 12389 1157 12398 1209
rect 12450 1157 12462 1209
rect 12514 1157 12526 1209
rect 12578 1157 12585 1209
rect 12389 1147 12585 1157
rect 12680 1209 12876 1217
rect 12680 1157 12689 1209
rect 12741 1157 12753 1209
rect 12805 1157 12817 1209
rect 12869 1157 12876 1209
rect 12680 1147 12876 1157
rect 5753 1075 5793 1131
rect 5849 1075 5873 1131
rect 5929 1075 5953 1131
rect 6009 1075 6929 1131
rect 6985 1075 7009 1131
rect 7065 1075 7089 1131
rect 7145 1075 7189 1131
rect 5753 1031 7189 1075
rect 5753 975 5793 1031
rect 5849 975 5873 1031
rect 5929 975 5953 1031
rect 6009 975 6929 1031
rect 6985 975 7009 1031
rect 7065 975 7089 1031
rect 7145 975 7189 1031
rect 8324 1040 8520 1048
rect 8324 988 8333 1040
rect 8385 988 8397 1040
rect 8449 988 8461 1040
rect 8513 988 8520 1040
rect 8324 978 8520 988
rect 16736 1040 16932 1048
rect 16736 988 16745 1040
rect 16797 988 16809 1040
rect 16861 988 16873 1040
rect 16925 988 16932 1040
rect 16736 978 16932 988
rect 5753 953 7189 975
rect -26532 304 -26232 316
rect -6105 304 -5805 316
rect -26532 294 -23206 304
rect -26532 238 -26492 294
rect -26436 238 -26412 294
rect -26356 238 -26332 294
rect -26276 238 -23206 294
rect -26532 216 -23206 238
rect -9131 294 -5805 304
rect -9131 238 -6061 294
rect -6005 238 -5981 294
rect -5925 238 -5901 294
rect -5845 238 -5805 294
rect -9131 216 -5805 238
rect -4750 304 -4450 316
rect 5753 304 6053 316
rect -4750 294 -1553 304
rect -4750 238 -4706 294
rect -4650 238 -4626 294
rect -4570 238 -4546 294
rect -4490 238 -1553 294
rect -4750 216 -1553 238
rect 2855 294 6053 304
rect 2855 238 5793 294
rect 5849 238 5873 294
rect 5929 238 5953 294
rect 6009 238 6053 294
rect 2855 216 6053 238
rect 9816 304 10116 316
rect 15130 304 15430 316
rect 9816 216 15430 304
rect -27032 -16 -26732 -5
rect -5606 -16 -5306 -5
rect 10784 -16 11084 -5
rect 14162 -16 14462 -5
rect -27032 -27 -23863 -16
rect -27032 -83 -26992 -27
rect -26936 -83 -26912 -27
rect -26856 -83 -26832 -27
rect -26776 -83 -23863 -27
rect -27032 -105 -23863 -83
rect -8474 -27 -5306 -16
rect -8474 -83 -5562 -27
rect -5506 -83 -5482 -27
rect -5426 -83 -5402 -27
rect -5346 -83 -5306 -27
rect -8474 -105 -5306 -83
rect -4712 -105 -1553 -16
rect 2855 -105 6015 -16
rect 10784 -105 14462 -16
rect 12376 -481 12572 -473
rect 12376 -533 12385 -481
rect 12437 -533 12449 -481
rect 12501 -533 12513 -481
rect 12565 -533 12572 -481
rect 12376 -543 12572 -533
rect 12661 -481 12857 -473
rect 12661 -533 12670 -481
rect 12722 -533 12734 -481
rect 12786 -533 12798 -481
rect 12850 -533 12857 -481
rect 12661 -543 12857 -533
rect 9816 -604 12150 -582
rect 9816 -660 9856 -604
rect 9912 -660 9936 -604
rect 9992 -660 10016 -604
rect 10072 -660 12150 -604
rect 9816 -682 12150 -660
rect 13101 -604 15430 -582
rect 13101 -660 15170 -604
rect 15226 -660 15250 -604
rect 15306 -660 15330 -604
rect 15386 -660 15430 -604
rect 13101 -682 15430 -660
rect 10784 -765 14468 -743
rect 10784 -821 10828 -765
rect 10884 -821 10908 -765
rect 10964 -821 10988 -765
rect 11044 -821 14206 -765
rect 14262 -821 14286 -765
rect 14342 -821 14366 -765
rect 14422 -821 14468 -765
rect 10784 -843 14468 -821
rect 8311 -926 8507 -918
rect 8311 -978 8320 -926
rect 8372 -978 8384 -926
rect 8436 -978 8448 -926
rect 8500 -978 8507 -926
rect 8311 -988 8507 -978
rect 16722 -926 16918 -918
rect 16722 -978 16731 -926
rect 16783 -978 16795 -926
rect 16847 -978 16859 -926
rect 16911 -978 16918 -926
rect 16722 -988 16918 -978
rect -27032 -1365 -23863 -1343
rect -27032 -1421 -26992 -1365
rect -26936 -1421 -26912 -1365
rect -26856 -1421 -26832 -1365
rect -26776 -1421 -23863 -1365
rect -27032 -1431 -23863 -1421
rect -8474 -1365 -5306 -1343
rect -8474 -1421 -5562 -1365
rect -5506 -1421 -5482 -1365
rect -5426 -1421 -5402 -1365
rect -5346 -1421 -5306 -1365
rect -8474 -1431 -5306 -1421
rect -4712 -1431 -1553 -1343
rect 2855 -1431 6015 -1343
rect 10784 -1431 14462 -1343
rect -27032 -1443 -26732 -1431
rect -5606 -1443 -5306 -1431
rect 10784 -1443 11084 -1431
rect 14162 -1443 14462 -1431
rect -26532 -1685 -23206 -1663
rect -26532 -1741 -26492 -1685
rect -26436 -1741 -26412 -1685
rect -26356 -1741 -26332 -1685
rect -26276 -1741 -23206 -1685
rect -26532 -1752 -23206 -1741
rect -9131 -1685 -5805 -1663
rect -9131 -1741 -6061 -1685
rect -6005 -1741 -5981 -1685
rect -5925 -1741 -5901 -1685
rect -5845 -1741 -5805 -1685
rect -9131 -1752 -5805 -1741
rect -26532 -1763 -26232 -1752
rect -6105 -1763 -5805 -1752
rect -4750 -1685 -1553 -1663
rect -4750 -1741 -4706 -1685
rect -4650 -1741 -4626 -1685
rect -4570 -1741 -4546 -1685
rect -4490 -1741 -1553 -1685
rect -4750 -1752 -1553 -1741
rect 2855 -1685 6053 -1663
rect 2855 -1741 5793 -1685
rect 5849 -1741 5873 -1685
rect 5929 -1741 5953 -1685
rect 6009 -1741 6053 -1685
rect 2855 -1752 6053 -1741
rect -4750 -1763 -4450 -1752
rect 5753 -1763 6053 -1752
rect 9816 -1752 15430 -1663
rect 9816 -1763 10116 -1752
rect 15130 -1763 15430 -1752
rect 9816 -2117 12150 -2095
rect 9816 -2173 9856 -2117
rect 9912 -2173 9936 -2117
rect 9992 -2173 10016 -2117
rect 10072 -2173 12150 -2117
rect 9816 -2195 12150 -2173
rect 13101 -2117 15430 -2095
rect 13101 -2173 15170 -2117
rect 15226 -2173 15250 -2117
rect 15306 -2173 15330 -2117
rect 15386 -2173 15430 -2117
rect 13101 -2195 15430 -2173
rect 10784 -2285 14462 -2263
rect 10784 -2341 10828 -2285
rect 10884 -2341 10908 -2285
rect 10964 -2341 10988 -2285
rect 11044 -2341 14206 -2285
rect 14262 -2341 14286 -2285
rect 14342 -2341 14366 -2285
rect 14422 -2341 14462 -2285
rect 10784 -2363 14462 -2341
rect 8314 -2436 8510 -2426
rect 8314 -2488 8323 -2436
rect 8375 -2488 8387 -2436
rect 8439 -2488 8451 -2436
rect 8503 -2488 8510 -2436
rect 8314 -2496 8510 -2488
rect 16725 -2436 16921 -2426
rect 16725 -2488 16734 -2436
rect 16786 -2488 16798 -2436
rect 16850 -2488 16862 -2436
rect 16914 -2488 16921 -2436
rect 16725 -2496 16921 -2488
rect 12375 -2605 12571 -2595
rect 12375 -2657 12384 -2605
rect 12436 -2657 12448 -2605
rect 12500 -2657 12512 -2605
rect 12564 -2657 12571 -2605
rect 12375 -2665 12571 -2657
rect 12676 -2605 12872 -2595
rect 12676 -2657 12685 -2605
rect 12737 -2657 12749 -2605
rect 12801 -2657 12813 -2605
rect 12865 -2657 12872 -2605
rect 12676 -2665 12872 -2657
rect 12354 -3664 12550 -3656
rect 12354 -3716 12363 -3664
rect 12415 -3716 12427 -3664
rect 12479 -3716 12491 -3664
rect 12543 -3716 12550 -3664
rect 12354 -3726 12550 -3716
rect 12665 -3664 12861 -3656
rect 12665 -3716 12674 -3664
rect 12726 -3716 12738 -3664
rect 12790 -3716 12802 -3664
rect 12854 -3716 12861 -3664
rect 12665 -3726 12861 -3716
rect 8310 -3833 8506 -3825
rect 8310 -3885 8319 -3833
rect 8371 -3885 8383 -3833
rect 8435 -3885 8447 -3833
rect 8499 -3885 8506 -3833
rect 8310 -3895 8506 -3885
rect 16721 -3833 16917 -3825
rect 16721 -3885 16730 -3833
rect 16782 -3885 16794 -3833
rect 16846 -3885 16858 -3833
rect 16910 -3885 16917 -3833
rect 16721 -3895 16917 -3885
rect 10784 -3979 14462 -3957
rect 10784 -4035 10828 -3979
rect 10884 -4035 10908 -3979
rect 10964 -4035 10988 -3979
rect 11044 -4035 14206 -3979
rect 14262 -4035 14286 -3979
rect 14342 -4035 14366 -3979
rect 14422 -4035 14462 -3979
rect 10784 -4057 14462 -4035
rect 9816 -4148 12150 -4126
rect 9816 -4204 9856 -4148
rect 9912 -4204 9936 -4148
rect 9992 -4204 10016 -4148
rect 10072 -4204 12150 -4148
rect 9816 -4226 12150 -4204
rect 13101 -4148 15430 -4126
rect 13101 -4204 15170 -4148
rect 15226 -4204 15250 -4148
rect 15306 -4204 15330 -4148
rect 15386 -4204 15430 -4148
rect 13101 -4226 15430 -4204
rect -26532 -4569 -26232 -4558
rect -6105 -4569 -5805 -4558
rect -26532 -4580 -23206 -4569
rect -26532 -4636 -26492 -4580
rect -26436 -4636 -26412 -4580
rect -26356 -4636 -26332 -4580
rect -26276 -4636 -23206 -4580
rect -26532 -4658 -23206 -4636
rect -9131 -4580 -5805 -4569
rect -9131 -4636 -6061 -4580
rect -6005 -4636 -5981 -4580
rect -5925 -4636 -5901 -4580
rect -5845 -4636 -5805 -4580
rect -9131 -4658 -5805 -4636
rect -4750 -4569 -4450 -4558
rect 5753 -4569 6053 -4558
rect -4750 -4580 -1553 -4569
rect -4750 -4636 -4706 -4580
rect -4650 -4636 -4626 -4580
rect -4570 -4636 -4546 -4580
rect -4490 -4636 -1553 -4580
rect -4750 -4658 -1553 -4636
rect 2855 -4580 6053 -4569
rect 2855 -4636 5793 -4580
rect 5849 -4636 5873 -4580
rect 5929 -4636 5953 -4580
rect 6009 -4636 6053 -4580
rect 2855 -4658 6053 -4636
rect 9816 -4569 10116 -4558
rect 15130 -4569 15430 -4558
rect 9816 -4658 15430 -4569
rect -27032 -4889 -26732 -4878
rect -5606 -4889 -5306 -4878
rect -27032 -4900 -23863 -4889
rect -27032 -4956 -26992 -4900
rect -26936 -4956 -26912 -4900
rect -26856 -4956 -26832 -4900
rect -26776 -4956 -23863 -4900
rect -27032 -4978 -23863 -4956
rect -8474 -4900 -5306 -4889
rect -8474 -4956 -5562 -4900
rect -5506 -4956 -5482 -4900
rect -5426 -4956 -5402 -4900
rect -5346 -4956 -5306 -4900
rect -8474 -4978 -5306 -4956
rect -4750 -4889 -4450 -4878
rect 5753 -4889 6053 -4878
rect -4750 -4900 -1553 -4889
rect -4750 -4956 -4706 -4900
rect -4650 -4956 -4626 -4900
rect -4570 -4956 -4546 -4900
rect -4490 -4956 -1553 -4900
rect -4750 -4978 -1553 -4956
rect 2855 -4900 6053 -4889
rect 2855 -4956 5793 -4900
rect 5849 -4956 5873 -4900
rect 5929 -4956 5953 -4900
rect 6009 -4956 6053 -4900
rect 2855 -4978 6053 -4956
rect 10784 -4889 11084 -4878
rect 14162 -4889 14462 -4878
rect 10784 -4978 14462 -4889
rect 8297 -5343 8493 -5333
rect 8297 -5395 8306 -5343
rect 8358 -5395 8370 -5343
rect 8422 -5395 8434 -5343
rect 8486 -5395 8493 -5343
rect 8297 -5403 8493 -5395
rect 16709 -5343 16905 -5333
rect 16709 -5395 16718 -5343
rect 16770 -5395 16782 -5343
rect 16834 -5395 16846 -5343
rect 16898 -5395 16905 -5343
rect 16709 -5403 16905 -5395
rect 10784 -5499 14462 -5477
rect 10784 -5555 10828 -5499
rect 10884 -5555 10908 -5499
rect 10964 -5555 10988 -5499
rect 11044 -5555 14206 -5499
rect 14262 -5555 14286 -5499
rect 14342 -5555 14366 -5499
rect 14422 -5555 14462 -5499
rect 10784 -5577 14462 -5555
rect 9816 -5660 12150 -5638
rect 9816 -5716 9856 -5660
rect 9912 -5716 9936 -5660
rect 9992 -5716 10016 -5660
rect 10072 -5716 12150 -5660
rect 9816 -5738 12150 -5716
rect 13101 -5660 15430 -5638
rect 13101 -5716 15170 -5660
rect 15226 -5716 15250 -5660
rect 15306 -5716 15330 -5660
rect 15386 -5716 15430 -5660
rect 13101 -5738 15430 -5716
rect 12383 -5788 12579 -5778
rect 12383 -5840 12392 -5788
rect 12444 -5840 12456 -5788
rect 12508 -5840 12520 -5788
rect 12572 -5840 12579 -5788
rect 12383 -5848 12579 -5840
rect 12690 -5788 12886 -5778
rect 12690 -5840 12699 -5788
rect 12751 -5840 12763 -5788
rect 12815 -5840 12827 -5788
rect 12879 -5840 12886 -5788
rect 12690 -5848 12886 -5840
rect -27032 -6238 -23863 -6216
rect -27032 -6294 -26992 -6238
rect -26936 -6294 -26912 -6238
rect -26856 -6294 -26832 -6238
rect -26776 -6294 -23863 -6238
rect -27032 -6305 -23863 -6294
rect -8474 -6238 -5306 -6216
rect -8474 -6294 -5562 -6238
rect -5506 -6294 -5482 -6238
rect -5426 -6294 -5402 -6238
rect -5346 -6294 -5306 -6238
rect -8474 -6305 -5306 -6294
rect -27032 -6316 -26732 -6305
rect -5606 -6316 -5306 -6305
rect -4750 -6238 -1553 -6216
rect -4750 -6294 -4706 -6238
rect -4650 -6294 -4626 -6238
rect -4570 -6294 -4546 -6238
rect -4490 -6294 -1553 -6238
rect -4750 -6305 -1553 -6294
rect 2855 -6238 6053 -6216
rect 2855 -6294 5793 -6238
rect 5849 -6294 5873 -6238
rect 5929 -6294 5953 -6238
rect 6009 -6294 6053 -6238
rect 2855 -6305 6053 -6294
rect -4750 -6316 -4450 -6305
rect 5753 -6316 6053 -6305
rect 10784 -6305 14462 -6216
rect 10784 -6316 11084 -6305
rect 14162 -6316 14462 -6305
rect -26532 -6558 -23206 -6536
rect -26532 -6614 -26492 -6558
rect -26436 -6614 -26412 -6558
rect -26356 -6614 -26332 -6558
rect -26276 -6614 -23206 -6558
rect -26532 -6625 -23206 -6614
rect -9131 -6558 -5805 -6536
rect -9131 -6614 -6061 -6558
rect -6005 -6614 -5981 -6558
rect -5925 -6614 -5901 -6558
rect -5845 -6614 -5805 -6558
rect -9131 -6625 -5805 -6614
rect -26532 -6636 -26232 -6625
rect -6105 -6636 -5805 -6625
rect -4750 -6558 -1553 -6536
rect -4750 -6614 -4706 -6558
rect -4650 -6614 -4626 -6558
rect -4570 -6614 -4546 -6558
rect -4490 -6614 -1553 -6558
rect -4750 -6625 -1553 -6614
rect 2855 -6558 6053 -6536
rect 2855 -6614 5793 -6558
rect 5849 -6614 5873 -6558
rect 5929 -6614 5953 -6558
rect 6009 -6614 6053 -6558
rect 2855 -6625 6053 -6614
rect -4750 -6636 -4450 -6625
rect 5753 -6636 6053 -6625
rect 9816 -6625 15430 -6536
rect 9816 -6636 10116 -6625
rect 15130 -6636 15430 -6625
rect 8324 -7309 8520 -7299
rect 8324 -7361 8333 -7309
rect 8385 -7361 8397 -7309
rect 8449 -7361 8461 -7309
rect 8513 -7361 8520 -7309
rect 8324 -7369 8520 -7361
rect 16679 -7309 16979 -7299
rect 16679 -7361 16744 -7309
rect 16796 -7361 16808 -7309
rect 16860 -7361 16872 -7309
rect 16924 -7361 16979 -7309
rect 16679 -7399 16979 -7361
rect 12367 -7478 12563 -7468
rect 12367 -7530 12376 -7478
rect 12428 -7530 12440 -7478
rect 12492 -7530 12504 -7478
rect 12556 -7530 12563 -7478
rect 12367 -7538 12563 -7530
rect 12664 -7478 12860 -7468
rect 12664 -7530 12673 -7478
rect 12725 -7530 12737 -7478
rect 12789 -7530 12801 -7478
rect 12853 -7530 12860 -7478
rect 12664 -7538 12860 -7530
rect 11645 -7780 13348 -7758
rect 11645 -7836 11796 -7780
rect 11852 -7836 11876 -7780
rect 11932 -7836 11956 -7780
rect 12012 -7836 13088 -7780
rect 13144 -7836 13168 -7780
rect 13224 -7836 13248 -7780
rect 13304 -7836 13348 -7780
rect 11645 -7880 13348 -7836
rect 11645 -7936 11796 -7880
rect 11852 -7936 11876 -7880
rect 11932 -7936 11956 -7880
rect 12012 -7936 13088 -7880
rect 13144 -7936 13168 -7880
rect 13224 -7936 13248 -7880
rect 13304 -7936 13348 -7880
rect 11645 -7980 13348 -7936
rect -24932 -8018 -10561 -7996
rect -24932 -8074 -24892 -8018
rect -24836 -8074 -24812 -8018
rect -24756 -8074 -24732 -8018
rect -24676 -8074 -17326 -8018
rect -17270 -8074 -17246 -8018
rect -17190 -8074 -17166 -8018
rect -17110 -8074 -11972 -8018
rect -11916 -8074 -11892 -8018
rect -11836 -8074 -11812 -8018
rect -11756 -8074 -10821 -8018
rect -10765 -8074 -10741 -8018
rect -10685 -8074 -10661 -8018
rect -10605 -8074 -10561 -8018
rect -24932 -8118 -10561 -8074
rect -24932 -8174 -24892 -8118
rect -24836 -8174 -24812 -8118
rect -24756 -8174 -24732 -8118
rect -24676 -8174 -17326 -8118
rect -17270 -8174 -17246 -8118
rect -17190 -8174 -17166 -8118
rect -17110 -8174 -11972 -8118
rect -11916 -8174 -11892 -8118
rect -11836 -8174 -11812 -8118
rect -11756 -8174 -10821 -8118
rect -10765 -8174 -10741 -8118
rect -10685 -8174 -10661 -8118
rect -10605 -8174 -10561 -8118
rect 11645 -8036 11796 -7980
rect 11852 -8036 11876 -7980
rect 11932 -8036 11956 -7980
rect 12012 -8036 13088 -7980
rect 13144 -8036 13168 -7980
rect 13224 -8036 13248 -7980
rect 13304 -8036 13348 -7980
rect 11645 -8080 13348 -8036
rect 11645 -8136 11796 -8080
rect 11852 -8136 11876 -8080
rect 11932 -8136 11956 -8080
rect 12012 -8136 13088 -8080
rect 13144 -8136 13168 -8080
rect 13224 -8136 13248 -8080
rect 13304 -8136 13348 -8080
rect 11645 -8158 13348 -8136
rect -24932 -8218 -10561 -8174
rect -24932 -8274 -24892 -8218
rect -24836 -8274 -24812 -8218
rect -24756 -8274 -24732 -8218
rect -24676 -8274 -17326 -8218
rect -17270 -8274 -17246 -8218
rect -17190 -8274 -17166 -8218
rect -17110 -8274 -11972 -8218
rect -11916 -8274 -11892 -8218
rect -11836 -8274 -11812 -8218
rect -11756 -8274 -10821 -8218
rect -10765 -8274 -10741 -8218
rect -10685 -8274 -10661 -8218
rect -10605 -8274 -10561 -8218
rect -24932 -8318 -10561 -8274
rect -24932 -8374 -24892 -8318
rect -24836 -8374 -24812 -8318
rect -24756 -8374 -24732 -8318
rect -24676 -8374 -17326 -8318
rect -17270 -8374 -17246 -8318
rect -17190 -8374 -17166 -8318
rect -17110 -8374 -11972 -8318
rect -11916 -8374 -11892 -8318
rect -11836 -8374 -11812 -8318
rect -11756 -8374 -10821 -8318
rect -10765 -8374 -10741 -8318
rect -10685 -8374 -10661 -8318
rect -10605 -8374 -10561 -8318
rect -24932 -8396 -10561 -8374
rect -46 -8349 8265 -8327
rect -46 -8405 -6 -8349
rect 50 -8405 74 -8349
rect 130 -8405 154 -8349
rect 210 -8405 1144 -8349
rect 1200 -8405 1224 -8349
rect 1280 -8405 1304 -8349
rect 1360 -8405 1990 -8349
rect 2046 -8405 2070 -8349
rect 2126 -8405 2150 -8349
rect 2206 -8405 8265 -8349
rect -46 -8449 8265 -8405
rect -46 -8505 -6 -8449
rect 50 -8505 74 -8449
rect 130 -8505 154 -8449
rect 210 -8505 1144 -8449
rect 1200 -8505 1224 -8449
rect 1280 -8505 1304 -8449
rect 1360 -8505 1990 -8449
rect 2046 -8505 2070 -8449
rect 2126 -8505 2150 -8449
rect 2206 -8505 8265 -8449
rect -46 -8549 8265 -8505
rect -46 -8605 -6 -8549
rect 50 -8605 74 -8549
rect 130 -8605 154 -8549
rect 210 -8605 1144 -8549
rect 1200 -8605 1224 -8549
rect 1280 -8605 1304 -8549
rect 1360 -8605 1990 -8549
rect 2046 -8605 2070 -8549
rect 2126 -8605 2150 -8549
rect 2206 -8605 8265 -8549
rect -46 -8649 8265 -8605
rect -46 -8705 -6 -8649
rect 50 -8705 74 -8649
rect 130 -8705 154 -8649
rect 210 -8705 1144 -8649
rect 1200 -8705 1224 -8649
rect 1280 -8705 1304 -8649
rect 1360 -8705 1990 -8649
rect 2046 -8705 2070 -8649
rect 2126 -8705 2150 -8649
rect 2206 -8705 8265 -8649
rect -21724 -8736 -7353 -8714
rect -46 -8727 8265 -8705
rect -21724 -8792 -21680 -8736
rect -21624 -8792 -21600 -8736
rect -21544 -8792 -21520 -8736
rect -21464 -8792 -20529 -8736
rect -20473 -8792 -20449 -8736
rect -20393 -8792 -20369 -8736
rect -20313 -8792 -15175 -8736
rect -15119 -8792 -15095 -8736
rect -15039 -8792 -15015 -8736
rect -14959 -8792 -7609 -8736
rect -7553 -8792 -7529 -8736
rect -7473 -8792 -7449 -8736
rect -7393 -8792 -7353 -8736
rect -21724 -8836 -7353 -8792
rect -21724 -8892 -21680 -8836
rect -21624 -8892 -21600 -8836
rect -21544 -8892 -21520 -8836
rect -21464 -8892 -20529 -8836
rect -20473 -8892 -20449 -8836
rect -20393 -8892 -20369 -8836
rect -20313 -8892 -15175 -8836
rect -15119 -8892 -15095 -8836
rect -15039 -8892 -15015 -8836
rect -14959 -8892 -7609 -8836
rect -7553 -8892 -7529 -8836
rect -7473 -8892 -7449 -8836
rect -7393 -8892 -7353 -8836
rect -21724 -8936 -7353 -8892
rect -21724 -8992 -21680 -8936
rect -21624 -8992 -21600 -8936
rect -21544 -8992 -21520 -8936
rect -21464 -8992 -20529 -8936
rect -20473 -8992 -20449 -8936
rect -20393 -8992 -20369 -8936
rect -20313 -8992 -15175 -8936
rect -15119 -8992 -15095 -8936
rect -15039 -8992 -15015 -8936
rect -14959 -8992 -7609 -8936
rect -7553 -8992 -7529 -8936
rect -7473 -8992 -7449 -8936
rect -7393 -8992 -7353 -8936
rect -21724 -9036 -7353 -8992
rect -21724 -9092 -21680 -9036
rect -21624 -9092 -21600 -9036
rect -21544 -9092 -21520 -9036
rect -21464 -9092 -20529 -9036
rect -20473 -9092 -20449 -9036
rect -20393 -9092 -20369 -9036
rect -20313 -9092 -15175 -9036
rect -15119 -9092 -15095 -9036
rect -15039 -9092 -15015 -9036
rect -14959 -9092 -7609 -9036
rect -7553 -9092 -7529 -9036
rect -7473 -9092 -7449 -9036
rect -7393 -9092 -7353 -9036
rect -21724 -9114 -7353 -9092
rect -3254 -8899 17620 -8877
rect -3254 -8955 -3214 -8899
rect -3158 -8955 -3134 -8899
rect -3078 -8955 -3054 -8899
rect -2998 -8955 -468 -8899
rect -412 -8955 -388 -8899
rect -332 -8955 -308 -8899
rect -252 -8955 4352 -8899
rect 4408 -8955 4432 -8899
rect 4488 -8955 4512 -8899
rect 4568 -8955 17360 -8899
rect 17416 -8955 17440 -8899
rect 17496 -8955 17520 -8899
rect 17576 -8955 17620 -8899
rect -3254 -8999 17620 -8955
rect -3254 -9055 -3214 -8999
rect -3158 -9055 -3134 -8999
rect -3078 -9055 -3054 -8999
rect -2998 -9055 -468 -8999
rect -412 -9055 -388 -8999
rect -332 -9055 -308 -8999
rect -252 -9055 4352 -8999
rect 4408 -9055 4432 -8999
rect 4488 -9055 4512 -8999
rect 4568 -9055 17360 -8999
rect 17416 -9055 17440 -8999
rect 17496 -9055 17520 -8999
rect 17576 -9055 17620 -8999
rect -3254 -9099 17620 -9055
rect -3254 -9155 -3214 -9099
rect -3158 -9155 -3134 -9099
rect -3078 -9155 -3054 -9099
rect -2998 -9155 -468 -9099
rect -412 -9155 -388 -9099
rect -332 -9155 -308 -9099
rect -252 -9155 4352 -9099
rect 4408 -9155 4432 -9099
rect 4488 -9155 4512 -9099
rect 4568 -9155 17360 -9099
rect 17416 -9155 17440 -9099
rect 17496 -9155 17520 -9099
rect 17576 -9155 17620 -9099
rect -3254 -9199 17620 -9155
rect -3254 -9255 -3214 -9199
rect -3158 -9255 -3134 -9199
rect -3078 -9255 -3054 -9199
rect -2998 -9255 -468 -9199
rect -412 -9255 -388 -9199
rect -332 -9255 -308 -9199
rect -252 -9255 4352 -9199
rect 4408 -9255 4432 -9199
rect 4488 -9255 4512 -9199
rect 4568 -9255 17360 -9199
rect 17416 -9255 17440 -9199
rect 17496 -9255 17520 -9199
rect 17576 -9255 17620 -9199
rect -3254 -9277 17620 -9255
rect 8690 -9528 16556 -9506
rect 8690 -9584 8730 -9528
rect 8786 -9584 8810 -9528
rect 8866 -9584 8890 -9528
rect 8946 -9584 13633 -9528
rect 13689 -9584 13713 -9528
rect 13769 -9584 13793 -9528
rect 13849 -9584 16296 -9528
rect 16352 -9584 16376 -9528
rect 16432 -9584 16456 -9528
rect 16512 -9584 16556 -9528
rect 8690 -9628 16556 -9584
rect 8690 -9684 8730 -9628
rect 8786 -9684 8810 -9628
rect 8866 -9684 8890 -9628
rect 8946 -9684 13633 -9628
rect 13689 -9684 13713 -9628
rect 13769 -9684 13793 -9628
rect 13849 -9684 16296 -9628
rect 16352 -9684 16376 -9628
rect 16432 -9684 16456 -9628
rect 16512 -9684 16556 -9628
rect 8690 -9728 16556 -9684
rect 8690 -9784 8730 -9728
rect 8786 -9784 8810 -9728
rect 8866 -9784 8890 -9728
rect 8946 -9784 13633 -9728
rect 13689 -9784 13713 -9728
rect 13769 -9784 13793 -9728
rect 13849 -9784 16296 -9728
rect 16352 -9784 16376 -9728
rect 16432 -9784 16456 -9728
rect 16512 -9784 16556 -9728
rect 8690 -9828 16556 -9784
rect 8690 -9884 8730 -9828
rect 8786 -9884 8810 -9828
rect 8866 -9884 8890 -9828
rect 8946 -9884 13633 -9828
rect 13689 -9884 13713 -9828
rect 13769 -9884 13793 -9828
rect 13849 -9884 16296 -9828
rect 16352 -9884 16376 -9828
rect 16432 -9884 16456 -9828
rect 16512 -9884 16556 -9828
rect -10861 -9908 -1978 -9886
rect 8690 -9906 16556 -9884
rect -10861 -9964 -10821 -9908
rect -10765 -9964 -10741 -9908
rect -10685 -9964 -10661 -9908
rect -10605 -9964 -2238 -9908
rect -2182 -9964 -2158 -9908
rect -2102 -9964 -2078 -9908
rect -2022 -9964 -1978 -9908
rect -10861 -10008 -1978 -9964
rect -10861 -10064 -10821 -10008
rect -10765 -10064 -10741 -10008
rect -10685 -10064 -10661 -10008
rect -10605 -10064 -2238 -10008
rect -2182 -10064 -2158 -10008
rect -2102 -10064 -2078 -10008
rect -2022 -10064 -1978 -10008
rect -10861 -10108 -1978 -10064
rect -10861 -10164 -10821 -10108
rect -10765 -10164 -10741 -10108
rect -10685 -10164 -10661 -10108
rect -10605 -10164 -2238 -10108
rect -2182 -10164 -2158 -10108
rect -2102 -10164 -2078 -10108
rect -2022 -10164 -1978 -10108
rect -10861 -10208 -1978 -10164
rect -10861 -10264 -10821 -10208
rect -10765 -10264 -10741 -10208
rect -10685 -10264 -10661 -10208
rect -10605 -10264 -2238 -10208
rect -2182 -10264 -2158 -10208
rect -2102 -10264 -2078 -10208
rect -2022 -10264 -1978 -10208
rect -10861 -10286 -1978 -10264
rect 6889 -10039 7441 -10017
rect 6889 -10095 6929 -10039
rect 6985 -10095 7009 -10039
rect 7065 -10095 7089 -10039
rect 7145 -10095 7441 -10039
rect 6889 -10117 7441 -10095
rect 18143 -10039 18695 -10017
rect 18143 -10095 18439 -10039
rect 18495 -10095 18519 -10039
rect 18575 -10095 18599 -10039
rect 18655 -10095 18695 -10039
rect 18143 -10117 18695 -10095
rect 6889 -10139 7749 -10117
rect 6889 -10195 6929 -10139
rect 6985 -10195 7009 -10139
rect 7065 -10195 7089 -10139
rect 7145 -10195 7749 -10139
rect 6889 -10217 7749 -10195
rect 17836 -10139 18695 -10117
rect 17836 -10195 18439 -10139
rect 18495 -10195 18519 -10139
rect 18575 -10195 18599 -10139
rect 18655 -10195 18695 -10139
rect 17836 -10217 18695 -10195
rect 6889 -10239 9486 -10217
rect 6889 -10295 6929 -10239
rect 6985 -10295 7009 -10239
rect 7065 -10295 7089 -10239
rect 7145 -10295 9486 -10239
rect 6889 -10317 9486 -10295
rect 16098 -10239 18695 -10217
rect 16098 -10295 18439 -10239
rect 18495 -10295 18519 -10239
rect 18575 -10295 18599 -10239
rect 18655 -10295 18695 -10239
rect 16098 -10317 18695 -10295
rect 6889 -10339 7749 -10317
rect 6889 -10395 6929 -10339
rect 6985 -10395 7009 -10339
rect 7065 -10395 7089 -10339
rect 7145 -10395 7749 -10339
rect 6889 -10417 7749 -10395
rect 17836 -10339 18695 -10317
rect 17836 -10395 18439 -10339
rect 18495 -10395 18519 -10339
rect 18575 -10395 18599 -10339
rect 18655 -10395 18695 -10339
rect 17836 -10417 18695 -10395
rect 6889 -10439 7441 -10417
rect 6889 -10495 6933 -10439
rect 6989 -10495 7013 -10439
rect 7069 -10495 7093 -10439
rect 7149 -10495 7441 -10439
rect 6889 -10517 7441 -10495
rect 18143 -10439 18695 -10417
rect 18143 -10495 18435 -10439
rect 18491 -10495 18515 -10439
rect 18571 -10495 18595 -10439
rect 18651 -10495 18695 -10439
rect 18143 -10517 18695 -10495
rect -7653 -10626 -2898 -10604
rect -7653 -10682 -7609 -10626
rect -7553 -10682 -7529 -10626
rect -7473 -10682 -7449 -10626
rect -7393 -10682 -3158 -10626
rect -3102 -10682 -3078 -10626
rect -3022 -10682 -2998 -10626
rect -2942 -10682 -2898 -10626
rect -7653 -10726 -2898 -10682
rect -7653 -10782 -7609 -10726
rect -7553 -10782 -7529 -10726
rect -7473 -10782 -7449 -10726
rect -7393 -10782 -3158 -10726
rect -3102 -10782 -3078 -10726
rect -3022 -10782 -2998 -10726
rect -2942 -10782 -2898 -10726
rect -1730 -10675 -1430 -10671
rect 3160 -10675 3460 -10671
rect -1730 -10693 508 -10675
rect -1730 -10749 -1690 -10693
rect -1634 -10749 -1610 -10693
rect -1554 -10749 -1530 -10693
rect -1474 -10749 508 -10693
rect -1730 -10771 508 -10749
rect 1222 -10693 3460 -10675
rect 1222 -10749 3204 -10693
rect 3260 -10749 3284 -10693
rect 3340 -10749 3364 -10693
rect 3420 -10749 3460 -10693
rect 1222 -10771 3460 -10749
rect 7965 -10675 8265 -10671
rect 17320 -10675 17620 -10671
rect 7965 -10693 10202 -10675
rect 7965 -10749 8005 -10693
rect 8061 -10749 8085 -10693
rect 8141 -10749 8165 -10693
rect 8221 -10749 10202 -10693
rect 7965 -10771 10202 -10749
rect 15383 -10693 17620 -10675
rect 15383 -10749 17364 -10693
rect 17420 -10749 17444 -10693
rect 17500 -10749 17524 -10693
rect 17580 -10749 17620 -10693
rect 15383 -10771 17620 -10749
rect -7653 -10826 -2898 -10782
rect -7653 -10882 -7609 -10826
rect -7553 -10882 -7529 -10826
rect -7473 -10882 -7449 -10826
rect -7393 -10882 -3158 -10826
rect -3102 -10882 -3078 -10826
rect -3022 -10882 -2998 -10826
rect -2942 -10882 -2898 -10826
rect -7653 -10926 -2898 -10882
rect -7653 -10982 -7609 -10926
rect -7553 -10982 -7529 -10926
rect -7473 -10982 -7449 -10926
rect -7393 -10982 -3158 -10926
rect -3102 -10982 -3078 -10926
rect -3022 -10982 -2998 -10926
rect -2942 -10982 -2898 -10926
rect -7653 -11004 -2898 -10982
rect -1730 -11010 508 -10988
rect -1730 -11066 -1690 -11010
rect -1634 -11066 -1610 -11010
rect -1554 -11066 -1530 -11010
rect -1474 -11066 508 -11010
rect -1730 -11084 508 -11066
rect 1222 -11010 3460 -10988
rect 1222 -11066 3204 -11010
rect 3260 -11066 3284 -11010
rect 3340 -11066 3364 -11010
rect 3420 -11066 3460 -11010
rect 1222 -11084 3460 -11066
rect -1730 -11088 -1430 -11084
rect 3160 -11088 3460 -11084
rect 7477 -11010 9715 -10988
rect 7477 -11066 7517 -11010
rect 7573 -11066 7597 -11010
rect 7653 -11066 7677 -11010
rect 7733 -11066 9715 -11010
rect 7477 -11084 9715 -11066
rect 11678 -11011 13916 -10988
rect 11678 -11067 12672 -11011
rect 12728 -11067 12752 -11011
rect 12808 -11067 12832 -11011
rect 12888 -11067 13916 -11011
rect 11678 -11084 13916 -11067
rect 15870 -11010 18107 -10988
rect 15870 -11066 17851 -11010
rect 17907 -11066 17931 -11010
rect 17987 -11066 18011 -11010
rect 18067 -11066 18107 -11010
rect 15870 -11084 18107 -11066
rect 7477 -11088 7777 -11084
rect 12632 -11089 12932 -11084
rect 17807 -11088 18107 -11084
rect -1730 -12073 -1430 -12068
rect 3160 -12073 3460 -12068
rect -1730 -12090 508 -12073
rect -1730 -12146 -1690 -12090
rect -1634 -12146 -1610 -12090
rect -1554 -12146 -1530 -12090
rect -1474 -12146 508 -12090
rect -1730 -12168 508 -12146
rect 1222 -12090 3460 -12073
rect 1222 -12146 3204 -12090
rect 3260 -12146 3284 -12090
rect 3340 -12146 3364 -12090
rect 3420 -12146 3460 -12090
rect 1222 -12168 3460 -12146
rect 7477 -12073 7777 -12068
rect 12632 -12073 12932 -12068
rect 17807 -12073 18107 -12068
rect 7477 -12090 9715 -12073
rect 7477 -12146 7517 -12090
rect 7573 -12146 7597 -12090
rect 7653 -12146 7677 -12090
rect 7733 -12146 9715 -12090
rect 7477 -12168 9715 -12146
rect 11678 -12090 13916 -12073
rect 11678 -12146 12672 -12090
rect 12728 -12146 12752 -12090
rect 12808 -12146 12832 -12090
rect 12888 -12146 13916 -12090
rect 11678 -12168 13916 -12146
rect 15870 -12090 18107 -12073
rect 15870 -12146 17851 -12090
rect 17907 -12146 17931 -12090
rect 17987 -12146 18011 -12090
rect 18067 -12146 18107 -12090
rect 15870 -12168 18107 -12146
rect -1730 -12408 508 -12386
rect -1730 -12464 -1690 -12408
rect -1634 -12464 -1610 -12408
rect -1554 -12464 -1530 -12408
rect -1474 -12464 508 -12408
rect -1730 -12481 508 -12464
rect 1222 -12408 3460 -12386
rect 1222 -12464 3204 -12408
rect 3260 -12464 3284 -12408
rect 3340 -12464 3364 -12408
rect 3420 -12464 3460 -12408
rect 1222 -12481 3460 -12464
rect -1730 -12486 -1430 -12481
rect 3160 -12486 3460 -12481
rect 7965 -12408 10202 -12386
rect 7965 -12464 8005 -12408
rect 8061 -12464 8085 -12408
rect 8141 -12464 8165 -12408
rect 8221 -12464 10202 -12408
rect 7965 -12481 10202 -12464
rect 15383 -12408 17620 -12386
rect 15383 -12464 17364 -12408
rect 17420 -12464 17444 -12408
rect 17500 -12464 17524 -12408
rect 17580 -12464 17620 -12408
rect 15383 -12481 17620 -12464
rect 7965 -12486 8265 -12481
rect 17320 -12486 17620 -12481
rect 8754 -13150 12377 -12981
rect 13161 -13150 16785 -12981
rect -3198 -13365 2682 -13343
rect -3198 -13421 -3158 -13365
rect -3102 -13421 -3078 -13365
rect -3022 -13421 -2998 -13365
rect -2942 -13421 220 -13365
rect 276 -13421 300 -13365
rect 356 -13421 380 -13365
rect 436 -13421 1301 -13365
rect 1357 -13421 1381 -13365
rect 1437 -13421 1461 -13365
rect 1517 -13421 2422 -13365
rect 2478 -13421 2502 -13365
rect 2558 -13421 2582 -13365
rect 2638 -13421 2682 -13365
rect -3198 -13465 2682 -13421
rect -3198 -13521 -3158 -13465
rect -3102 -13521 -3078 -13465
rect -3022 -13521 -2998 -13465
rect -2942 -13521 220 -13465
rect 276 -13521 300 -13465
rect 356 -13521 380 -13465
rect 436 -13521 1301 -13465
rect 1357 -13521 1381 -13465
rect 1437 -13521 1461 -13465
rect 1517 -13521 2422 -13465
rect 2478 -13521 2502 -13465
rect 2558 -13521 2582 -13465
rect 2638 -13521 2682 -13465
rect -3198 -13565 2682 -13521
rect -3198 -13621 -3158 -13565
rect -3102 -13621 -3078 -13565
rect -3022 -13621 -2998 -13565
rect -2942 -13621 220 -13565
rect 276 -13621 300 -13565
rect 356 -13621 380 -13565
rect 436 -13621 1301 -13565
rect 1357 -13621 1381 -13565
rect 1437 -13621 1461 -13565
rect 1517 -13621 2422 -13565
rect 2478 -13621 2502 -13565
rect 2558 -13621 2582 -13565
rect 2638 -13621 2682 -13565
rect -3198 -13665 2682 -13621
rect -3198 -13721 -3158 -13665
rect -3102 -13721 -3078 -13665
rect -3022 -13721 -2998 -13665
rect -2942 -13721 220 -13665
rect 276 -13721 300 -13665
rect 356 -13721 380 -13665
rect 436 -13721 1301 -13665
rect 1357 -13721 1381 -13665
rect 1437 -13721 1461 -13665
rect 1517 -13721 2422 -13665
rect 2478 -13721 2502 -13665
rect 2558 -13721 2582 -13665
rect 2638 -13721 2682 -13665
rect -3198 -13743 2682 -13721
rect 9622 -13484 15920 -13462
rect 9622 -13540 9662 -13484
rect 9718 -13540 9742 -13484
rect 9798 -13540 9822 -13484
rect 9878 -13540 13201 -13484
rect 13257 -13540 13281 -13484
rect 13337 -13540 13361 -13484
rect 13417 -13540 15660 -13484
rect 15716 -13540 15740 -13484
rect 15796 -13540 15820 -13484
rect 15876 -13540 15920 -13484
rect 9622 -13584 15920 -13540
rect 9622 -13640 9662 -13584
rect 9718 -13640 9742 -13584
rect 9798 -13640 9822 -13584
rect 9878 -13640 13201 -13584
rect 13257 -13640 13281 -13584
rect 13337 -13640 13361 -13584
rect 13417 -13640 15660 -13584
rect 15716 -13640 15740 -13584
rect 15796 -13640 15820 -13584
rect 15876 -13640 15920 -13584
rect 9622 -13684 15920 -13640
rect 9622 -13740 9662 -13684
rect 9718 -13740 9742 -13684
rect 9798 -13740 9822 -13684
rect 9878 -13740 13201 -13684
rect 13257 -13740 13281 -13684
rect 13337 -13740 13361 -13684
rect 13417 -13740 15660 -13684
rect 15716 -13740 15740 -13684
rect 15796 -13740 15820 -13684
rect 15876 -13740 15920 -13684
rect 9622 -13784 15920 -13740
rect 9622 -13840 9662 -13784
rect 9718 -13840 9742 -13784
rect 9798 -13840 9822 -13784
rect 9878 -13840 13201 -13784
rect 13257 -13840 13281 -13784
rect 13337 -13840 13361 -13784
rect 13417 -13840 15660 -13784
rect 15716 -13840 15740 -13784
rect 15796 -13840 15820 -13784
rect 15876 -13840 15920 -13784
rect 9622 -13862 15920 -13840
rect -2308 -14025 4019 -14003
rect -2308 -14081 -2238 -14025
rect -2182 -14081 -2158 -14025
rect -2102 -14081 -2078 -14025
rect -2022 -14081 -901 -14025
rect -845 -14081 -821 -14025
rect -765 -14081 -741 -14025
rect -685 -14081 3759 -14025
rect 3815 -14081 3839 -14025
rect 3895 -14081 3919 -14025
rect 3975 -14081 4019 -14025
rect -2308 -14125 4019 -14081
rect -2308 -14181 -2238 -14125
rect -2182 -14181 -2158 -14125
rect -2102 -14181 -2078 -14125
rect -2022 -14181 -901 -14125
rect -845 -14181 -821 -14125
rect -765 -14181 -741 -14125
rect -685 -14181 3759 -14125
rect 3815 -14181 3839 -14125
rect 3895 -14181 3919 -14125
rect 3975 -14181 4019 -14125
rect -2308 -14225 4019 -14181
rect -2308 -14281 -2238 -14225
rect -2182 -14281 -2158 -14225
rect -2102 -14281 -2078 -14225
rect -2022 -14281 -901 -14225
rect -845 -14281 -821 -14225
rect -765 -14281 -741 -14225
rect -685 -14281 3759 -14225
rect 3815 -14281 3839 -14225
rect 3895 -14281 3919 -14225
rect 3975 -14281 4019 -14225
rect -2308 -14325 4019 -14281
rect -2308 -14381 -2238 -14325
rect -2182 -14381 -2158 -14325
rect -2102 -14381 -2078 -14325
rect -2022 -14381 -901 -14325
rect -845 -14381 -821 -14325
rect -765 -14381 -741 -14325
rect -685 -14381 3759 -14325
rect 3815 -14381 3839 -14325
rect 3895 -14381 3919 -14325
rect 3975 -14381 4019 -14325
rect -2308 -14403 4019 -14381
rect 12081 -14040 13461 -14018
rect 12081 -14096 12121 -14040
rect 12177 -14096 12201 -14040
rect 12257 -14096 12281 -14040
rect 12337 -14096 13201 -14040
rect 13257 -14096 13281 -14040
rect 13337 -14096 13361 -14040
rect 13417 -14096 13461 -14040
rect 12081 -14140 13461 -14096
rect 12081 -14196 12121 -14140
rect 12177 -14196 12201 -14140
rect 12257 -14196 12281 -14140
rect 12337 -14196 13201 -14140
rect 13257 -14196 13281 -14140
rect 13337 -14196 13361 -14140
rect 13417 -14196 13461 -14140
rect 12081 -14240 13461 -14196
rect 12081 -14296 12121 -14240
rect 12177 -14296 12201 -14240
rect 12257 -14296 12281 -14240
rect 12337 -14296 13201 -14240
rect 13257 -14296 13281 -14240
rect 13337 -14296 13361 -14240
rect 13417 -14296 13461 -14240
rect 12081 -14340 13461 -14296
rect 12081 -14396 12121 -14340
rect 12177 -14396 12201 -14340
rect 12257 -14396 12281 -14340
rect 12337 -14396 13201 -14340
rect 13257 -14396 13281 -14340
rect 13337 -14396 13361 -14340
rect 13417 -14396 13461 -14340
rect 12081 -14418 13461 -14396
rect -2631 -14619 -2435 -14611
rect -2631 -14671 -2622 -14619
rect -2570 -14671 -2558 -14619
rect -2506 -14671 -2494 -14619
rect -2442 -14671 -2435 -14619
rect -2631 -14681 -2435 -14671
rect 4199 -14619 4395 -14611
rect 4199 -14671 4208 -14619
rect 4260 -14671 4272 -14619
rect 4324 -14671 4336 -14619
rect 4388 -14671 4395 -14619
rect 4199 -14681 4395 -14671
rect 9232 -14619 9428 -14611
rect 9232 -14671 9241 -14619
rect 9293 -14671 9305 -14619
rect 9357 -14671 9369 -14619
rect 9421 -14671 9428 -14619
rect 9232 -14681 9428 -14671
rect 16098 -14619 16294 -14611
rect 16098 -14671 16107 -14619
rect 16159 -14671 16171 -14619
rect 16223 -14671 16235 -14619
rect 16287 -14671 16294 -14619
rect 16098 -14681 16294 -14671
rect 649 -14734 845 -14726
rect 649 -14786 658 -14734
rect 710 -14786 722 -14734
rect 774 -14786 786 -14734
rect 838 -14786 845 -14734
rect 649 -14796 845 -14786
rect 1030 -14734 1226 -14726
rect 1030 -14786 1039 -14734
rect 1091 -14786 1103 -14734
rect 1155 -14786 1167 -14734
rect 1219 -14786 1226 -14734
rect 1030 -14796 1226 -14786
rect 12495 -14734 12691 -14726
rect 12495 -14786 12504 -14734
rect 12556 -14786 12568 -14734
rect 12620 -14786 12632 -14734
rect 12684 -14786 12691 -14734
rect 12495 -14796 12691 -14786
rect 12909 -14734 13105 -14726
rect 12909 -14786 12918 -14734
rect 12970 -14786 12982 -14734
rect 13034 -14786 13046 -14734
rect 13098 -14786 13105 -14734
rect 12909 -14796 13105 -14786
rect -3497 -15310 -3197 -15306
rect 4894 -15310 5194 -15306
rect 8404 -15310 8704 -15306
rect 16794 -15310 17094 -15306
rect -3497 -15328 -1259 -15310
rect -3497 -15384 -3457 -15328
rect -3401 -15384 -3377 -15328
rect -3321 -15384 -3297 -15328
rect -3241 -15384 -1259 -15328
rect -3497 -15406 -1259 -15384
rect 2957 -15328 11293 -15310
rect 2957 -15384 4938 -15328
rect 4994 -15384 5018 -15328
rect 5074 -15384 5098 -15328
rect 5154 -15384 8444 -15328
rect 8500 -15384 8524 -15328
rect 8580 -15384 8604 -15328
rect 8660 -15384 11293 -15328
rect 2957 -15406 11293 -15384
rect 14857 -15328 17094 -15310
rect 14857 -15384 16838 -15328
rect 16894 -15384 16918 -15328
rect 16974 -15384 16998 -15328
rect 17054 -15384 17094 -15328
rect 14857 -15406 17094 -15384
rect -3497 -15645 -1259 -15623
rect -3497 -15701 -3457 -15645
rect -3401 -15701 -3377 -15645
rect -3321 -15701 -3297 -15645
rect -3241 -15701 -1259 -15645
rect -3497 -15719 -1259 -15701
rect 2957 -15645 11293 -15623
rect 2957 -15701 4938 -15645
rect 4994 -15701 5018 -15645
rect 5074 -15701 5098 -15645
rect 5154 -15701 8444 -15645
rect 8500 -15701 8524 -15645
rect 8580 -15701 8604 -15645
rect 8660 -15701 11293 -15645
rect 2957 -15719 11293 -15701
rect 14857 -15645 17094 -15623
rect 14857 -15701 16838 -15645
rect 16894 -15701 16918 -15645
rect 16974 -15701 16998 -15645
rect 17054 -15701 17094 -15645
rect 14857 -15719 17094 -15701
rect -3497 -15723 -3197 -15719
rect 4894 -15723 5194 -15719
rect 8404 -15723 8704 -15719
rect 16794 -15723 17094 -15719
rect -2640 -16244 -2444 -16234
rect -2640 -16296 -2633 -16244
rect -2581 -16296 -2569 -16244
rect -2517 -16296 -2505 -16244
rect -2453 -16296 -2444 -16244
rect -2640 -16304 -2444 -16296
rect 4190 -16244 4386 -16234
rect 4190 -16296 4197 -16244
rect 4249 -16296 4261 -16244
rect 4313 -16296 4325 -16244
rect 4377 -16296 4386 -16244
rect 4190 -16304 4386 -16296
rect 9223 -16244 9419 -16234
rect 9223 -16296 9230 -16244
rect 9282 -16296 9294 -16244
rect 9346 -16296 9358 -16244
rect 9410 -16296 9419 -16244
rect 9223 -16304 9419 -16296
rect 16089 -16244 16285 -16234
rect 16089 -16296 16096 -16244
rect 16148 -16296 16160 -16244
rect 16212 -16296 16224 -16244
rect 16276 -16296 16285 -16244
rect 16089 -16304 16285 -16296
rect 623 -16343 819 -16333
rect 623 -16395 630 -16343
rect 682 -16395 694 -16343
rect 746 -16395 758 -16343
rect 810 -16395 819 -16343
rect 623 -16403 819 -16395
rect 1004 -16343 1200 -16333
rect 1004 -16395 1011 -16343
rect 1063 -16395 1075 -16343
rect 1127 -16395 1139 -16343
rect 1191 -16395 1200 -16343
rect 1004 -16403 1200 -16395
rect 12469 -16343 12665 -16333
rect 12469 -16395 12476 -16343
rect 12528 -16395 12540 -16343
rect 12592 -16395 12604 -16343
rect 12656 -16395 12665 -16343
rect 12469 -16403 12665 -16395
rect 12883 -16343 13079 -16333
rect 12883 -16395 12890 -16343
rect 12942 -16395 12954 -16343
rect 13006 -16395 13018 -16343
rect 13070 -16395 13079 -16343
rect 12883 -16403 13079 -16395
rect -3497 -16707 -3197 -16703
rect 4894 -16707 5194 -16703
rect 8404 -16707 8704 -16703
rect 16794 -16707 17094 -16703
rect -3497 -16725 -1259 -16707
rect -3497 -16781 -3457 -16725
rect -3401 -16781 -3377 -16725
rect -3321 -16781 -3297 -16725
rect -3241 -16781 -1259 -16725
rect -3497 -16803 -1259 -16781
rect 2957 -16725 11293 -16707
rect 2957 -16781 4938 -16725
rect 4994 -16781 5018 -16725
rect 5074 -16781 5098 -16725
rect 5154 -16781 8444 -16725
rect 8500 -16781 8524 -16725
rect 8580 -16781 8604 -16725
rect 8660 -16781 11293 -16725
rect 2957 -16803 11293 -16781
rect 14857 -16725 17094 -16707
rect 14857 -16781 16838 -16725
rect 16894 -16781 16918 -16725
rect 16974 -16781 16998 -16725
rect 17054 -16781 17094 -16725
rect 14857 -16803 17094 -16781
rect -3497 -17042 -1259 -17020
rect -3497 -17098 -3457 -17042
rect -3401 -17098 -3377 -17042
rect -3321 -17098 -3297 -17042
rect -3241 -17098 -1259 -17042
rect -3497 -17116 -1259 -17098
rect 2957 -17042 11293 -17020
rect 2957 -17098 4938 -17042
rect 4994 -17098 5018 -17042
rect 5074 -17098 5098 -17042
rect 5154 -17098 8444 -17042
rect 8500 -17098 8524 -17042
rect 8580 -17098 8604 -17042
rect 8660 -17098 11293 -17042
rect 2957 -17116 11293 -17098
rect 14857 -17042 17094 -17020
rect 14857 -17098 16838 -17042
rect 16894 -17098 16918 -17042
rect 16974 -17098 16998 -17042
rect 17054 -17098 17094 -17042
rect 14857 -17116 17094 -17098
rect -3497 -17120 -3197 -17116
rect 4894 -17120 5194 -17116
rect 8404 -17120 8704 -17116
rect 16794 -17120 17094 -17116
rect 601 -17626 797 -17616
rect 601 -17678 608 -17626
rect 660 -17678 672 -17626
rect 724 -17678 736 -17626
rect 788 -17678 797 -17626
rect 601 -17686 797 -17678
rect 981 -17626 1177 -17616
rect 981 -17678 988 -17626
rect 1040 -17678 1052 -17626
rect 1104 -17678 1116 -17626
rect 1168 -17678 1177 -17626
rect 981 -17686 1177 -17678
rect 12446 -17626 12642 -17616
rect 12446 -17678 12453 -17626
rect 12505 -17678 12517 -17626
rect 12569 -17678 12581 -17626
rect 12633 -17678 12642 -17626
rect 12446 -17686 12642 -17678
rect 12860 -17626 13056 -17616
rect 12860 -17678 12867 -17626
rect 12919 -17678 12931 -17626
rect 12983 -17678 12995 -17626
rect 13047 -17678 13056 -17626
rect 12860 -17686 13056 -17678
rect -2633 -17725 -2437 -17715
rect -2633 -17777 -2626 -17725
rect -2574 -17777 -2562 -17725
rect -2510 -17777 -2498 -17725
rect -2446 -17777 -2437 -17725
rect -2633 -17785 -2437 -17777
rect 4197 -17725 4393 -17715
rect 4197 -17777 4204 -17725
rect 4256 -17777 4268 -17725
rect 4320 -17777 4332 -17725
rect 4384 -17777 4393 -17725
rect 4197 -17785 4393 -17777
rect 9230 -17725 9426 -17715
rect 9230 -17777 9237 -17725
rect 9289 -17777 9301 -17725
rect 9353 -17777 9365 -17725
rect 9417 -17777 9426 -17725
rect 9230 -17785 9426 -17777
rect 16096 -17725 16292 -17715
rect 16096 -17777 16103 -17725
rect 16155 -17777 16167 -17725
rect 16219 -17777 16231 -17725
rect 16283 -17777 16292 -17725
rect 16096 -17785 16292 -17777
<< via2 >>
rect -25719 10432 -25663 10488
rect -25639 10432 -25583 10488
rect -25559 10432 -25503 10488
rect -6573 10432 -6517 10488
rect -6493 10432 -6437 10488
rect -6413 10432 -6357 10488
rect -4706 10432 -4650 10488
rect -4626 10432 -4570 10488
rect -4546 10432 -4490 10488
rect 5793 10432 5849 10488
rect 5873 10432 5929 10488
rect 5953 10432 6009 10488
rect 6929 10432 6985 10488
rect 7009 10432 7065 10488
rect 7089 10432 7145 10488
rect 18435 10432 18491 10488
rect 18515 10432 18571 10488
rect 18595 10432 18651 10488
rect -25719 10112 -25663 10168
rect -25639 10112 -25583 10168
rect -25559 10112 -25503 10168
rect -6573 10112 -6517 10168
rect -6493 10112 -6437 10168
rect -6413 10112 -6357 10168
rect 5793 10111 5849 10167
rect 5873 10111 5929 10167
rect 5953 10111 6009 10167
rect 6929 10111 6985 10167
rect 7009 10111 7065 10167
rect 7089 10111 7145 10167
rect 18435 10111 18491 10167
rect 18515 10111 18571 10167
rect 18595 10111 18651 10167
rect 9856 9534 9912 9590
rect 9936 9534 9992 9590
rect 10016 9534 10072 9590
rect 15170 9534 15226 9590
rect 15250 9534 15306 9590
rect 15330 9534 15386 9590
rect 10828 9373 10884 9429
rect 10908 9373 10964 9429
rect 10988 9373 11044 9429
rect 14206 9373 14262 9429
rect 14286 9373 14342 9429
rect 14366 9373 14422 9429
rect -25719 8785 -25663 8841
rect -25639 8785 -25583 8841
rect -25559 8785 -25503 8841
rect -6573 8785 -6517 8841
rect -6493 8785 -6437 8841
rect -6413 8785 -6357 8841
rect 5793 8785 5849 8841
rect 5873 8785 5929 8841
rect 5953 8785 6009 8841
rect 6929 8785 6985 8841
rect 7009 8785 7065 8841
rect 7089 8785 7145 8841
rect 18435 8785 18491 8841
rect 18515 8785 18571 8841
rect 18595 8785 18651 8841
rect -25719 8453 -25663 8509
rect -25639 8453 -25583 8509
rect -25559 8453 -25503 8509
rect -6573 8453 -6517 8509
rect -6493 8453 -6437 8509
rect -6413 8453 -6357 8509
rect -4706 8453 -4650 8509
rect -4626 8453 -4570 8509
rect -4546 8453 -4490 8509
rect 5793 8453 5849 8509
rect 5873 8453 5929 8509
rect 5953 8453 6009 8509
rect 6929 8453 6985 8509
rect 7009 8453 7065 8509
rect 7089 8453 7145 8509
rect 18435 8453 18491 8509
rect 18515 8453 18571 8509
rect 18595 8453 18651 8509
rect 9856 8021 9912 8077
rect 9936 8021 9992 8077
rect 10016 8021 10072 8077
rect 15170 8021 15226 8077
rect 15250 8021 15306 8077
rect 15330 8021 15386 8077
rect 10828 7853 10884 7909
rect 10908 7853 10964 7909
rect 10988 7853 11044 7909
rect 14206 7853 14262 7909
rect 14286 7853 14342 7909
rect 14366 7853 14422 7909
rect 10828 6159 10884 6215
rect 10908 6159 10964 6215
rect 10988 6159 11044 6215
rect 14206 6159 14262 6215
rect 14286 6159 14342 6215
rect 14366 6159 14422 6215
rect 9856 5990 9912 6046
rect 9936 5990 9992 6046
rect 10016 5990 10072 6046
rect 15170 5990 15226 6046
rect 15250 5990 15306 6046
rect 15330 5990 15386 6046
rect -25719 5559 -25663 5615
rect -25639 5559 -25583 5615
rect -25559 5559 -25503 5615
rect -6573 5559 -6517 5615
rect -6493 5559 -6437 5615
rect -6413 5559 -6357 5615
rect -4706 5558 -4650 5614
rect -4626 5558 -4570 5614
rect -4546 5558 -4490 5614
rect 5793 5558 5849 5614
rect 5873 5558 5929 5614
rect 5953 5558 6009 5614
rect 6929 5558 6985 5614
rect 7009 5558 7065 5614
rect 7089 5558 7145 5614
rect 18435 5558 18491 5614
rect 18515 5558 18571 5614
rect 18595 5558 18651 5614
rect -25719 5227 -25663 5283
rect -25639 5227 -25583 5283
rect -25559 5227 -25503 5283
rect -6573 5227 -6517 5283
rect -6493 5227 -6437 5283
rect -6413 5227 -6357 5283
rect -4706 5238 -4650 5294
rect -4626 5238 -4570 5294
rect -4546 5238 -4490 5294
rect 5793 5232 5849 5288
rect 5873 5232 5929 5288
rect 5953 5232 6009 5288
rect 6929 5232 6985 5288
rect 7009 5232 7065 5288
rect 7089 5232 7145 5288
rect 18435 5232 18491 5288
rect 18515 5232 18571 5288
rect 18595 5232 18651 5288
rect 10828 4639 10884 4695
rect 10908 4639 10964 4695
rect 10988 4639 11044 4695
rect 14206 4639 14262 4695
rect 14286 4639 14342 4695
rect 14366 4639 14422 4695
rect 9856 4478 9912 4534
rect 9936 4478 9992 4534
rect 10016 4478 10072 4534
rect 15170 4478 15226 4534
rect 15250 4478 15306 4534
rect 15330 4478 15386 4534
rect -25719 3900 -25663 3956
rect -25639 3900 -25583 3956
rect -25559 3900 -25503 3956
rect -6573 3900 -6517 3956
rect -6493 3900 -6437 3956
rect -6413 3900 -6357 3956
rect -4706 3900 -4650 3956
rect -4626 3900 -4570 3956
rect -4546 3900 -4490 3956
rect 5793 3900 5849 3956
rect 5873 3900 5929 3956
rect 5953 3900 6009 3956
rect 6929 3900 6985 3956
rect 7009 3900 7065 3956
rect 7089 3900 7145 3956
rect 18435 3900 18491 3956
rect 18515 3900 18571 3956
rect 18595 3900 18651 3956
rect -25719 3580 -25663 3636
rect -25639 3580 -25583 3636
rect -25559 3580 -25503 3636
rect -6573 3580 -6517 3636
rect -6493 3580 -6437 3636
rect -6413 3580 -6357 3636
rect -4706 3580 -4650 3636
rect -4626 3580 -4570 3636
rect -4546 3580 -4490 3636
rect 5793 3580 5849 3636
rect 5873 3580 5929 3636
rect 5953 3580 6009 3636
rect 6929 3580 6985 3636
rect 7009 3580 7065 3636
rect 7089 3580 7145 3636
rect 18435 3580 18491 3636
rect 18515 3580 18571 3636
rect 18595 3580 18651 3636
rect -11240 2441 -11184 2497
rect -11160 2441 -11104 2497
rect -11080 2441 -11024 2497
rect -10531 2441 -10475 2497
rect -10451 2441 -10395 2497
rect -10371 2441 -10315 2497
rect -11240 2341 -11184 2397
rect -11160 2341 -11104 2397
rect -11080 2341 -11024 2397
rect -10531 2341 -10475 2397
rect -10451 2341 -10395 2397
rect -10371 2341 -10315 2397
rect -6 2358 50 2414
rect 74 2358 130 2414
rect 154 2358 210 2414
rect 562 2358 618 2414
rect 642 2358 698 2414
rect 722 2358 778 2414
rect 1144 2358 1200 2414
rect 1224 2358 1280 2414
rect 1304 2358 1360 2414
rect -6 2258 50 2314
rect 74 2258 130 2314
rect 154 2258 210 2314
rect 562 2258 618 2314
rect 642 2258 698 2314
rect 722 2258 778 2314
rect 1144 2258 1200 2314
rect 1224 2258 1280 2314
rect 1304 2258 1360 2314
rect -24315 2084 -24259 2140
rect -24235 2084 -24179 2140
rect -24155 2084 -24099 2140
rect -16749 2084 -16693 2140
rect -16669 2084 -16613 2140
rect -16589 2084 -16533 2140
rect -15598 2084 -15542 2140
rect -15518 2084 -15462 2140
rect -15438 2084 -15382 2140
rect -11400 2084 -11344 2140
rect -11320 2084 -11264 2140
rect -11240 2084 -11184 2140
rect -8032 2084 -7976 2140
rect -7952 2084 -7896 2140
rect -7872 2084 -7816 2140
rect -7187 2084 -7131 2140
rect -7107 2084 -7051 2140
rect -7027 2084 -6971 2140
rect -24315 1984 -24259 2040
rect -24235 1984 -24179 2040
rect -24155 1984 -24099 2040
rect -16749 1984 -16693 2040
rect -16669 1984 -16613 2040
rect -16589 1984 -16533 2040
rect -15598 1984 -15542 2040
rect -15518 1984 -15462 2040
rect -15438 1984 -15382 2040
rect -11400 1984 -11344 2040
rect -11320 1984 -11264 2040
rect -11240 1984 -11184 2040
rect -8032 1984 -7976 2040
rect -7952 1984 -7896 2040
rect -7872 1984 -7816 2040
rect -7187 1984 -7131 2040
rect -7107 1984 -7051 2040
rect -7027 1984 -6971 2040
rect -6 2158 50 2214
rect 74 2158 130 2214
rect 154 2158 210 2214
rect 562 2158 618 2214
rect 642 2158 698 2214
rect 722 2158 778 2214
rect 1144 2158 1200 2214
rect 1224 2158 1280 2214
rect 1304 2158 1360 2214
rect -6 2058 50 2114
rect 74 2058 130 2114
rect 154 2058 210 2114
rect 562 2058 618 2114
rect 642 2058 698 2114
rect 722 2058 778 2114
rect 1144 2058 1200 2114
rect 1224 2058 1280 2114
rect 1304 2058 1360 2114
rect -25310 1735 -25254 1791
rect -25230 1735 -25174 1791
rect -25150 1735 -25094 1791
rect -21107 1735 -21051 1791
rect -21027 1735 -20971 1791
rect -20947 1735 -20891 1791
rect -19957 1735 -19901 1791
rect -19877 1735 -19821 1791
rect -19797 1735 -19741 1791
rect -16899 1735 -16843 1791
rect -16819 1735 -16763 1791
rect -16739 1735 -16683 1791
rect -12390 1735 -12334 1791
rect -12310 1735 -12254 1791
rect -12230 1735 -12174 1791
rect -10531 1735 -10475 1791
rect -10451 1735 -10395 1791
rect -10371 1735 -10315 1791
rect -25310 1635 -25254 1691
rect -25230 1635 -25174 1691
rect -25150 1635 -25094 1691
rect -21107 1635 -21051 1691
rect -21027 1635 -20971 1691
rect -20947 1635 -20891 1691
rect -19957 1635 -19901 1691
rect -19877 1635 -19821 1691
rect -19797 1635 -19741 1691
rect -16899 1635 -16843 1691
rect -16819 1635 -16763 1691
rect -16739 1635 -16683 1691
rect -12390 1635 -12334 1691
rect -12310 1635 -12254 1691
rect -12230 1635 -12174 1691
rect -10531 1635 -10475 1691
rect -10451 1635 -10395 1691
rect -10371 1635 -10315 1691
rect -3636 1752 -3580 1808
rect -3556 1752 -3500 1808
rect -3476 1752 -3420 1808
rect -3214 1752 -3158 1808
rect -3134 1752 -3078 1808
rect -3054 1752 -2998 1808
rect 4352 1752 4408 1808
rect 4432 1752 4488 1808
rect 4512 1752 4568 1808
rect 4775 1752 4831 1808
rect 4855 1752 4911 1808
rect 4935 1752 4991 1808
rect -3636 1652 -3580 1708
rect -3556 1652 -3500 1708
rect -3476 1652 -3420 1708
rect -3214 1652 -3158 1708
rect -3134 1652 -3078 1708
rect -3054 1652 -2998 1708
rect 4352 1652 4408 1708
rect 4432 1652 4488 1708
rect 4512 1652 4568 1708
rect 4775 1652 4831 1708
rect 4855 1652 4911 1708
rect 4935 1652 4991 1708
rect -3636 1552 -3580 1608
rect -3556 1552 -3500 1608
rect -3476 1552 -3420 1608
rect -3214 1552 -3158 1608
rect -3134 1552 -3078 1608
rect -3054 1552 -2998 1608
rect 4352 1552 4408 1608
rect 4432 1552 4488 1608
rect 4512 1552 4568 1608
rect 4775 1552 4831 1608
rect 4855 1552 4911 1608
rect 4935 1552 4991 1608
rect -3636 1452 -3580 1508
rect -3556 1452 -3500 1508
rect -3476 1452 -3420 1508
rect -3214 1452 -3158 1508
rect -3134 1452 -3078 1508
rect -3054 1452 -2998 1508
rect 4352 1452 4408 1508
rect 4432 1452 4488 1508
rect 4512 1452 4568 1508
rect 4775 1452 4831 1508
rect 4855 1452 4911 1508
rect 4935 1452 4991 1508
rect 5793 1275 5849 1331
rect 5873 1275 5929 1331
rect 5953 1275 6009 1331
rect 6929 1275 6985 1331
rect 7009 1275 7065 1331
rect 7089 1275 7145 1331
rect 5793 1175 5849 1231
rect 5873 1175 5929 1231
rect 5953 1175 6009 1231
rect 6929 1175 6985 1231
rect 7009 1175 7065 1231
rect 7089 1175 7145 1231
rect 5793 1075 5849 1131
rect 5873 1075 5929 1131
rect 5953 1075 6009 1131
rect 6929 1075 6985 1131
rect 7009 1075 7065 1131
rect 7089 1075 7145 1131
rect 5793 975 5849 1031
rect 5873 975 5929 1031
rect 5953 975 6009 1031
rect 6929 975 6985 1031
rect 7009 975 7065 1031
rect 7089 975 7145 1031
rect -26492 238 -26436 294
rect -26412 238 -26356 294
rect -26332 238 -26276 294
rect -6061 238 -6005 294
rect -5981 238 -5925 294
rect -5901 238 -5845 294
rect -4706 238 -4650 294
rect -4626 238 -4570 294
rect -4546 238 -4490 294
rect 5793 238 5849 294
rect 5873 238 5929 294
rect 5953 238 6009 294
rect -26992 -83 -26936 -27
rect -26912 -83 -26856 -27
rect -26832 -83 -26776 -27
rect -5562 -83 -5506 -27
rect -5482 -83 -5426 -27
rect -5402 -83 -5346 -27
rect 9856 -660 9912 -604
rect 9936 -660 9992 -604
rect 10016 -660 10072 -604
rect 15170 -660 15226 -604
rect 15250 -660 15306 -604
rect 15330 -660 15386 -604
rect 10828 -821 10884 -765
rect 10908 -821 10964 -765
rect 10988 -821 11044 -765
rect 14206 -821 14262 -765
rect 14286 -821 14342 -765
rect 14366 -821 14422 -765
rect -26992 -1421 -26936 -1365
rect -26912 -1421 -26856 -1365
rect -26832 -1421 -26776 -1365
rect -5562 -1421 -5506 -1365
rect -5482 -1421 -5426 -1365
rect -5402 -1421 -5346 -1365
rect -26492 -1741 -26436 -1685
rect -26412 -1741 -26356 -1685
rect -26332 -1741 -26276 -1685
rect -6061 -1741 -6005 -1685
rect -5981 -1741 -5925 -1685
rect -5901 -1741 -5845 -1685
rect -4706 -1741 -4650 -1685
rect -4626 -1741 -4570 -1685
rect -4546 -1741 -4490 -1685
rect 5793 -1741 5849 -1685
rect 5873 -1741 5929 -1685
rect 5953 -1741 6009 -1685
rect 9856 -2173 9912 -2117
rect 9936 -2173 9992 -2117
rect 10016 -2173 10072 -2117
rect 15170 -2173 15226 -2117
rect 15250 -2173 15306 -2117
rect 15330 -2173 15386 -2117
rect 10828 -2341 10884 -2285
rect 10908 -2341 10964 -2285
rect 10988 -2341 11044 -2285
rect 14206 -2341 14262 -2285
rect 14286 -2341 14342 -2285
rect 14366 -2341 14422 -2285
rect 10828 -4035 10884 -3979
rect 10908 -4035 10964 -3979
rect 10988 -4035 11044 -3979
rect 14206 -4035 14262 -3979
rect 14286 -4035 14342 -3979
rect 14366 -4035 14422 -3979
rect 9856 -4204 9912 -4148
rect 9936 -4204 9992 -4148
rect 10016 -4204 10072 -4148
rect 15170 -4204 15226 -4148
rect 15250 -4204 15306 -4148
rect 15330 -4204 15386 -4148
rect -26492 -4636 -26436 -4580
rect -26412 -4636 -26356 -4580
rect -26332 -4636 -26276 -4580
rect -6061 -4636 -6005 -4580
rect -5981 -4636 -5925 -4580
rect -5901 -4636 -5845 -4580
rect -4706 -4636 -4650 -4580
rect -4626 -4636 -4570 -4580
rect -4546 -4636 -4490 -4580
rect 5793 -4636 5849 -4580
rect 5873 -4636 5929 -4580
rect 5953 -4636 6009 -4580
rect -26992 -4956 -26936 -4900
rect -26912 -4956 -26856 -4900
rect -26832 -4956 -26776 -4900
rect -5562 -4956 -5506 -4900
rect -5482 -4956 -5426 -4900
rect -5402 -4956 -5346 -4900
rect -4706 -4956 -4650 -4900
rect -4626 -4956 -4570 -4900
rect -4546 -4956 -4490 -4900
rect 5793 -4956 5849 -4900
rect 5873 -4956 5929 -4900
rect 5953 -4956 6009 -4900
rect 10828 -5555 10884 -5499
rect 10908 -5555 10964 -5499
rect 10988 -5555 11044 -5499
rect 14206 -5555 14262 -5499
rect 14286 -5555 14342 -5499
rect 14366 -5555 14422 -5499
rect 9856 -5716 9912 -5660
rect 9936 -5716 9992 -5660
rect 10016 -5716 10072 -5660
rect 15170 -5716 15226 -5660
rect 15250 -5716 15306 -5660
rect 15330 -5716 15386 -5660
rect -26992 -6294 -26936 -6238
rect -26912 -6294 -26856 -6238
rect -26832 -6294 -26776 -6238
rect -5562 -6294 -5506 -6238
rect -5482 -6294 -5426 -6238
rect -5402 -6294 -5346 -6238
rect -4706 -6294 -4650 -6238
rect -4626 -6294 -4570 -6238
rect -4546 -6294 -4490 -6238
rect 5793 -6294 5849 -6238
rect 5873 -6294 5929 -6238
rect 5953 -6294 6009 -6238
rect -26492 -6614 -26436 -6558
rect -26412 -6614 -26356 -6558
rect -26332 -6614 -26276 -6558
rect -6061 -6614 -6005 -6558
rect -5981 -6614 -5925 -6558
rect -5901 -6614 -5845 -6558
rect -4706 -6614 -4650 -6558
rect -4626 -6614 -4570 -6558
rect -4546 -6614 -4490 -6558
rect 5793 -6614 5849 -6558
rect 5873 -6614 5929 -6558
rect 5953 -6614 6009 -6558
rect 11796 -7836 11852 -7780
rect 11876 -7836 11932 -7780
rect 11956 -7836 12012 -7780
rect 13088 -7836 13144 -7780
rect 13168 -7836 13224 -7780
rect 13248 -7836 13304 -7780
rect 11796 -7936 11852 -7880
rect 11876 -7936 11932 -7880
rect 11956 -7936 12012 -7880
rect 13088 -7936 13144 -7880
rect 13168 -7936 13224 -7880
rect 13248 -7936 13304 -7880
rect -24892 -8074 -24836 -8018
rect -24812 -8074 -24756 -8018
rect -24732 -8074 -24676 -8018
rect -17326 -8074 -17270 -8018
rect -17246 -8074 -17190 -8018
rect -17166 -8074 -17110 -8018
rect -11972 -8074 -11916 -8018
rect -11892 -8074 -11836 -8018
rect -11812 -8074 -11756 -8018
rect -10821 -8074 -10765 -8018
rect -10741 -8074 -10685 -8018
rect -10661 -8074 -10605 -8018
rect -24892 -8174 -24836 -8118
rect -24812 -8174 -24756 -8118
rect -24732 -8174 -24676 -8118
rect -17326 -8174 -17270 -8118
rect -17246 -8174 -17190 -8118
rect -17166 -8174 -17110 -8118
rect -11972 -8174 -11916 -8118
rect -11892 -8174 -11836 -8118
rect -11812 -8174 -11756 -8118
rect -10821 -8174 -10765 -8118
rect -10741 -8174 -10685 -8118
rect -10661 -8174 -10605 -8118
rect 11796 -8036 11852 -7980
rect 11876 -8036 11932 -7980
rect 11956 -8036 12012 -7980
rect 13088 -8036 13144 -7980
rect 13168 -8036 13224 -7980
rect 13248 -8036 13304 -7980
rect 11796 -8136 11852 -8080
rect 11876 -8136 11932 -8080
rect 11956 -8136 12012 -8080
rect 13088 -8136 13144 -8080
rect 13168 -8136 13224 -8080
rect 13248 -8136 13304 -8080
rect -24892 -8274 -24836 -8218
rect -24812 -8274 -24756 -8218
rect -24732 -8274 -24676 -8218
rect -17326 -8274 -17270 -8218
rect -17246 -8274 -17190 -8218
rect -17166 -8274 -17110 -8218
rect -11972 -8274 -11916 -8218
rect -11892 -8274 -11836 -8218
rect -11812 -8274 -11756 -8218
rect -10821 -8274 -10765 -8218
rect -10741 -8274 -10685 -8218
rect -10661 -8274 -10605 -8218
rect -24892 -8374 -24836 -8318
rect -24812 -8374 -24756 -8318
rect -24732 -8374 -24676 -8318
rect -17326 -8374 -17270 -8318
rect -17246 -8374 -17190 -8318
rect -17166 -8374 -17110 -8318
rect -11972 -8374 -11916 -8318
rect -11892 -8374 -11836 -8318
rect -11812 -8374 -11756 -8318
rect -10821 -8374 -10765 -8318
rect -10741 -8374 -10685 -8318
rect -10661 -8374 -10605 -8318
rect -6 -8405 50 -8349
rect 74 -8405 130 -8349
rect 154 -8405 210 -8349
rect 1144 -8405 1200 -8349
rect 1224 -8405 1280 -8349
rect 1304 -8405 1360 -8349
rect 1990 -8405 2046 -8349
rect 2070 -8405 2126 -8349
rect 2150 -8405 2206 -8349
rect -6 -8505 50 -8449
rect 74 -8505 130 -8449
rect 154 -8505 210 -8449
rect 1144 -8505 1200 -8449
rect 1224 -8505 1280 -8449
rect 1304 -8505 1360 -8449
rect 1990 -8505 2046 -8449
rect 2070 -8505 2126 -8449
rect 2150 -8505 2206 -8449
rect -6 -8605 50 -8549
rect 74 -8605 130 -8549
rect 154 -8605 210 -8549
rect 1144 -8605 1200 -8549
rect 1224 -8605 1280 -8549
rect 1304 -8605 1360 -8549
rect 1990 -8605 2046 -8549
rect 2070 -8605 2126 -8549
rect 2150 -8605 2206 -8549
rect -6 -8705 50 -8649
rect 74 -8705 130 -8649
rect 154 -8705 210 -8649
rect 1144 -8705 1200 -8649
rect 1224 -8705 1280 -8649
rect 1304 -8705 1360 -8649
rect 1990 -8705 2046 -8649
rect 2070 -8705 2126 -8649
rect 2150 -8705 2206 -8649
rect -21680 -8792 -21624 -8736
rect -21600 -8792 -21544 -8736
rect -21520 -8792 -21464 -8736
rect -20529 -8792 -20473 -8736
rect -20449 -8792 -20393 -8736
rect -20369 -8792 -20313 -8736
rect -15175 -8792 -15119 -8736
rect -15095 -8792 -15039 -8736
rect -15015 -8792 -14959 -8736
rect -7609 -8792 -7553 -8736
rect -7529 -8792 -7473 -8736
rect -7449 -8792 -7393 -8736
rect -21680 -8892 -21624 -8836
rect -21600 -8892 -21544 -8836
rect -21520 -8892 -21464 -8836
rect -20529 -8892 -20473 -8836
rect -20449 -8892 -20393 -8836
rect -20369 -8892 -20313 -8836
rect -15175 -8892 -15119 -8836
rect -15095 -8892 -15039 -8836
rect -15015 -8892 -14959 -8836
rect -7609 -8892 -7553 -8836
rect -7529 -8892 -7473 -8836
rect -7449 -8892 -7393 -8836
rect -21680 -8992 -21624 -8936
rect -21600 -8992 -21544 -8936
rect -21520 -8992 -21464 -8936
rect -20529 -8992 -20473 -8936
rect -20449 -8992 -20393 -8936
rect -20369 -8992 -20313 -8936
rect -15175 -8992 -15119 -8936
rect -15095 -8992 -15039 -8936
rect -15015 -8992 -14959 -8936
rect -7609 -8992 -7553 -8936
rect -7529 -8992 -7473 -8936
rect -7449 -8992 -7393 -8936
rect -21680 -9092 -21624 -9036
rect -21600 -9092 -21544 -9036
rect -21520 -9092 -21464 -9036
rect -20529 -9092 -20473 -9036
rect -20449 -9092 -20393 -9036
rect -20369 -9092 -20313 -9036
rect -15175 -9092 -15119 -9036
rect -15095 -9092 -15039 -9036
rect -15015 -9092 -14959 -9036
rect -7609 -9092 -7553 -9036
rect -7529 -9092 -7473 -9036
rect -7449 -9092 -7393 -9036
rect -3214 -8955 -3158 -8899
rect -3134 -8955 -3078 -8899
rect -3054 -8955 -2998 -8899
rect -468 -8955 -412 -8899
rect -388 -8955 -332 -8899
rect -308 -8955 -252 -8899
rect 4352 -8955 4408 -8899
rect 4432 -8955 4488 -8899
rect 4512 -8955 4568 -8899
rect 17360 -8955 17416 -8899
rect 17440 -8955 17496 -8899
rect 17520 -8955 17576 -8899
rect -3214 -9055 -3158 -8999
rect -3134 -9055 -3078 -8999
rect -3054 -9055 -2998 -8999
rect -468 -9055 -412 -8999
rect -388 -9055 -332 -8999
rect -308 -9055 -252 -8999
rect 4352 -9055 4408 -8999
rect 4432 -9055 4488 -8999
rect 4512 -9055 4568 -8999
rect 17360 -9055 17416 -8999
rect 17440 -9055 17496 -8999
rect 17520 -9055 17576 -8999
rect -3214 -9155 -3158 -9099
rect -3134 -9155 -3078 -9099
rect -3054 -9155 -2998 -9099
rect -468 -9155 -412 -9099
rect -388 -9155 -332 -9099
rect -308 -9155 -252 -9099
rect 4352 -9155 4408 -9099
rect 4432 -9155 4488 -9099
rect 4512 -9155 4568 -9099
rect 17360 -9155 17416 -9099
rect 17440 -9155 17496 -9099
rect 17520 -9155 17576 -9099
rect -3214 -9255 -3158 -9199
rect -3134 -9255 -3078 -9199
rect -3054 -9255 -2998 -9199
rect -468 -9255 -412 -9199
rect -388 -9255 -332 -9199
rect -308 -9255 -252 -9199
rect 4352 -9255 4408 -9199
rect 4432 -9255 4488 -9199
rect 4512 -9255 4568 -9199
rect 17360 -9255 17416 -9199
rect 17440 -9255 17496 -9199
rect 17520 -9255 17576 -9199
rect 8730 -9584 8786 -9528
rect 8810 -9584 8866 -9528
rect 8890 -9584 8946 -9528
rect 13633 -9584 13689 -9528
rect 13713 -9584 13769 -9528
rect 13793 -9584 13849 -9528
rect 16296 -9584 16352 -9528
rect 16376 -9584 16432 -9528
rect 16456 -9584 16512 -9528
rect 8730 -9684 8786 -9628
rect 8810 -9684 8866 -9628
rect 8890 -9684 8946 -9628
rect 13633 -9684 13689 -9628
rect 13713 -9684 13769 -9628
rect 13793 -9684 13849 -9628
rect 16296 -9684 16352 -9628
rect 16376 -9684 16432 -9628
rect 16456 -9684 16512 -9628
rect 8730 -9784 8786 -9728
rect 8810 -9784 8866 -9728
rect 8890 -9784 8946 -9728
rect 13633 -9784 13689 -9728
rect 13713 -9784 13769 -9728
rect 13793 -9784 13849 -9728
rect 16296 -9784 16352 -9728
rect 16376 -9784 16432 -9728
rect 16456 -9784 16512 -9728
rect 8730 -9884 8786 -9828
rect 8810 -9884 8866 -9828
rect 8890 -9884 8946 -9828
rect 13633 -9884 13689 -9828
rect 13713 -9884 13769 -9828
rect 13793 -9884 13849 -9828
rect 16296 -9884 16352 -9828
rect 16376 -9884 16432 -9828
rect 16456 -9884 16512 -9828
rect -10821 -9964 -10765 -9908
rect -10741 -9964 -10685 -9908
rect -10661 -9964 -10605 -9908
rect -2238 -9964 -2182 -9908
rect -2158 -9964 -2102 -9908
rect -2078 -9964 -2022 -9908
rect -10821 -10064 -10765 -10008
rect -10741 -10064 -10685 -10008
rect -10661 -10064 -10605 -10008
rect -2238 -10064 -2182 -10008
rect -2158 -10064 -2102 -10008
rect -2078 -10064 -2022 -10008
rect -10821 -10164 -10765 -10108
rect -10741 -10164 -10685 -10108
rect -10661 -10164 -10605 -10108
rect -2238 -10164 -2182 -10108
rect -2158 -10164 -2102 -10108
rect -2078 -10164 -2022 -10108
rect -10821 -10264 -10765 -10208
rect -10741 -10264 -10685 -10208
rect -10661 -10264 -10605 -10208
rect -2238 -10264 -2182 -10208
rect -2158 -10264 -2102 -10208
rect -2078 -10264 -2022 -10208
rect 6929 -10095 6985 -10039
rect 7009 -10095 7065 -10039
rect 7089 -10095 7145 -10039
rect 18439 -10095 18495 -10039
rect 18519 -10095 18575 -10039
rect 18599 -10095 18655 -10039
rect 6929 -10195 6985 -10139
rect 7009 -10195 7065 -10139
rect 7089 -10195 7145 -10139
rect 18439 -10195 18495 -10139
rect 18519 -10195 18575 -10139
rect 18599 -10195 18655 -10139
rect 6929 -10295 6985 -10239
rect 7009 -10295 7065 -10239
rect 7089 -10295 7145 -10239
rect 18439 -10295 18495 -10239
rect 18519 -10295 18575 -10239
rect 18599 -10295 18655 -10239
rect 6929 -10395 6985 -10339
rect 7009 -10395 7065 -10339
rect 7089 -10395 7145 -10339
rect 18439 -10395 18495 -10339
rect 18519 -10395 18575 -10339
rect 18599 -10395 18655 -10339
rect 6933 -10495 6989 -10439
rect 7013 -10495 7069 -10439
rect 7093 -10495 7149 -10439
rect 18435 -10495 18491 -10439
rect 18515 -10495 18571 -10439
rect 18595 -10495 18651 -10439
rect -7609 -10682 -7553 -10626
rect -7529 -10682 -7473 -10626
rect -7449 -10682 -7393 -10626
rect -3158 -10682 -3102 -10626
rect -3078 -10682 -3022 -10626
rect -2998 -10682 -2942 -10626
rect -7609 -10782 -7553 -10726
rect -7529 -10782 -7473 -10726
rect -7449 -10782 -7393 -10726
rect -3158 -10782 -3102 -10726
rect -3078 -10782 -3022 -10726
rect -2998 -10782 -2942 -10726
rect -1690 -10749 -1634 -10693
rect -1610 -10749 -1554 -10693
rect -1530 -10749 -1474 -10693
rect 3204 -10749 3260 -10693
rect 3284 -10749 3340 -10693
rect 3364 -10749 3420 -10693
rect 8005 -10749 8061 -10693
rect 8085 -10749 8141 -10693
rect 8165 -10749 8221 -10693
rect 17364 -10749 17420 -10693
rect 17444 -10749 17500 -10693
rect 17524 -10749 17580 -10693
rect -7609 -10882 -7553 -10826
rect -7529 -10882 -7473 -10826
rect -7449 -10882 -7393 -10826
rect -3158 -10882 -3102 -10826
rect -3078 -10882 -3022 -10826
rect -2998 -10882 -2942 -10826
rect -7609 -10982 -7553 -10926
rect -7529 -10982 -7473 -10926
rect -7449 -10982 -7393 -10926
rect -3158 -10982 -3102 -10926
rect -3078 -10982 -3022 -10926
rect -2998 -10982 -2942 -10926
rect -1690 -11066 -1634 -11010
rect -1610 -11066 -1554 -11010
rect -1530 -11066 -1474 -11010
rect 3204 -11066 3260 -11010
rect 3284 -11066 3340 -11010
rect 3364 -11066 3420 -11010
rect 7517 -11066 7573 -11010
rect 7597 -11066 7653 -11010
rect 7677 -11066 7733 -11010
rect 12672 -11067 12728 -11011
rect 12752 -11067 12808 -11011
rect 12832 -11067 12888 -11011
rect 17851 -11066 17907 -11010
rect 17931 -11066 17987 -11010
rect 18011 -11066 18067 -11010
rect -1690 -12146 -1634 -12090
rect -1610 -12146 -1554 -12090
rect -1530 -12146 -1474 -12090
rect 3204 -12146 3260 -12090
rect 3284 -12146 3340 -12090
rect 3364 -12146 3420 -12090
rect 7517 -12146 7573 -12090
rect 7597 -12146 7653 -12090
rect 7677 -12146 7733 -12090
rect 12672 -12146 12728 -12090
rect 12752 -12146 12808 -12090
rect 12832 -12146 12888 -12090
rect 17851 -12146 17907 -12090
rect 17931 -12146 17987 -12090
rect 18011 -12146 18067 -12090
rect -1690 -12464 -1634 -12408
rect -1610 -12464 -1554 -12408
rect -1530 -12464 -1474 -12408
rect 3204 -12464 3260 -12408
rect 3284 -12464 3340 -12408
rect 3364 -12464 3420 -12408
rect 8005 -12464 8061 -12408
rect 8085 -12464 8141 -12408
rect 8165 -12464 8221 -12408
rect 17364 -12464 17420 -12408
rect 17444 -12464 17500 -12408
rect 17524 -12464 17580 -12408
rect -3158 -13421 -3102 -13365
rect -3078 -13421 -3022 -13365
rect -2998 -13421 -2942 -13365
rect 220 -13421 276 -13365
rect 300 -13421 356 -13365
rect 380 -13421 436 -13365
rect 1301 -13421 1357 -13365
rect 1381 -13421 1437 -13365
rect 1461 -13421 1517 -13365
rect 2422 -13421 2478 -13365
rect 2502 -13421 2558 -13365
rect 2582 -13421 2638 -13365
rect -3158 -13521 -3102 -13465
rect -3078 -13521 -3022 -13465
rect -2998 -13521 -2942 -13465
rect 220 -13521 276 -13465
rect 300 -13521 356 -13465
rect 380 -13521 436 -13465
rect 1301 -13521 1357 -13465
rect 1381 -13521 1437 -13465
rect 1461 -13521 1517 -13465
rect 2422 -13521 2478 -13465
rect 2502 -13521 2558 -13465
rect 2582 -13521 2638 -13465
rect -3158 -13621 -3102 -13565
rect -3078 -13621 -3022 -13565
rect -2998 -13621 -2942 -13565
rect 220 -13621 276 -13565
rect 300 -13621 356 -13565
rect 380 -13621 436 -13565
rect 1301 -13621 1357 -13565
rect 1381 -13621 1437 -13565
rect 1461 -13621 1517 -13565
rect 2422 -13621 2478 -13565
rect 2502 -13621 2558 -13565
rect 2582 -13621 2638 -13565
rect -3158 -13721 -3102 -13665
rect -3078 -13721 -3022 -13665
rect -2998 -13721 -2942 -13665
rect 220 -13721 276 -13665
rect 300 -13721 356 -13665
rect 380 -13721 436 -13665
rect 1301 -13721 1357 -13665
rect 1381 -13721 1437 -13665
rect 1461 -13721 1517 -13665
rect 2422 -13721 2478 -13665
rect 2502 -13721 2558 -13665
rect 2582 -13721 2638 -13665
rect 9662 -13540 9718 -13484
rect 9742 -13540 9798 -13484
rect 9822 -13540 9878 -13484
rect 13201 -13540 13257 -13484
rect 13281 -13540 13337 -13484
rect 13361 -13540 13417 -13484
rect 15660 -13540 15716 -13484
rect 15740 -13540 15796 -13484
rect 15820 -13540 15876 -13484
rect 9662 -13640 9718 -13584
rect 9742 -13640 9798 -13584
rect 9822 -13640 9878 -13584
rect 13201 -13640 13257 -13584
rect 13281 -13640 13337 -13584
rect 13361 -13640 13417 -13584
rect 15660 -13640 15716 -13584
rect 15740 -13640 15796 -13584
rect 15820 -13640 15876 -13584
rect 9662 -13740 9718 -13684
rect 9742 -13740 9798 -13684
rect 9822 -13740 9878 -13684
rect 13201 -13740 13257 -13684
rect 13281 -13740 13337 -13684
rect 13361 -13740 13417 -13684
rect 15660 -13740 15716 -13684
rect 15740 -13740 15796 -13684
rect 15820 -13740 15876 -13684
rect 9662 -13840 9718 -13784
rect 9742 -13840 9798 -13784
rect 9822 -13840 9878 -13784
rect 13201 -13840 13257 -13784
rect 13281 -13840 13337 -13784
rect 13361 -13840 13417 -13784
rect 15660 -13840 15716 -13784
rect 15740 -13840 15796 -13784
rect 15820 -13840 15876 -13784
rect -2238 -14081 -2182 -14025
rect -2158 -14081 -2102 -14025
rect -2078 -14081 -2022 -14025
rect -901 -14081 -845 -14025
rect -821 -14081 -765 -14025
rect -741 -14081 -685 -14025
rect 3759 -14081 3815 -14025
rect 3839 -14081 3895 -14025
rect 3919 -14081 3975 -14025
rect -2238 -14181 -2182 -14125
rect -2158 -14181 -2102 -14125
rect -2078 -14181 -2022 -14125
rect -901 -14181 -845 -14125
rect -821 -14181 -765 -14125
rect -741 -14181 -685 -14125
rect 3759 -14181 3815 -14125
rect 3839 -14181 3895 -14125
rect 3919 -14181 3975 -14125
rect -2238 -14281 -2182 -14225
rect -2158 -14281 -2102 -14225
rect -2078 -14281 -2022 -14225
rect -901 -14281 -845 -14225
rect -821 -14281 -765 -14225
rect -741 -14281 -685 -14225
rect 3759 -14281 3815 -14225
rect 3839 -14281 3895 -14225
rect 3919 -14281 3975 -14225
rect -2238 -14381 -2182 -14325
rect -2158 -14381 -2102 -14325
rect -2078 -14381 -2022 -14325
rect -901 -14381 -845 -14325
rect -821 -14381 -765 -14325
rect -741 -14381 -685 -14325
rect 3759 -14381 3815 -14325
rect 3839 -14381 3895 -14325
rect 3919 -14381 3975 -14325
rect 12121 -14096 12177 -14040
rect 12201 -14096 12257 -14040
rect 12281 -14096 12337 -14040
rect 13201 -14096 13257 -14040
rect 13281 -14096 13337 -14040
rect 13361 -14096 13417 -14040
rect 12121 -14196 12177 -14140
rect 12201 -14196 12257 -14140
rect 12281 -14196 12337 -14140
rect 13201 -14196 13257 -14140
rect 13281 -14196 13337 -14140
rect 13361 -14196 13417 -14140
rect 12121 -14296 12177 -14240
rect 12201 -14296 12257 -14240
rect 12281 -14296 12337 -14240
rect 13201 -14296 13257 -14240
rect 13281 -14296 13337 -14240
rect 13361 -14296 13417 -14240
rect 12121 -14396 12177 -14340
rect 12201 -14396 12257 -14340
rect 12281 -14396 12337 -14340
rect 13201 -14396 13257 -14340
rect 13281 -14396 13337 -14340
rect 13361 -14396 13417 -14340
rect -3457 -15384 -3401 -15328
rect -3377 -15384 -3321 -15328
rect -3297 -15384 -3241 -15328
rect 4938 -15384 4994 -15328
rect 5018 -15384 5074 -15328
rect 5098 -15384 5154 -15328
rect 8444 -15384 8500 -15328
rect 8524 -15384 8580 -15328
rect 8604 -15384 8660 -15328
rect 16838 -15384 16894 -15328
rect 16918 -15384 16974 -15328
rect 16998 -15384 17054 -15328
rect -3457 -15701 -3401 -15645
rect -3377 -15701 -3321 -15645
rect -3297 -15701 -3241 -15645
rect 4938 -15701 4994 -15645
rect 5018 -15701 5074 -15645
rect 5098 -15701 5154 -15645
rect 8444 -15701 8500 -15645
rect 8524 -15701 8580 -15645
rect 8604 -15701 8660 -15645
rect 16838 -15701 16894 -15645
rect 16918 -15701 16974 -15645
rect 16998 -15701 17054 -15645
rect -3457 -16781 -3401 -16725
rect -3377 -16781 -3321 -16725
rect -3297 -16781 -3241 -16725
rect 4938 -16781 4994 -16725
rect 5018 -16781 5074 -16725
rect 5098 -16781 5154 -16725
rect 8444 -16781 8500 -16725
rect 8524 -16781 8580 -16725
rect 8604 -16781 8660 -16725
rect 16838 -16781 16894 -16725
rect 16918 -16781 16974 -16725
rect 16998 -16781 17054 -16725
rect -3457 -17098 -3401 -17042
rect -3377 -17098 -3321 -17042
rect -3297 -17098 -3241 -17042
rect 4938 -17098 4994 -17042
rect 5018 -17098 5074 -17042
rect 5098 -17098 5154 -17042
rect 8444 -17098 8500 -17042
rect 8524 -17098 8580 -17042
rect 8604 -17098 8660 -17042
rect 16838 -17098 16894 -17042
rect 16918 -17098 16974 -17042
rect 16998 -17098 17054 -17042
<< metal3 >>
rect -25759 10488 -25459 10510
rect -25759 10432 -25719 10488
rect -25663 10432 -25639 10488
rect -25583 10432 -25559 10488
rect -25503 10432 -25459 10488
rect -25759 10168 -25459 10432
rect -25759 10112 -25719 10168
rect -25663 10112 -25639 10168
rect -25583 10112 -25559 10168
rect -25503 10112 -25459 10168
rect -25759 8841 -25459 10112
rect -25759 8785 -25719 8841
rect -25663 8785 -25639 8841
rect -25583 8785 -25559 8841
rect -25503 8785 -25459 8841
rect -25759 8509 -25459 8785
rect -25759 8453 -25719 8509
rect -25663 8453 -25639 8509
rect -25583 8453 -25559 8509
rect -25503 8453 -25459 8509
rect -25759 5615 -25459 8453
rect -25759 5559 -25719 5615
rect -25663 5559 -25639 5615
rect -25583 5559 -25559 5615
rect -25503 5559 -25459 5615
rect -6617 10488 -6317 10510
rect -6617 10432 -6573 10488
rect -6517 10432 -6493 10488
rect -6437 10432 -6413 10488
rect -6357 10432 -6317 10488
rect -6617 10168 -6317 10432
rect -6617 10112 -6573 10168
rect -6517 10112 -6493 10168
rect -6437 10112 -6413 10168
rect -6357 10112 -6317 10168
rect -6617 8841 -6317 10112
rect -6617 8785 -6573 8841
rect -6517 8785 -6493 8841
rect -6437 8785 -6413 8841
rect -6357 8785 -6317 8841
rect -6617 8509 -6317 8785
rect -6617 8453 -6573 8509
rect -6517 8453 -6493 8509
rect -6437 8453 -6413 8509
rect -6357 8453 -6317 8509
rect -6617 5615 -6317 8453
rect -25759 5283 -25459 5559
rect -25759 5227 -25719 5283
rect -25663 5227 -25639 5283
rect -25583 5227 -25559 5283
rect -25503 5227 -25459 5283
rect -25759 3956 -25459 5227
rect -25759 3900 -25719 3956
rect -25663 3900 -25639 3956
rect -25583 3900 -25559 3956
rect -25503 3900 -25459 3956
rect -25759 3636 -25459 3900
rect -25759 3580 -25719 3636
rect -25663 3580 -25639 3636
rect -25583 3580 -25559 3636
rect -25503 3580 -25459 3636
rect -25759 3558 -25459 3580
rect -24359 2140 -24059 3817
rect -24359 2084 -24315 2140
rect -24259 2084 -24235 2140
rect -24179 2084 -24155 2140
rect -24099 2084 -24059 2140
rect -24359 2040 -24059 2084
rect -24359 1984 -24315 2040
rect -24259 1984 -24235 2040
rect -24179 1984 -24155 2040
rect -24099 1984 -24059 2040
rect -24359 1962 -24059 1984
rect -25354 1791 -25054 1813
rect -25354 1735 -25310 1791
rect -25254 1735 -25230 1791
rect -25174 1735 -25150 1791
rect -25094 1735 -25054 1791
rect -25354 1691 -25054 1735
rect -25354 1635 -25310 1691
rect -25254 1635 -25230 1691
rect -25174 1635 -25150 1691
rect -25094 1635 -25054 1691
rect -26532 294 -26232 316
rect -26532 238 -26492 294
rect -26436 238 -26412 294
rect -26356 238 -26332 294
rect -26276 238 -26232 294
rect -27032 -27 -26732 -5
rect -27032 -83 -26992 -27
rect -26936 -83 -26912 -27
rect -26856 -83 -26832 -27
rect -26776 -83 -26732 -27
rect -27032 -1365 -26732 -83
rect -27032 -1421 -26992 -1365
rect -26936 -1421 -26912 -1365
rect -26856 -1421 -26832 -1365
rect -26776 -1421 -26732 -1365
rect -27032 -4900 -26732 -1421
rect -27032 -4956 -26992 -4900
rect -26936 -4956 -26912 -4900
rect -26856 -4956 -26832 -4900
rect -26776 -4956 -26732 -4900
rect -27032 -6238 -26732 -4956
rect -27032 -6294 -26992 -6238
rect -26936 -6294 -26912 -6238
rect -26856 -6294 -26832 -6238
rect -26776 -6294 -26732 -6238
rect -27032 -6316 -26732 -6294
rect -26532 -1685 -26232 238
rect -25354 -62 -25054 1635
rect -21151 1791 -20851 3468
rect -21151 1735 -21107 1791
rect -21051 1735 -21027 1791
rect -20971 1735 -20947 1791
rect -20891 1735 -20851 1791
rect -21151 1691 -20851 1735
rect -21151 1635 -21107 1691
rect -21051 1635 -21027 1691
rect -20971 1635 -20947 1691
rect -20891 1635 -20851 1691
rect -21151 -62 -20851 1635
rect -20001 1791 -19701 3468
rect -16793 2140 -16493 3817
rect -16793 2084 -16749 2140
rect -16693 2084 -16669 2140
rect -16613 2084 -16589 2140
rect -16533 2084 -16493 2140
rect -16793 2040 -16493 2084
rect -16793 1984 -16749 2040
rect -16693 1984 -16669 2040
rect -16613 1984 -16589 2040
rect -16533 1984 -16493 2040
rect -16793 1962 -16493 1984
rect -15642 2140 -15342 3817
rect -15642 2084 -15598 2140
rect -15542 2084 -15518 2140
rect -15462 2084 -15438 2140
rect -15382 2084 -15342 2140
rect -15642 2040 -15342 2084
rect -15642 1984 -15598 2040
rect -15542 1984 -15518 2040
rect -15462 1984 -15438 2040
rect -15382 1984 -15342 2040
rect -20001 1735 -19957 1791
rect -19901 1735 -19877 1791
rect -19821 1735 -19797 1791
rect -19741 1735 -19701 1791
rect -20001 1691 -19701 1735
rect -20001 1635 -19957 1691
rect -19901 1635 -19877 1691
rect -19821 1635 -19797 1691
rect -19741 1635 -19701 1691
rect -20001 1613 -19701 1635
rect -16943 1791 -16643 1813
rect -16943 1735 -16899 1791
rect -16843 1735 -16819 1791
rect -16763 1735 -16739 1791
rect -16683 1735 -16643 1791
rect -16943 1691 -16643 1735
rect -16943 1635 -16899 1691
rect -16843 1635 -16819 1691
rect -16763 1635 -16739 1691
rect -16683 1635 -16643 1691
rect -16943 -62 -16643 1635
rect -15642 -874 -15342 1984
rect -12434 1791 -12134 3468
rect -11284 2497 -10984 5598
rect -6617 5559 -6573 5615
rect -6517 5559 -6493 5615
rect -6437 5559 -6413 5615
rect -6357 5559 -6317 5615
rect -6617 5283 -6317 5559
rect -6617 5227 -6573 5283
rect -6517 5227 -6493 5283
rect -6437 5227 -6413 5283
rect -6357 5227 -6317 5283
rect -6617 3956 -6317 5227
rect -6617 3900 -6573 3956
rect -6517 3900 -6493 3956
rect -6437 3900 -6413 3956
rect -6357 3900 -6317 3956
rect -11284 2441 -11240 2497
rect -11184 2441 -11160 2497
rect -11104 2441 -11080 2497
rect -11024 2441 -10984 2497
rect -11284 2397 -10984 2441
rect -11284 2341 -11240 2397
rect -11184 2341 -11160 2397
rect -11104 2341 -11080 2397
rect -11024 2341 -10984 2397
rect -11284 2319 -10984 2341
rect -10575 2497 -10275 2519
rect -10575 2441 -10531 2497
rect -10475 2441 -10451 2497
rect -10395 2441 -10371 2497
rect -10315 2441 -10275 2497
rect -10575 2397 -10275 2441
rect -10575 2341 -10531 2397
rect -10475 2341 -10451 2397
rect -10395 2341 -10371 2397
rect -10315 2341 -10275 2397
rect -12434 1735 -12390 1791
rect -12334 1735 -12310 1791
rect -12254 1735 -12230 1791
rect -12174 1735 -12134 1791
rect -12434 1691 -12134 1735
rect -12434 1635 -12390 1691
rect -12334 1635 -12310 1691
rect -12254 1635 -12230 1691
rect -12174 1635 -12134 1691
rect -12434 1613 -12134 1635
rect -11444 2140 -11144 2162
rect -11444 2084 -11400 2140
rect -11344 2084 -11320 2140
rect -11264 2084 -11240 2140
rect -11184 2084 -11144 2140
rect -11444 2040 -11144 2084
rect -11444 1984 -11400 2040
rect -11344 1984 -11320 2040
rect -11264 1984 -11240 2040
rect -11184 1984 -11144 2040
rect -11444 307 -11144 1984
rect -10575 1791 -10275 2341
rect -8076 2140 -7776 3817
rect -6617 3636 -6317 3900
rect -6617 3580 -6573 3636
rect -6517 3580 -6493 3636
rect -6437 3580 -6413 3636
rect -6357 3580 -6317 3636
rect -6617 3558 -6317 3580
rect -4750 10488 -4450 10510
rect -4750 10432 -4706 10488
rect -4650 10432 -4626 10488
rect -4570 10432 -4546 10488
rect -4490 10432 -4450 10488
rect -4750 8509 -4450 10432
rect -4750 8453 -4706 8509
rect -4650 8453 -4626 8509
rect -4570 8453 -4546 8509
rect -4490 8453 -4450 8509
rect -4750 5614 -4450 8453
rect 5753 10488 6053 10510
rect 5753 10432 5793 10488
rect 5849 10432 5873 10488
rect 5929 10432 5953 10488
rect 6009 10432 6053 10488
rect 5753 10167 6053 10432
rect 5753 10111 5793 10167
rect 5849 10111 5873 10167
rect 5929 10111 5953 10167
rect 6009 10111 6053 10167
rect 5753 8841 6053 10111
rect 5753 8785 5793 8841
rect 5849 8785 5873 8841
rect 5929 8785 5953 8841
rect 6009 8785 6053 8841
rect 5753 8509 6053 8785
rect 5753 8453 5793 8509
rect 5849 8453 5873 8509
rect 5929 8453 5953 8509
rect 6009 8453 6053 8509
rect -4750 5558 -4706 5614
rect -4650 5558 -4626 5614
rect -4570 5558 -4546 5614
rect -4490 5558 -4450 5614
rect -4750 5294 -4450 5558
rect -4750 5238 -4706 5294
rect -4650 5238 -4626 5294
rect -4570 5238 -4546 5294
rect -4490 5238 -4450 5294
rect -4750 3956 -4450 5238
rect -4750 3900 -4706 3956
rect -4650 3900 -4626 3956
rect -4570 3900 -4546 3956
rect -4490 3900 -4450 3956
rect -4750 3636 -4450 3900
rect -4750 3580 -4706 3636
rect -4650 3580 -4626 3636
rect -4570 3580 -4546 3636
rect -4490 3580 -4450 3636
rect -4750 3558 -4450 3580
rect -8076 2084 -8032 2140
rect -7976 2084 -7952 2140
rect -7896 2084 -7872 2140
rect -7816 2084 -7776 2140
rect -8076 2040 -7776 2084
rect -8076 1984 -8032 2040
rect -7976 1984 -7952 2040
rect -7896 1984 -7872 2040
rect -7816 1984 -7776 2040
rect -8076 1962 -7776 1984
rect -7231 2140 -6931 2162
rect -7231 2084 -7187 2140
rect -7131 2084 -7107 2140
rect -7051 2084 -7027 2140
rect -6971 2084 -6931 2140
rect -7231 2040 -6931 2084
rect -7231 1984 -7187 2040
rect -7131 1984 -7107 2040
rect -7051 1984 -7027 2040
rect -6971 1984 -6931 2040
rect -10575 1735 -10531 1791
rect -10475 1735 -10451 1791
rect -10395 1735 -10371 1791
rect -10315 1735 -10275 1791
rect -10575 1691 -10275 1735
rect -10575 1635 -10531 1691
rect -10475 1635 -10451 1691
rect -10395 1635 -10371 1691
rect -10315 1635 -10275 1691
rect -10575 1613 -10275 1635
rect -7231 287 -6931 1984
rect -3676 1808 -3376 1830
rect -3676 1752 -3636 1808
rect -3580 1752 -3556 1808
rect -3500 1752 -3476 1808
rect -3420 1752 -3376 1808
rect -3676 1708 -3376 1752
rect -3676 1652 -3636 1708
rect -3580 1652 -3556 1708
rect -3500 1652 -3476 1708
rect -3420 1652 -3376 1708
rect -3676 1608 -3376 1652
rect -3676 1552 -3636 1608
rect -3580 1552 -3556 1608
rect -3500 1552 -3476 1608
rect -3420 1552 -3376 1608
rect -3676 1508 -3376 1552
rect -3676 1452 -3636 1508
rect -3580 1452 -3556 1508
rect -3500 1452 -3476 1508
rect -3420 1452 -3376 1508
rect -6105 294 -5805 316
rect -6105 238 -6061 294
rect -6005 238 -5981 294
rect -5925 238 -5901 294
rect -5845 238 -5805 294
rect -26532 -1741 -26492 -1685
rect -26436 -1741 -26412 -1685
rect -26356 -1741 -26332 -1685
rect -26276 -1741 -26232 -1685
rect -26532 -4580 -26232 -1741
rect -26532 -4636 -26492 -4580
rect -26436 -4636 -26412 -4580
rect -26356 -4636 -26332 -4580
rect -26276 -4636 -26232 -4580
rect -26532 -6558 -26232 -4636
rect -6105 -1685 -5805 238
rect -4750 294 -4450 316
rect -4750 238 -4706 294
rect -4650 238 -4626 294
rect -4570 238 -4546 294
rect -4490 238 -4450 294
rect -6105 -1741 -6061 -1685
rect -6005 -1741 -5981 -1685
rect -5925 -1741 -5901 -1685
rect -5845 -1741 -5805 -1685
rect -6105 -4580 -5805 -1741
rect -6105 -4636 -6061 -4580
rect -6005 -4636 -5981 -4580
rect -5925 -4636 -5901 -4580
rect -5845 -4636 -5805 -4580
rect -26532 -6614 -26492 -6558
rect -26436 -6614 -26412 -6558
rect -26356 -6614 -26332 -6558
rect -26276 -6614 -26232 -6558
rect -26532 -6636 -26232 -6614
rect -24932 -8018 -24632 -5454
rect -24932 -8074 -24892 -8018
rect -24836 -8074 -24812 -8018
rect -24756 -8074 -24732 -8018
rect -24676 -8074 -24632 -8018
rect -24932 -8118 -24632 -8074
rect -24932 -8174 -24892 -8118
rect -24836 -8174 -24812 -8118
rect -24756 -8174 -24732 -8118
rect -24676 -8174 -24632 -8118
rect -24932 -8218 -24632 -8174
rect -24932 -8274 -24892 -8218
rect -24836 -8274 -24812 -8218
rect -24756 -8274 -24732 -8218
rect -24676 -8274 -24632 -8218
rect -24932 -8318 -24632 -8274
rect -24932 -8374 -24892 -8318
rect -24836 -8374 -24812 -8318
rect -24756 -8374 -24732 -8318
rect -24676 -8374 -24632 -8318
rect -24932 -8396 -24632 -8374
rect -21724 -8736 -21424 -5739
rect -21724 -8792 -21680 -8736
rect -21624 -8792 -21600 -8736
rect -21544 -8792 -21520 -8736
rect -21464 -8792 -21424 -8736
rect -21724 -8836 -21424 -8792
rect -21724 -8892 -21680 -8836
rect -21624 -8892 -21600 -8836
rect -21544 -8892 -21520 -8836
rect -21464 -8892 -21424 -8836
rect -21724 -8936 -21424 -8892
rect -21724 -8992 -21680 -8936
rect -21624 -8992 -21600 -8936
rect -21544 -8992 -21520 -8936
rect -21464 -8992 -21424 -8936
rect -21724 -9036 -21424 -8992
rect -20574 -8714 -20274 -5739
rect -17366 -8018 -17066 -5454
rect -17366 -8074 -17326 -8018
rect -17270 -8074 -17246 -8018
rect -17190 -8074 -17166 -8018
rect -17110 -8074 -17066 -8018
rect -17366 -8118 -17066 -8074
rect -17366 -8174 -17326 -8118
rect -17270 -8174 -17246 -8118
rect -17190 -8174 -17166 -8118
rect -17110 -8174 -17066 -8118
rect -17366 -8218 -17066 -8174
rect -17366 -8274 -17326 -8218
rect -17270 -8274 -17246 -8218
rect -17190 -8274 -17166 -8218
rect -17110 -8274 -17066 -8218
rect -17366 -8318 -17066 -8274
rect -17366 -8374 -17326 -8318
rect -17270 -8374 -17246 -8318
rect -17190 -8374 -17166 -8318
rect -17110 -8374 -17066 -8318
rect -17366 -8396 -17066 -8374
rect -15220 -8714 -14920 -5908
rect -12012 -8018 -11712 -5117
rect -12012 -8074 -11972 -8018
rect -11916 -8074 -11892 -8018
rect -11836 -8074 -11812 -8018
rect -11756 -8074 -11712 -8018
rect -12012 -8118 -11712 -8074
rect -12012 -8174 -11972 -8118
rect -11916 -8174 -11892 -8118
rect -11836 -8174 -11812 -8118
rect -11756 -8174 -11712 -8118
rect -12012 -8218 -11712 -8174
rect -12012 -8274 -11972 -8218
rect -11916 -8274 -11892 -8218
rect -11836 -8274 -11812 -8218
rect -11756 -8274 -11712 -8218
rect -12012 -8318 -11712 -8274
rect -12012 -8374 -11972 -8318
rect -11916 -8374 -11892 -8318
rect -11836 -8374 -11812 -8318
rect -11756 -8374 -11712 -8318
rect -12012 -8396 -11712 -8374
rect -10861 -8018 -10561 -5117
rect -10861 -8074 -10821 -8018
rect -10765 -8074 -10741 -8018
rect -10685 -8074 -10661 -8018
rect -10605 -8074 -10561 -8018
rect -10861 -8118 -10561 -8074
rect -10861 -8174 -10821 -8118
rect -10765 -8174 -10741 -8118
rect -10685 -8174 -10661 -8118
rect -10605 -8174 -10561 -8118
rect -10861 -8218 -10561 -8174
rect -10861 -8274 -10821 -8218
rect -10765 -8274 -10741 -8218
rect -10685 -8274 -10661 -8218
rect -10605 -8274 -10561 -8218
rect -10861 -8318 -10561 -8274
rect -10861 -8374 -10821 -8318
rect -10765 -8374 -10741 -8318
rect -10685 -8374 -10661 -8318
rect -10605 -8374 -10561 -8318
rect -20574 -8736 -20273 -8714
rect -20574 -8792 -20529 -8736
rect -20473 -8792 -20449 -8736
rect -20393 -8792 -20369 -8736
rect -20313 -8792 -20273 -8736
rect -20574 -8836 -20273 -8792
rect -20574 -8892 -20529 -8836
rect -20473 -8892 -20449 -8836
rect -20393 -8892 -20369 -8836
rect -20313 -8892 -20273 -8836
rect -15220 -8736 -14919 -8714
rect -15220 -8792 -15175 -8736
rect -15119 -8792 -15095 -8736
rect -15039 -8792 -15015 -8736
rect -14959 -8792 -14919 -8736
rect -15220 -8836 -14919 -8792
rect -15220 -8850 -15175 -8836
rect -20574 -8936 -20273 -8892
rect -20574 -8992 -20529 -8936
rect -20473 -8992 -20449 -8936
rect -20393 -8992 -20369 -8936
rect -20313 -8992 -20273 -8936
rect -20574 -9019 -20273 -8992
rect -21724 -9092 -21680 -9036
rect -21624 -9092 -21600 -9036
rect -21544 -9092 -21520 -9036
rect -21464 -9092 -21424 -9036
rect -21724 -9114 -21424 -9092
rect -20573 -9036 -20273 -9019
rect -20573 -9092 -20529 -9036
rect -20473 -9092 -20449 -9036
rect -20393 -9092 -20369 -9036
rect -20313 -9092 -20273 -9036
rect -20573 -9114 -20273 -9092
rect -15219 -8892 -15175 -8850
rect -15119 -8892 -15095 -8836
rect -15039 -8892 -15015 -8836
rect -14959 -8892 -14919 -8836
rect -15219 -8936 -14919 -8892
rect -15219 -8992 -15175 -8936
rect -15119 -8992 -15095 -8936
rect -15039 -8992 -15015 -8936
rect -14959 -8992 -14919 -8936
rect -15219 -9036 -14919 -8992
rect -15219 -9092 -15175 -9036
rect -15119 -9092 -15095 -9036
rect -15039 -9092 -15015 -9036
rect -14959 -9092 -14919 -9036
rect -15219 -9114 -14919 -9092
rect -10861 -9908 -10561 -8374
rect -10861 -9964 -10821 -9908
rect -10765 -9964 -10741 -9908
rect -10685 -9964 -10661 -9908
rect -10605 -9964 -10561 -9908
rect -10861 -10008 -10561 -9964
rect -10861 -10064 -10821 -10008
rect -10765 -10064 -10741 -10008
rect -10685 -10064 -10661 -10008
rect -10605 -10064 -10561 -10008
rect -10861 -10108 -10561 -10064
rect -10861 -10164 -10821 -10108
rect -10765 -10164 -10741 -10108
rect -10685 -10164 -10661 -10108
rect -10605 -10164 -10561 -10108
rect -10861 -10208 -10561 -10164
rect -10861 -10264 -10821 -10208
rect -10765 -10264 -10741 -10208
rect -10685 -10264 -10661 -10208
rect -10605 -10264 -10561 -10208
rect -10861 -10286 -10561 -10264
rect -7653 -8736 -7353 -5908
rect -6105 -6558 -5805 -4636
rect -5606 -27 -5306 -5
rect -5606 -83 -5562 -27
rect -5506 -83 -5482 -27
rect -5426 -83 -5402 -27
rect -5346 -83 -5306 -27
rect -5606 -1365 -5306 -83
rect -5606 -1421 -5562 -1365
rect -5506 -1421 -5482 -1365
rect -5426 -1421 -5402 -1365
rect -5346 -1421 -5306 -1365
rect -5606 -4900 -5306 -1421
rect -5606 -4956 -5562 -4900
rect -5506 -4956 -5482 -4900
rect -5426 -4956 -5402 -4900
rect -5346 -4956 -5306 -4900
rect -5606 -6238 -5306 -4956
rect -5606 -6294 -5562 -6238
rect -5506 -6294 -5482 -6238
rect -5426 -6294 -5402 -6238
rect -5346 -6294 -5306 -6238
rect -5606 -6316 -5306 -6294
rect -4750 -1685 -4450 238
rect -4750 -1741 -4706 -1685
rect -4650 -1741 -4626 -1685
rect -4570 -1741 -4546 -1685
rect -4490 -1741 -4450 -1685
rect -4750 -4580 -4450 -1741
rect -3676 -1775 -3376 1452
rect -3254 1808 -2954 4371
rect -46 2414 254 6237
rect -46 2358 -6 2414
rect 50 2358 74 2414
rect 130 2358 154 2414
rect 210 2358 254 2414
rect -46 2314 254 2358
rect -46 2258 -6 2314
rect 50 2258 74 2314
rect 130 2258 154 2314
rect 210 2258 254 2314
rect -46 2214 254 2258
rect -46 2158 -6 2214
rect 50 2158 74 2214
rect 130 2158 154 2214
rect 210 2158 254 2214
rect -46 2114 254 2158
rect -46 2058 -6 2114
rect 50 2058 74 2114
rect 130 2058 154 2114
rect 210 2058 254 2114
rect -46 2036 254 2058
rect 389 2414 970 2436
rect 389 2358 562 2414
rect 618 2358 642 2414
rect 698 2358 722 2414
rect 778 2358 970 2414
rect 389 2314 970 2358
rect 389 2258 562 2314
rect 618 2258 642 2314
rect 698 2258 722 2314
rect 778 2258 970 2314
rect 389 2214 970 2258
rect 389 2158 562 2214
rect 618 2158 642 2214
rect 698 2158 722 2214
rect 778 2158 970 2214
rect 389 2114 970 2158
rect 389 2058 562 2114
rect 618 2058 642 2114
rect 698 2058 722 2114
rect 778 2058 970 2114
rect -3254 1752 -3214 1808
rect -3158 1752 -3134 1808
rect -3078 1752 -3054 1808
rect -2998 1752 -2954 1808
rect -3254 1708 -2954 1752
rect -3254 1652 -3214 1708
rect -3158 1652 -3134 1708
rect -3078 1652 -3054 1708
rect -2998 1652 -2954 1708
rect -3254 1608 -2954 1652
rect -3254 1552 -3214 1608
rect -3158 1552 -3134 1608
rect -3078 1552 -3054 1608
rect -2998 1552 -2954 1608
rect -3254 1508 -2954 1552
rect -3254 1452 -3214 1508
rect -3158 1452 -3134 1508
rect -3078 1452 -3054 1508
rect -2998 1452 -2954 1508
rect -3254 1430 -2954 1452
rect 389 522 970 2058
rect 1104 2414 1404 6237
rect 5753 5614 6053 8453
rect 5753 5558 5793 5614
rect 5849 5558 5873 5614
rect 5929 5558 5953 5614
rect 6009 5558 6053 5614
rect 5753 5288 6053 5558
rect 5753 5232 5793 5288
rect 5849 5232 5873 5288
rect 5929 5232 5953 5288
rect 6009 5232 6053 5288
rect 1104 2358 1144 2414
rect 1200 2358 1224 2414
rect 1280 2358 1304 2414
rect 1360 2358 1404 2414
rect 1104 2314 1404 2358
rect 1104 2258 1144 2314
rect 1200 2258 1224 2314
rect 1280 2258 1304 2314
rect 1360 2258 1404 2314
rect 1104 2214 1404 2258
rect 1104 2158 1144 2214
rect 1200 2158 1224 2214
rect 1280 2158 1304 2214
rect 1360 2158 1404 2214
rect 1104 2114 1404 2158
rect 1104 2058 1144 2114
rect 1200 2058 1224 2114
rect 1280 2058 1304 2114
rect 1360 2058 1404 2114
rect 1104 2036 1404 2058
rect 4312 1808 4612 4371
rect 5753 3956 6053 5232
rect 5753 3900 5793 3956
rect 5849 3900 5873 3956
rect 5929 3900 5953 3956
rect 6009 3900 6053 3956
rect 5753 3636 6053 3900
rect 5753 3580 5793 3636
rect 5849 3580 5873 3636
rect 5929 3580 5953 3636
rect 6009 3580 6053 3636
rect 4312 1752 4352 1808
rect 4408 1752 4432 1808
rect 4488 1752 4512 1808
rect 4568 1752 4612 1808
rect 4312 1708 4612 1752
rect 4312 1652 4352 1708
rect 4408 1652 4432 1708
rect 4488 1652 4512 1708
rect 4568 1652 4612 1708
rect 4312 1608 4612 1652
rect 4312 1552 4352 1608
rect 4408 1552 4432 1608
rect 4488 1552 4512 1608
rect 4568 1552 4612 1608
rect 4312 1508 4612 1552
rect 4312 1452 4352 1508
rect 4408 1452 4432 1508
rect 4488 1452 4512 1508
rect 4568 1452 4612 1508
rect 4312 1430 4612 1452
rect 4735 1808 5035 1830
rect 4735 1752 4775 1808
rect 4831 1752 4855 1808
rect 4911 1752 4935 1808
rect 4991 1752 5035 1808
rect 4735 1708 5035 1752
rect 4735 1652 4775 1708
rect 4831 1652 4855 1708
rect 4911 1652 4935 1708
rect 4991 1652 5035 1708
rect 4735 1608 5035 1652
rect 4735 1552 4775 1608
rect 4831 1552 4855 1608
rect 4911 1552 4935 1608
rect 4991 1552 5035 1608
rect 4735 1508 5035 1552
rect 4735 1452 4775 1508
rect 4831 1452 4855 1508
rect 4911 1452 4935 1508
rect 4991 1452 5035 1508
rect 4735 -1775 5035 1452
rect 5753 1331 6053 3580
rect 5753 1275 5793 1331
rect 5849 1275 5873 1331
rect 5929 1275 5953 1331
rect 6009 1275 6053 1331
rect 5753 1231 6053 1275
rect 5753 1175 5793 1231
rect 5849 1175 5873 1231
rect 5929 1175 5953 1231
rect 6009 1175 6053 1231
rect 5753 1131 6053 1175
rect 5753 1075 5793 1131
rect 5849 1075 5873 1131
rect 5929 1075 5953 1131
rect 6009 1075 6053 1131
rect 5753 1031 6053 1075
rect 5753 975 5793 1031
rect 5849 975 5873 1031
rect 5929 975 5953 1031
rect 6009 975 6053 1031
rect 5753 953 6053 975
rect 6889 10488 7189 10510
rect 6889 10432 6929 10488
rect 6985 10432 7009 10488
rect 7065 10432 7089 10488
rect 7145 10432 7189 10488
rect 6889 10167 7189 10432
rect 6889 10111 6929 10167
rect 6985 10111 7009 10167
rect 7065 10111 7089 10167
rect 7145 10111 7189 10167
rect 6889 8841 7189 10111
rect 6889 8785 6929 8841
rect 6985 8785 7009 8841
rect 7065 8785 7089 8841
rect 7145 8785 7189 8841
rect 6889 8509 7189 8785
rect 6889 8453 6929 8509
rect 6985 8453 7009 8509
rect 7065 8453 7089 8509
rect 7145 8453 7189 8509
rect 6889 5614 7189 8453
rect 6889 5558 6929 5614
rect 6985 5558 7009 5614
rect 7065 5558 7089 5614
rect 7145 5558 7189 5614
rect 6889 5288 7189 5558
rect 6889 5232 6929 5288
rect 6985 5232 7009 5288
rect 7065 5232 7089 5288
rect 7145 5232 7189 5288
rect 6889 3956 7189 5232
rect 6889 3900 6929 3956
rect 6985 3900 7009 3956
rect 7065 3900 7089 3956
rect 7145 3900 7189 3956
rect 6889 3636 7189 3900
rect 9816 9590 10116 10510
rect 9816 9534 9856 9590
rect 9912 9534 9936 9590
rect 9992 9534 10016 9590
rect 10072 9534 10116 9590
rect 9816 8077 10116 9534
rect 9816 8021 9856 8077
rect 9912 8021 9936 8077
rect 9992 8021 10016 8077
rect 10072 8021 10116 8077
rect 9816 6046 10116 8021
rect 9816 5990 9856 6046
rect 9912 5990 9936 6046
rect 9992 5990 10016 6046
rect 10072 5990 10116 6046
rect 9816 4534 10116 5990
rect 9816 4478 9856 4534
rect 9912 4478 9936 4534
rect 9992 4478 10016 4534
rect 10072 4478 10116 4534
rect 6889 3580 6929 3636
rect 6985 3580 7009 3636
rect 7065 3580 7089 3636
rect 7145 3580 7189 3636
rect 6889 1331 7189 3580
rect 6889 1275 6929 1331
rect 6985 1275 7009 1331
rect 7065 1275 7089 1331
rect 7145 1275 7189 1331
rect 6889 1231 7189 1275
rect 6889 1175 6929 1231
rect 6985 1175 7009 1231
rect 7065 1175 7089 1231
rect 7145 1175 7189 1231
rect 6889 1131 7189 1175
rect 6889 1075 6929 1131
rect 6985 1075 7009 1131
rect 7065 1075 7089 1131
rect 7145 1075 7189 1131
rect 6889 1031 7189 1075
rect 6889 975 6929 1031
rect 6985 975 7009 1031
rect 7065 975 7089 1031
rect 7145 975 7189 1031
rect 5753 294 6053 316
rect 5753 238 5793 294
rect 5849 238 5873 294
rect 5929 238 5953 294
rect 6009 238 6053 294
rect 5753 -1685 6053 238
rect 5753 -1741 5793 -1685
rect 5849 -1741 5873 -1685
rect 5929 -1741 5953 -1685
rect 6009 -1741 6053 -1685
rect -4750 -4636 -4706 -4580
rect -4650 -4636 -4626 -4580
rect -4570 -4636 -4546 -4580
rect -4490 -4636 -4450 -4580
rect -4750 -4900 -4450 -4636
rect -4750 -4956 -4706 -4900
rect -4650 -4956 -4626 -4900
rect -4570 -4956 -4546 -4900
rect -4490 -4956 -4450 -4900
rect -4750 -6238 -4450 -4956
rect 5753 -4580 6053 -1741
rect 5753 -4636 5793 -4580
rect 5849 -4636 5873 -4580
rect 5929 -4636 5953 -4580
rect 6009 -4636 6053 -4580
rect 5753 -4900 6053 -4636
rect 5753 -4956 5793 -4900
rect 5849 -4956 5873 -4900
rect 5929 -4956 5953 -4900
rect 6009 -4956 6053 -4900
rect -4750 -6294 -4706 -6238
rect -4650 -6294 -4626 -6238
rect -4570 -6294 -4546 -6238
rect -4490 -6294 -4450 -6238
rect -6105 -6614 -6061 -6558
rect -6005 -6614 -5981 -6558
rect -5925 -6614 -5901 -6558
rect -5845 -6614 -5805 -6558
rect -6105 -6636 -5805 -6614
rect -4750 -6558 -4450 -6294
rect -4750 -6614 -4706 -6558
rect -4650 -6614 -4626 -6558
rect -4570 -6614 -4546 -6558
rect -4490 -6614 -4450 -6558
rect -4750 -6636 -4450 -6614
rect -7653 -8792 -7609 -8736
rect -7553 -8792 -7529 -8736
rect -7473 -8792 -7449 -8736
rect -7393 -8792 -7353 -8736
rect -7653 -8836 -7353 -8792
rect -7653 -8892 -7609 -8836
rect -7553 -8892 -7529 -8836
rect -7473 -8892 -7449 -8836
rect -7393 -8892 -7353 -8836
rect -7653 -8936 -7353 -8892
rect -7653 -8992 -7609 -8936
rect -7553 -8992 -7529 -8936
rect -7473 -8992 -7449 -8936
rect -7393 -8992 -7353 -8936
rect -7653 -9036 -7353 -8992
rect -7653 -9092 -7609 -9036
rect -7553 -9092 -7529 -9036
rect -7473 -9092 -7449 -9036
rect -7393 -9092 -7353 -9036
rect -7653 -10626 -7353 -9092
rect -3254 -8899 -2954 -6102
rect -46 -8349 254 -5448
rect -46 -8405 -6 -8349
rect 50 -8405 74 -8349
rect 130 -8405 154 -8349
rect 210 -8405 254 -8349
rect -46 -8449 254 -8405
rect -46 -8505 -6 -8449
rect 50 -8505 74 -8449
rect 130 -8505 154 -8449
rect 210 -8505 254 -8449
rect -46 -8549 254 -8505
rect -46 -8605 -6 -8549
rect 50 -8605 74 -8549
rect 130 -8605 154 -8549
rect 210 -8605 254 -8549
rect -46 -8649 254 -8605
rect -46 -8705 -6 -8649
rect 50 -8705 74 -8649
rect 130 -8705 154 -8649
rect 210 -8705 254 -8649
rect -46 -8728 254 -8705
rect 1104 -8349 1404 -5448
rect 1104 -8405 1144 -8349
rect 1200 -8405 1224 -8349
rect 1280 -8405 1304 -8349
rect 1360 -8405 1404 -8349
rect 1104 -8449 1404 -8405
rect 1104 -8505 1144 -8449
rect 1200 -8505 1224 -8449
rect 1280 -8505 1304 -8449
rect 1360 -8505 1404 -8449
rect 1104 -8549 1404 -8505
rect 1104 -8605 1144 -8549
rect 1200 -8605 1224 -8549
rect 1280 -8605 1304 -8549
rect 1360 -8605 1404 -8549
rect 1104 -8649 1404 -8605
rect 1104 -8705 1144 -8649
rect 1200 -8705 1224 -8649
rect 1280 -8705 1304 -8649
rect 1360 -8705 1404 -8649
rect 1104 -8728 1404 -8705
rect 1950 -8349 2250 -8327
rect 1950 -8405 1990 -8349
rect 2046 -8405 2070 -8349
rect 2126 -8405 2150 -8349
rect 2206 -8405 2250 -8349
rect 1950 -8449 2250 -8405
rect 1950 -8505 1990 -8449
rect 2046 -8505 2070 -8449
rect 2126 -8505 2150 -8449
rect 2206 -8505 2250 -8449
rect 1950 -8549 2250 -8505
rect 1950 -8605 1990 -8549
rect 2046 -8605 2070 -8549
rect 2126 -8605 2150 -8549
rect 2206 -8605 2250 -8549
rect 1950 -8649 2250 -8605
rect 1950 -8705 1990 -8649
rect 2046 -8705 2070 -8649
rect 2126 -8705 2150 -8649
rect 2206 -8705 2250 -8649
rect -3254 -8955 -3214 -8899
rect -3158 -8955 -3134 -8899
rect -3078 -8955 -3054 -8899
rect -2998 -8955 -2954 -8899
rect -3254 -8999 -2954 -8955
rect -3254 -9055 -3214 -8999
rect -3158 -9055 -3134 -8999
rect -3078 -9055 -3054 -8999
rect -2998 -9055 -2954 -8999
rect -3254 -9099 -2954 -9055
rect -3254 -9155 -3214 -9099
rect -3158 -9155 -3134 -9099
rect -3078 -9155 -3054 -9099
rect -2998 -9155 -2954 -9099
rect -3254 -9199 -2954 -9155
rect -3254 -9255 -3214 -9199
rect -3158 -9255 -3134 -9199
rect -3078 -9255 -3054 -9199
rect -2998 -9255 -2954 -9199
rect -3254 -9277 -2954 -9255
rect -508 -8899 -208 -8870
rect -508 -8955 -468 -8899
rect -412 -8955 -388 -8899
rect -332 -8955 -308 -8899
rect -252 -8955 -208 -8899
rect -508 -8999 -208 -8955
rect -508 -9055 -468 -8999
rect -412 -9055 -388 -8999
rect -332 -9055 -308 -8999
rect -252 -9055 -208 -8999
rect -508 -9099 -208 -9055
rect -508 -9155 -468 -9099
rect -412 -9155 -388 -9099
rect -332 -9155 -308 -9099
rect -252 -9155 -208 -9099
rect -508 -9199 -208 -9155
rect -508 -9255 -468 -9199
rect -412 -9255 -388 -9199
rect -332 -9255 -308 -9199
rect -252 -9255 -208 -9199
rect -2278 -9908 -1978 -9886
rect -2278 -9964 -2238 -9908
rect -2182 -9964 -2158 -9908
rect -2102 -9964 -2078 -9908
rect -2022 -9964 -1978 -9908
rect -2278 -10008 -1978 -9964
rect -2278 -10064 -2238 -10008
rect -2182 -10064 -2158 -10008
rect -2102 -10064 -2078 -10008
rect -2022 -10064 -1978 -10008
rect -2278 -10108 -1978 -10064
rect -2278 -10164 -2238 -10108
rect -2182 -10164 -2158 -10108
rect -2102 -10164 -2078 -10108
rect -2022 -10164 -1978 -10108
rect -2278 -10208 -1978 -10164
rect -2278 -10264 -2238 -10208
rect -2182 -10264 -2158 -10208
rect -2102 -10264 -2078 -10208
rect -2022 -10264 -1978 -10208
rect -7653 -10682 -7609 -10626
rect -7553 -10682 -7529 -10626
rect -7473 -10682 -7449 -10626
rect -7393 -10682 -7353 -10626
rect -7653 -10726 -7353 -10682
rect -7653 -10782 -7609 -10726
rect -7553 -10782 -7529 -10726
rect -7473 -10782 -7449 -10726
rect -7393 -10782 -7353 -10726
rect -7653 -10826 -7353 -10782
rect -7653 -10882 -7609 -10826
rect -7553 -10882 -7529 -10826
rect -7473 -10882 -7449 -10826
rect -7393 -10882 -7353 -10826
rect -7653 -10926 -7353 -10882
rect -7653 -10982 -7609 -10926
rect -7553 -10982 -7529 -10926
rect -7473 -10982 -7449 -10926
rect -7393 -10982 -7353 -10926
rect -7653 -11004 -7353 -10982
rect -3198 -10626 -2898 -10604
rect -3198 -10682 -3158 -10626
rect -3102 -10682 -3078 -10626
rect -3022 -10682 -2998 -10626
rect -2942 -10682 -2898 -10626
rect -3198 -10726 -2898 -10682
rect -3198 -10782 -3158 -10726
rect -3102 -10782 -3078 -10726
rect -3022 -10782 -2998 -10726
rect -2942 -10782 -2898 -10726
rect -3198 -10826 -2898 -10782
rect -3198 -10882 -3158 -10826
rect -3102 -10882 -3078 -10826
rect -3022 -10882 -2998 -10826
rect -2942 -10882 -2898 -10826
rect -3198 -10926 -2898 -10882
rect -3198 -10982 -3158 -10926
rect -3102 -10982 -3078 -10926
rect -3022 -10982 -2998 -10926
rect -2942 -10982 -2898 -10926
rect -3198 -13365 -2898 -10982
rect -3198 -13421 -3158 -13365
rect -3102 -13421 -3078 -13365
rect -3022 -13421 -2998 -13365
rect -2942 -13421 -2898 -13365
rect -3198 -13465 -2898 -13421
rect -3198 -13521 -3158 -13465
rect -3102 -13521 -3078 -13465
rect -3022 -13521 -2998 -13465
rect -2942 -13521 -2898 -13465
rect -3198 -13565 -2898 -13521
rect -3198 -13621 -3158 -13565
rect -3102 -13621 -3078 -13565
rect -3022 -13621 -2998 -13565
rect -2942 -13621 -2898 -13565
rect -3198 -13665 -2898 -13621
rect -3198 -13721 -3158 -13665
rect -3102 -13721 -3078 -13665
rect -3022 -13721 -2998 -13665
rect -2942 -13721 -2898 -13665
rect -3198 -13743 -2898 -13721
rect -2278 -14025 -1978 -10264
rect -1730 -10693 -1430 -10671
rect -1730 -10749 -1690 -10693
rect -1634 -10749 -1610 -10693
rect -1554 -10749 -1530 -10693
rect -1474 -10749 -1430 -10693
rect -1730 -11010 -1430 -10749
rect -1730 -11066 -1690 -11010
rect -1634 -11066 -1610 -11010
rect -1554 -11066 -1530 -11010
rect -1474 -11066 -1430 -11010
rect -1730 -12090 -1430 -11066
rect -1730 -12146 -1690 -12090
rect -1634 -12146 -1610 -12090
rect -1554 -12146 -1530 -12090
rect -1474 -12146 -1430 -12090
rect -1730 -12408 -1430 -12146
rect -1730 -12464 -1690 -12408
rect -1634 -12464 -1610 -12408
rect -1554 -12464 -1530 -12408
rect -1474 -12464 -1430 -12408
rect -1730 -12486 -1430 -12464
rect -2278 -14081 -2238 -14025
rect -2182 -14081 -2158 -14025
rect -2102 -14081 -2078 -14025
rect -2022 -14081 -1978 -14025
rect -2278 -14125 -1978 -14081
rect -2278 -14181 -2238 -14125
rect -2182 -14181 -2158 -14125
rect -2102 -14181 -2078 -14125
rect -2022 -14181 -1978 -14125
rect -2278 -14225 -1978 -14181
rect -2278 -14281 -2238 -14225
rect -2182 -14281 -2158 -14225
rect -2102 -14281 -2078 -14225
rect -2022 -14281 -1978 -14225
rect -2278 -14325 -1978 -14281
rect -2278 -14381 -2238 -14325
rect -2182 -14381 -2158 -14325
rect -2102 -14381 -2078 -14325
rect -2022 -14381 -1978 -14325
rect -3497 -15328 -3196 -15306
rect -3497 -15384 -3457 -15328
rect -3401 -15384 -3377 -15328
rect -3321 -15384 -3297 -15328
rect -3241 -15384 -3196 -15328
rect -3497 -15645 -3196 -15384
rect -3497 -15701 -3457 -15645
rect -3401 -15701 -3377 -15645
rect -3321 -15701 -3297 -15645
rect -3241 -15701 -3196 -15645
rect -3497 -16725 -3196 -15701
rect -3497 -16781 -3457 -16725
rect -3401 -16781 -3377 -16725
rect -3321 -16781 -3297 -16725
rect -3241 -16781 -3196 -16725
rect -2278 -16727 -1978 -14381
rect -941 -14025 -641 -11259
rect -508 -11593 -208 -9255
rect 1950 -10852 2250 -8705
rect 4312 -8899 4612 -6102
rect 5753 -6238 6053 -4956
rect 5753 -6294 5793 -6238
rect 5849 -6294 5873 -6238
rect 5929 -6294 5953 -6238
rect 6009 -6294 6053 -6238
rect 5753 -6558 6053 -6294
rect 5753 -6614 5793 -6558
rect 5849 -6614 5873 -6558
rect 5929 -6614 5953 -6558
rect 6009 -6614 6053 -6558
rect 5753 -6636 6053 -6614
rect 4312 -8955 4352 -8899
rect 4408 -8955 4432 -8899
rect 4488 -8955 4512 -8899
rect 4568 -8955 4612 -8899
rect 4312 -8999 4612 -8955
rect 4312 -9055 4352 -8999
rect 4408 -9055 4432 -8999
rect 4488 -9055 4512 -8999
rect 4568 -9055 4612 -8999
rect 4312 -9099 4612 -9055
rect 4312 -9155 4352 -9099
rect 4408 -9155 4432 -9099
rect 4488 -9155 4512 -9099
rect 4568 -9155 4612 -9099
rect 4312 -9199 4612 -9155
rect 4312 -9255 4352 -9199
rect 4408 -9255 4432 -9199
rect 4488 -9255 4512 -9199
rect 4568 -9255 4612 -9199
rect 4312 -9277 4612 -9255
rect 6889 -10039 7189 975
rect 8267 151 8567 3756
rect 9816 3558 10116 4478
rect 10784 9429 11084 10189
rect 10784 9373 10828 9429
rect 10884 9373 10908 9429
rect 10964 9373 10988 9429
rect 11044 9373 11084 9429
rect 10784 7909 11084 9373
rect 10784 7853 10828 7909
rect 10884 7853 10908 7909
rect 10964 7853 10988 7909
rect 11044 7853 11084 7909
rect 10784 6215 11084 7853
rect 10784 6159 10828 6215
rect 10884 6159 10908 6215
rect 10964 6159 10988 6215
rect 11044 6159 11084 6215
rect 10784 4695 11084 6159
rect 10784 4639 10828 4695
rect 10884 4639 10908 4695
rect 10964 4639 10988 4695
rect 11044 4639 11084 4695
rect 10784 3878 11084 4639
rect 14162 9429 14462 10189
rect 14162 9373 14206 9429
rect 14262 9373 14286 9429
rect 14342 9373 14366 9429
rect 14422 9373 14462 9429
rect 14162 7909 14462 9373
rect 14162 7853 14206 7909
rect 14262 7853 14286 7909
rect 14342 7853 14366 7909
rect 14422 7853 14462 7909
rect 14162 6215 14462 7853
rect 14162 6159 14206 6215
rect 14262 6159 14286 6215
rect 14342 6159 14366 6215
rect 14422 6159 14462 6215
rect 14162 4695 14462 6159
rect 14162 4639 14206 4695
rect 14262 4639 14286 4695
rect 14342 4639 14366 4695
rect 14422 4639 14462 4695
rect 14162 3878 14462 4639
rect 15130 9590 15430 10510
rect 15130 9534 15170 9590
rect 15226 9534 15250 9590
rect 15306 9534 15330 9590
rect 15386 9534 15430 9590
rect 15130 8077 15430 9534
rect 15130 8021 15170 8077
rect 15226 8021 15250 8077
rect 15306 8021 15330 8077
rect 15386 8021 15430 8077
rect 15130 6046 15430 8021
rect 15130 5990 15170 6046
rect 15226 5990 15250 6046
rect 15306 5990 15330 6046
rect 15386 5990 15430 6046
rect 15130 4534 15430 5990
rect 15130 4478 15170 4534
rect 15226 4478 15250 4534
rect 15306 4478 15330 4534
rect 15386 4478 15430 4534
rect 9816 -604 10116 316
rect 9816 -660 9856 -604
rect 9912 -660 9936 -604
rect 9992 -660 10016 -604
rect 10072 -660 10116 -604
rect 9816 -2117 10116 -660
rect 9816 -2173 9856 -2117
rect 9912 -2173 9936 -2117
rect 9992 -2173 10016 -2117
rect 10072 -2173 10116 -2117
rect 9816 -4148 10116 -2173
rect 9816 -4204 9856 -4148
rect 9912 -4204 9936 -4148
rect 9992 -4204 10016 -4148
rect 10072 -4204 10116 -4148
rect 9816 -5660 10116 -4204
rect 9816 -5716 9856 -5660
rect 9912 -5716 9936 -5660
rect 9992 -5716 10016 -5660
rect 10072 -5716 10116 -5660
rect 9816 -6636 10116 -5716
rect 10784 -765 11084 -5
rect 12332 -182 12914 3760
rect 15130 3558 15430 4478
rect 18395 10488 18695 10510
rect 18395 10432 18435 10488
rect 18491 10432 18515 10488
rect 18571 10432 18595 10488
rect 18651 10432 18695 10488
rect 18395 10167 18695 10432
rect 18395 10111 18435 10167
rect 18491 10111 18515 10167
rect 18571 10111 18595 10167
rect 18651 10111 18695 10167
rect 18395 8841 18695 10111
rect 18395 8785 18435 8841
rect 18491 8785 18515 8841
rect 18571 8785 18595 8841
rect 18651 8785 18695 8841
rect 18395 8509 18695 8785
rect 18395 8453 18435 8509
rect 18491 8453 18515 8509
rect 18571 8453 18595 8509
rect 18651 8453 18695 8509
rect 18395 5614 18695 8453
rect 18395 5558 18435 5614
rect 18491 5558 18515 5614
rect 18571 5558 18595 5614
rect 18651 5558 18695 5614
rect 18395 5288 18695 5558
rect 18395 5232 18435 5288
rect 18491 5232 18515 5288
rect 18571 5232 18595 5288
rect 18651 5232 18695 5288
rect 18395 3956 18695 5232
rect 18395 3900 18435 3956
rect 18491 3900 18515 3956
rect 18571 3900 18595 3956
rect 18651 3900 18695 3956
rect 10784 -821 10828 -765
rect 10884 -821 10908 -765
rect 10964 -821 10988 -765
rect 11044 -821 11084 -765
rect 10784 -2285 11084 -821
rect 10784 -2341 10828 -2285
rect 10884 -2341 10908 -2285
rect 10964 -2341 10988 -2285
rect 11044 -2341 11084 -2285
rect 10784 -3979 11084 -2341
rect 10784 -4035 10828 -3979
rect 10884 -4035 10908 -3979
rect 10964 -4035 10988 -3979
rect 11044 -4035 11084 -3979
rect 10784 -5499 11084 -4035
rect 14162 -765 14462 -5
rect 14162 -821 14206 -765
rect 14262 -821 14286 -765
rect 14342 -821 14366 -765
rect 14422 -821 14462 -765
rect 14162 -2285 14462 -821
rect 14162 -2341 14206 -2285
rect 14262 -2341 14286 -2285
rect 14342 -2341 14366 -2285
rect 14422 -2341 14462 -2285
rect 14162 -3979 14462 -2341
rect 14162 -4035 14206 -3979
rect 14262 -4035 14286 -3979
rect 14342 -4035 14366 -3979
rect 14422 -4035 14462 -3979
rect 10784 -5555 10828 -5499
rect 10884 -5555 10908 -5499
rect 10964 -5555 10988 -5499
rect 11044 -5555 11084 -5499
rect 10784 -6316 11084 -5555
rect 6889 -10095 6929 -10039
rect 6985 -10095 7009 -10039
rect 7065 -10095 7089 -10039
rect 7145 -10095 7189 -10039
rect 6889 -10139 7189 -10095
rect 6889 -10195 6929 -10139
rect 6985 -10195 7009 -10139
rect 7065 -10195 7089 -10139
rect 7145 -10195 7189 -10139
rect 6889 -10239 7189 -10195
rect 6889 -10295 6929 -10239
rect 6985 -10295 7009 -10239
rect 7065 -10295 7089 -10239
rect 7145 -10295 7189 -10239
rect 6889 -10339 7189 -10295
rect 6889 -10395 6929 -10339
rect 6985 -10395 7009 -10339
rect 7065 -10395 7089 -10339
rect 7145 -10395 7189 -10339
rect 6889 -10439 7189 -10395
rect 6889 -10495 6933 -10439
rect 6989 -10495 7013 -10439
rect 7069 -10495 7093 -10439
rect 7149 -10495 7189 -10439
rect 6889 -10517 7189 -10495
rect 3160 -10693 3460 -10671
rect 3160 -10749 3204 -10693
rect 3260 -10749 3284 -10693
rect 3340 -10749 3364 -10693
rect 3420 -10749 3460 -10693
rect -941 -14081 -901 -14025
rect -845 -14081 -821 -14025
rect -765 -14081 -741 -14025
rect -685 -14081 -641 -14025
rect -941 -14125 -641 -14081
rect -941 -14181 -901 -14125
rect -845 -14181 -821 -14125
rect -765 -14181 -741 -14125
rect -685 -14181 -641 -14125
rect -941 -14225 -641 -14181
rect -941 -14281 -901 -14225
rect -845 -14281 -821 -14225
rect -765 -14281 -741 -14225
rect -685 -14281 -641 -14225
rect -941 -14325 -641 -14281
rect -941 -14381 -901 -14325
rect -845 -14381 -821 -14325
rect -765 -14381 -741 -14325
rect -685 -14381 -641 -14325
rect -941 -14403 -641 -14381
rect 180 -13359 480 -13343
rect 180 -13365 481 -13359
rect 180 -13421 220 -13365
rect 276 -13421 300 -13365
rect 356 -13421 380 -13365
rect 436 -13421 481 -13365
rect 180 -13465 481 -13421
rect 180 -13521 220 -13465
rect 276 -13521 300 -13465
rect 356 -13521 380 -13465
rect 436 -13521 481 -13465
rect 180 -13565 481 -13521
rect 180 -13621 220 -13565
rect 276 -13621 300 -13565
rect 356 -13621 380 -13565
rect 436 -13621 481 -13565
rect 180 -13665 481 -13621
rect 180 -13721 220 -13665
rect 276 -13721 300 -13665
rect 356 -13721 380 -13665
rect 436 -13721 481 -13665
rect 180 -15883 481 -13721
rect 1261 -13365 1561 -13343
rect 1261 -13421 1301 -13365
rect 1357 -13421 1381 -13365
rect 1437 -13421 1461 -13365
rect 1517 -13421 1561 -13365
rect 1261 -13465 1561 -13421
rect 1261 -13521 1301 -13465
rect 1357 -13521 1381 -13465
rect 1437 -13521 1461 -13465
rect 1517 -13521 1561 -13465
rect 1261 -13565 1561 -13521
rect 1261 -13621 1301 -13565
rect 1357 -13621 1381 -13565
rect 1437 -13621 1461 -13565
rect 1517 -13621 1561 -13565
rect 1261 -13665 1561 -13621
rect 1261 -13721 1301 -13665
rect 1357 -13721 1381 -13665
rect 1437 -13721 1461 -13665
rect 1517 -13721 1561 -13665
rect 1261 -15883 1561 -13721
rect 2382 -13365 2682 -10798
rect 3160 -11010 3460 -10749
rect 7965 -10693 8265 -8327
rect 8690 -9528 8990 -6715
rect 11898 -7758 12198 -4879
rect 11756 -7780 12198 -7758
rect 11756 -7836 11796 -7780
rect 11852 -7836 11876 -7780
rect 11932 -7836 11956 -7780
rect 12012 -7836 12198 -7780
rect 11756 -7880 12198 -7836
rect 11756 -7936 11796 -7880
rect 11852 -7936 11876 -7880
rect 11932 -7936 11956 -7880
rect 12012 -7936 12198 -7880
rect 11756 -7974 12198 -7936
rect 8690 -9584 8730 -9528
rect 8786 -9584 8810 -9528
rect 8866 -9584 8890 -9528
rect 8946 -9584 8990 -9528
rect 8690 -9628 8990 -9584
rect 8690 -9684 8730 -9628
rect 8786 -9684 8810 -9628
rect 8866 -9684 8890 -9628
rect 8946 -9684 8990 -9628
rect 8690 -9728 8990 -9684
rect 8690 -9784 8730 -9728
rect 8786 -9784 8810 -9728
rect 8866 -9784 8890 -9728
rect 8946 -9784 8990 -9728
rect 8690 -9828 8990 -9784
rect 8690 -9884 8730 -9828
rect 8786 -9884 8810 -9828
rect 8866 -9884 8890 -9828
rect 8946 -9884 8990 -9828
rect 8690 -9906 8990 -9884
rect 11645 -7980 12198 -7974
rect 11645 -8036 11796 -7980
rect 11852 -8036 11876 -7980
rect 11932 -8036 11956 -7980
rect 12012 -8036 12198 -7980
rect 11645 -8080 12198 -8036
rect 11645 -8136 11796 -8080
rect 11852 -8136 11876 -8080
rect 11932 -8136 11956 -8080
rect 12012 -8136 12198 -8080
rect 11645 -8158 12198 -8136
rect 13048 -7780 13348 -4879
rect 14162 -5499 14462 -4035
rect 14162 -5555 14206 -5499
rect 14262 -5555 14286 -5499
rect 14342 -5555 14366 -5499
rect 14422 -5555 14462 -5499
rect 14162 -6316 14462 -5555
rect 15130 -604 15430 316
rect 16679 151 16979 3756
rect 18395 3636 18695 3900
rect 18395 3580 18435 3636
rect 18491 3580 18515 3636
rect 18571 3580 18595 3636
rect 18651 3580 18695 3636
rect 15130 -660 15170 -604
rect 15226 -660 15250 -604
rect 15306 -660 15330 -604
rect 15386 -660 15430 -604
rect 15130 -2117 15430 -660
rect 15130 -2173 15170 -2117
rect 15226 -2173 15250 -2117
rect 15306 -2173 15330 -2117
rect 15386 -2173 15430 -2117
rect 15130 -4148 15430 -2173
rect 15130 -4204 15170 -4148
rect 15226 -4204 15250 -4148
rect 15306 -4204 15330 -4148
rect 15386 -4204 15430 -4148
rect 15130 -5660 15430 -4204
rect 15130 -5716 15170 -5660
rect 15226 -5716 15250 -5660
rect 15306 -5716 15330 -5660
rect 15386 -5716 15430 -5660
rect 15130 -6636 15430 -5716
rect 13048 -7836 13088 -7780
rect 13144 -7836 13168 -7780
rect 13224 -7836 13248 -7780
rect 13304 -7836 13348 -7780
rect 13048 -7880 13348 -7836
rect 13048 -7936 13088 -7880
rect 13144 -7936 13168 -7880
rect 13224 -7936 13248 -7880
rect 13304 -7936 13348 -7880
rect 13048 -7980 13348 -7936
rect 13048 -8036 13088 -7980
rect 13144 -8036 13168 -7980
rect 13224 -8036 13248 -7980
rect 13304 -8036 13348 -7980
rect 13048 -8080 13348 -8036
rect 13048 -8136 13088 -8080
rect 13144 -8136 13168 -8080
rect 13224 -8136 13248 -8080
rect 13304 -8136 13348 -8080
rect 13048 -8158 13348 -8136
rect 11645 -10498 11945 -8158
rect 13593 -9528 13894 -9496
rect 13593 -9584 13633 -9528
rect 13689 -9584 13713 -9528
rect 13769 -9584 13793 -9528
rect 13849 -9584 13894 -9528
rect 13593 -9628 13894 -9584
rect 13593 -9684 13633 -9628
rect 13689 -9684 13713 -9628
rect 13769 -9684 13793 -9628
rect 13849 -9684 13894 -9628
rect 13593 -9728 13894 -9684
rect 13593 -9784 13633 -9728
rect 13689 -9784 13713 -9728
rect 13769 -9784 13793 -9728
rect 13849 -9784 13894 -9728
rect 13593 -9828 13894 -9784
rect 13593 -9884 13633 -9828
rect 13689 -9884 13713 -9828
rect 13769 -9884 13793 -9828
rect 13849 -9884 13894 -9828
rect 7965 -10749 8005 -10693
rect 8061 -10749 8085 -10693
rect 8141 -10749 8165 -10693
rect 8221 -10749 8265 -10693
rect 3160 -11066 3204 -11010
rect 3260 -11066 3284 -11010
rect 3340 -11066 3364 -11010
rect 3420 -11066 3460 -11010
rect 3160 -12090 3460 -11066
rect 3160 -12146 3204 -12090
rect 3260 -12146 3284 -12090
rect 3340 -12146 3364 -12090
rect 3420 -12146 3460 -12090
rect 3160 -12408 3460 -12146
rect 7477 -11010 7777 -10988
rect 7477 -11066 7517 -11010
rect 7573 -11066 7597 -11010
rect 7653 -11066 7677 -11010
rect 7733 -11066 7777 -11010
rect 7477 -12090 7777 -11066
rect 7477 -12146 7517 -12090
rect 7573 -12146 7597 -12090
rect 7653 -12146 7677 -12090
rect 7733 -12146 7777 -12090
rect 7477 -12168 7777 -12146
rect 3160 -12464 3204 -12408
rect 3260 -12464 3284 -12408
rect 3340 -12464 3364 -12408
rect 3420 -12464 3460 -12408
rect 3160 -12486 3460 -12464
rect 7965 -12408 8265 -10749
rect 12632 -11011 12933 -10989
rect 12632 -11067 12672 -11011
rect 12728 -11067 12752 -11011
rect 12808 -11067 12832 -11011
rect 12888 -11067 12933 -11011
rect 12632 -12090 12933 -11067
rect 12632 -12146 12672 -12090
rect 12728 -12146 12752 -12090
rect 12808 -12146 12832 -12090
rect 12888 -12146 12933 -12090
rect 12632 -12168 12933 -12146
rect 7965 -12464 8005 -12408
rect 8061 -12464 8085 -12408
rect 8141 -12464 8165 -12408
rect 8221 -12464 8265 -12408
rect 7965 -12486 8265 -12464
rect 2382 -13421 2422 -13365
rect 2478 -13421 2502 -13365
rect 2558 -13421 2582 -13365
rect 2638 -13421 2682 -13365
rect 2382 -13465 2682 -13421
rect 2382 -13521 2422 -13465
rect 2478 -13521 2502 -13465
rect 2558 -13521 2582 -13465
rect 2638 -13521 2682 -13465
rect 2382 -13565 2682 -13521
rect 2382 -13621 2422 -13565
rect 2478 -13621 2502 -13565
rect 2558 -13621 2582 -13565
rect 2638 -13621 2682 -13565
rect 2382 -13665 2682 -13621
rect 2382 -13721 2422 -13665
rect 2478 -13721 2502 -13665
rect 2558 -13721 2582 -13665
rect 2638 -13721 2682 -13665
rect 2382 -13743 2682 -13721
rect 9622 -13484 9922 -13462
rect 9622 -13540 9662 -13484
rect 9718 -13540 9742 -13484
rect 9798 -13540 9822 -13484
rect 9878 -13540 9922 -13484
rect 9622 -13584 9922 -13540
rect 9622 -13640 9662 -13584
rect 9718 -13640 9742 -13584
rect 9798 -13640 9822 -13584
rect 9878 -13640 9922 -13584
rect 9622 -13684 9922 -13640
rect 9622 -13740 9662 -13684
rect 9718 -13740 9742 -13684
rect 9798 -13740 9822 -13684
rect 9878 -13740 9922 -13684
rect 9622 -13784 9922 -13740
rect 9622 -13840 9662 -13784
rect 9718 -13840 9742 -13784
rect 9798 -13840 9822 -13784
rect 9878 -13840 9922 -13784
rect 3719 -14025 4019 -14003
rect 3719 -14081 3759 -14025
rect 3815 -14081 3839 -14025
rect 3895 -14081 3919 -14025
rect 3975 -14081 4019 -14025
rect 3719 -14125 4019 -14081
rect 3719 -14181 3759 -14125
rect 3815 -14181 3839 -14125
rect 3895 -14181 3919 -14125
rect 3975 -14181 4019 -14125
rect 3719 -14225 4019 -14181
rect 3719 -14281 3759 -14225
rect 3815 -14281 3839 -14225
rect 3895 -14281 3919 -14225
rect 3975 -14281 4019 -14225
rect 3719 -14325 4019 -14281
rect 3719 -14381 3759 -14325
rect 3815 -14381 3839 -14325
rect 3895 -14381 3919 -14325
rect 3975 -14381 4019 -14325
rect 3719 -16727 4019 -14381
rect 4894 -15328 5194 -15306
rect 4894 -15384 4938 -15328
rect 4994 -15384 5018 -15328
rect 5074 -15384 5098 -15328
rect 5154 -15384 5194 -15328
rect 4894 -15645 5194 -15384
rect 4894 -15701 4938 -15645
rect 4994 -15701 5018 -15645
rect 5074 -15701 5098 -15645
rect 5154 -15701 5194 -15645
rect 4894 -16725 5194 -15701
rect -3497 -17042 -3196 -16781
rect -3497 -17098 -3457 -17042
rect -3401 -17098 -3377 -17042
rect -3321 -17098 -3297 -17042
rect -3241 -17098 -3196 -17042
rect -3497 -17120 -3196 -17098
rect 4894 -16781 4938 -16725
rect 4994 -16781 5018 -16725
rect 5074 -16781 5098 -16725
rect 5154 -16781 5194 -16725
rect 4894 -17042 5194 -16781
rect 4894 -17098 4938 -17042
rect 4994 -17098 5018 -17042
rect 5074 -17098 5098 -17042
rect 5154 -17098 5194 -17042
rect 4894 -17120 5194 -17098
rect 8404 -15328 8704 -15306
rect 8404 -15384 8444 -15328
rect 8500 -15384 8524 -15328
rect 8580 -15384 8604 -15328
rect 8660 -15384 8704 -15328
rect 8404 -15645 8704 -15384
rect 8404 -15701 8444 -15645
rect 8500 -15701 8524 -15645
rect 8580 -15701 8604 -15645
rect 8660 -15701 8704 -15645
rect 8404 -16725 8704 -15701
rect 9622 -16186 9922 -13840
rect 12081 -14040 12381 -12910
rect 13161 -13484 13461 -11338
rect 13593 -12021 13894 -9884
rect 16256 -9528 16556 -6715
rect 16679 -7399 16979 -7299
rect 16256 -9584 16296 -9528
rect 16352 -9584 16376 -9528
rect 16432 -9584 16456 -9528
rect 16512 -9584 16556 -9528
rect 16256 -9628 16556 -9584
rect 16256 -9684 16296 -9628
rect 16352 -9684 16376 -9628
rect 16432 -9684 16456 -9628
rect 16512 -9684 16556 -9628
rect 16256 -9728 16556 -9684
rect 16256 -9784 16296 -9728
rect 16352 -9784 16376 -9728
rect 16432 -9784 16456 -9728
rect 16512 -9784 16556 -9728
rect 16256 -9828 16556 -9784
rect 16256 -9884 16296 -9828
rect 16352 -9884 16376 -9828
rect 16432 -9884 16456 -9828
rect 16512 -9884 16556 -9828
rect 16256 -9906 16556 -9884
rect 17320 -8899 17620 -8644
rect 17320 -8955 17360 -8899
rect 17416 -8955 17440 -8899
rect 17496 -8955 17520 -8899
rect 17576 -8955 17620 -8899
rect 17320 -8999 17620 -8955
rect 17320 -9055 17360 -8999
rect 17416 -9055 17440 -8999
rect 17496 -9055 17520 -8999
rect 17576 -9055 17620 -8999
rect 17320 -9099 17620 -9055
rect 17320 -9155 17360 -9099
rect 17416 -9155 17440 -9099
rect 17496 -9155 17520 -9099
rect 17576 -9155 17620 -9099
rect 17320 -9199 17620 -9155
rect 17320 -9255 17360 -9199
rect 17416 -9255 17440 -9199
rect 17496 -9255 17520 -9199
rect 17576 -9255 17620 -9199
rect 17320 -10693 17620 -9255
rect 18395 -10039 18695 3580
rect 18395 -10095 18439 -10039
rect 18495 -10095 18519 -10039
rect 18575 -10095 18599 -10039
rect 18655 -10095 18695 -10039
rect 18395 -10139 18695 -10095
rect 18395 -10195 18439 -10139
rect 18495 -10195 18519 -10139
rect 18575 -10195 18599 -10139
rect 18655 -10195 18695 -10139
rect 18395 -10239 18695 -10195
rect 18395 -10295 18439 -10239
rect 18495 -10295 18519 -10239
rect 18575 -10295 18599 -10239
rect 18655 -10295 18695 -10239
rect 18395 -10339 18695 -10295
rect 18395 -10395 18439 -10339
rect 18495 -10395 18519 -10339
rect 18575 -10395 18599 -10339
rect 18655 -10395 18695 -10339
rect 18395 -10439 18695 -10395
rect 18395 -10495 18435 -10439
rect 18491 -10495 18515 -10439
rect 18571 -10495 18595 -10439
rect 18651 -10495 18695 -10439
rect 18395 -10517 18695 -10495
rect 17320 -10749 17364 -10693
rect 17420 -10749 17444 -10693
rect 17500 -10749 17524 -10693
rect 17580 -10749 17620 -10693
rect 17320 -12408 17620 -10749
rect 17807 -10989 18107 -10988
rect 17807 -11010 18108 -10989
rect 17807 -11066 17851 -11010
rect 17907 -11066 17931 -11010
rect 17987 -11066 18011 -11010
rect 18067 -11066 18108 -11010
rect 17807 -12090 18108 -11066
rect 17807 -12146 17851 -12090
rect 17907 -12146 17931 -12090
rect 17987 -12146 18011 -12090
rect 18067 -12146 18108 -12090
rect 17807 -12168 18108 -12146
rect 17320 -12464 17364 -12408
rect 17420 -12464 17444 -12408
rect 17500 -12464 17524 -12408
rect 17580 -12464 17620 -12408
rect 17320 -12486 17620 -12464
rect 13161 -13540 13201 -13484
rect 13257 -13540 13281 -13484
rect 13337 -13540 13361 -13484
rect 13417 -13540 13461 -13484
rect 13161 -13584 13461 -13540
rect 13161 -13640 13201 -13584
rect 13257 -13640 13281 -13584
rect 13337 -13640 13361 -13584
rect 13417 -13640 13461 -13584
rect 13161 -13684 13461 -13640
rect 13161 -13740 13201 -13684
rect 13257 -13740 13281 -13684
rect 13337 -13740 13361 -13684
rect 13417 -13740 13461 -13684
rect 13161 -13784 13461 -13740
rect 13161 -13840 13201 -13784
rect 13257 -13840 13281 -13784
rect 13337 -13840 13361 -13784
rect 13417 -13840 13461 -13784
rect 13161 -13862 13461 -13840
rect 15620 -13484 15920 -13462
rect 15620 -13540 15660 -13484
rect 15716 -13540 15740 -13484
rect 15796 -13540 15820 -13484
rect 15876 -13540 15920 -13484
rect 15620 -13584 15920 -13540
rect 15620 -13640 15660 -13584
rect 15716 -13640 15740 -13584
rect 15796 -13640 15820 -13584
rect 15876 -13640 15920 -13584
rect 15620 -13684 15920 -13640
rect 15620 -13740 15660 -13684
rect 15716 -13740 15740 -13684
rect 15796 -13740 15820 -13684
rect 15876 -13740 15920 -13684
rect 15620 -13784 15920 -13740
rect 15620 -13840 15660 -13784
rect 15716 -13840 15740 -13784
rect 15796 -13840 15820 -13784
rect 15876 -13840 15920 -13784
rect 12081 -14096 12121 -14040
rect 12177 -14096 12201 -14040
rect 12257 -14096 12281 -14040
rect 12337 -14096 12381 -14040
rect 12081 -14140 12381 -14096
rect 12081 -14196 12121 -14140
rect 12177 -14196 12201 -14140
rect 12257 -14196 12281 -14140
rect 12337 -14196 12381 -14140
rect 12081 -14240 12381 -14196
rect 12081 -14296 12121 -14240
rect 12177 -14296 12201 -14240
rect 12257 -14296 12281 -14240
rect 12337 -14296 12381 -14240
rect 12081 -14340 12381 -14296
rect 12081 -14396 12121 -14340
rect 12177 -14396 12201 -14340
rect 12257 -14396 12281 -14340
rect 12337 -14396 12381 -14340
rect 12081 -15435 12381 -14396
rect 13161 -14040 13461 -14018
rect 13161 -14096 13201 -14040
rect 13257 -14096 13281 -14040
rect 13337 -14096 13361 -14040
rect 13417 -14096 13461 -14040
rect 13161 -14140 13461 -14096
rect 13161 -14196 13201 -14140
rect 13257 -14196 13281 -14140
rect 13337 -14196 13361 -14140
rect 13417 -14196 13461 -14140
rect 13161 -14240 13461 -14196
rect 13161 -14296 13201 -14240
rect 13257 -14296 13281 -14240
rect 13337 -14296 13361 -14240
rect 13417 -14296 13461 -14240
rect 13161 -14340 13461 -14296
rect 13161 -14396 13201 -14340
rect 13257 -14396 13281 -14340
rect 13337 -14396 13361 -14340
rect 13417 -14396 13461 -14340
rect 13161 -16543 13461 -14396
rect 15620 -16186 15920 -13840
rect 16794 -15328 17094 -15306
rect 16794 -15384 16838 -15328
rect 16894 -15384 16918 -15328
rect 16974 -15384 16998 -15328
rect 17054 -15384 17094 -15328
rect 16794 -15645 17094 -15384
rect 16794 -15701 16838 -15645
rect 16894 -15701 16918 -15645
rect 16974 -15701 16998 -15645
rect 17054 -15701 17094 -15645
rect 8404 -16781 8444 -16725
rect 8500 -16781 8524 -16725
rect 8580 -16781 8604 -16725
rect 8660 -16781 8704 -16725
rect 8404 -17042 8704 -16781
rect 8404 -17098 8444 -17042
rect 8500 -17098 8524 -17042
rect 8580 -17098 8604 -17042
rect 8660 -17098 8704 -17042
rect 8404 -17120 8704 -17098
rect 16794 -16725 17094 -15701
rect 16794 -16781 16838 -16725
rect 16894 -16781 16918 -16725
rect 16974 -16781 16998 -16725
rect 17054 -16781 17094 -16725
rect 16794 -17042 17094 -16781
rect 16794 -17098 16838 -17042
rect 16894 -17098 16918 -17042
rect 16974 -17098 16998 -17042
rect 17054 -17098 17094 -17042
rect 16794 -17120 17094 -17098
use nfets_2x  nfets_2x_0
timestamp 1698888477
transform -1 0 16515 0 1 -10535
box -270 -3101 3355 1015
use nfets_2x  nfets_2x_1
timestamp 1698888477
transform 1 0 9027 0 1 -10535
box -270 -3101 3355 1015
use nfets_2x  nfets_2x_2
timestamp 1698888477
transform 1 0 -672 0 1 -10535
box -270 -3101 3355 1015
use nfets_4x  nfets_4x_0
timestamp 1698888477
transform 1 0 9459 0 1 -15170
box -270 -3101 6894 1015
use nfets_4x  nfets_4x_1
timestamp 1698888477
transform 1 0 -2441 0 1 -15170
box -270 -3101 6894 1015
use pfets_4x  pfets_4x_0
timestamp 1698888477
transform 1 0 7375 0 1 11122
box 816 -8987 9679 813
use pfets_4x  pfets_4x_1
timestamp 1698888477
transform 1 0 7375 0 1 928
box 816 -8987 9679 813
use pfets_4x  pfets_4x_2
timestamp 1698888477
transform 1 0 -4568 0 1 928
box 816 -8987 9679 813
use pfets_4x  pfets_4x_3
timestamp 1698888477
transform 1 0 -16534 0 1 928
box 816 -8987 9679 813
use pfets_4x  pfets_4x_4
timestamp 1698888477
transform 1 0 -4568 0 1 11122
box 816 -8987 9679 813
use pfets_4x  pfets_4x_5
timestamp 1698888477
transform 1 0 -26246 0 1 928
box 816 -8987 9679 813
use pfets_8x  pfets_8x_0
timestamp 1698888477
transform 1 0 -25658 0 1 11416
box 800 -9284 18380 520
<< labels >>
flabel metal3 s -355 -9356 -355 -9356 2 FreeSans 150 0 0 0 VO2
flabel metal3 s 11676 -8070 11676 -8070 2 FreeSans 3126 0 0 0 VD1
flabel metal3 s 2172 -8788 2172 -8788 2 FreeSans 150 0 0 0 VO1
flabel metal3 s 12781 -11528 12781 -11528 2 FreeSans 150 0 0 0 VCM
flabel metal3 s 7558 -11576 7558 -11576 2 FreeSans 150 0 0 0 VCM
flabel metal3 s 8502 -16196 8502 -16196 2 FreeSans 150 0 0 0 VB2
flabel metal3 s 12160 -14286 12160 -14286 2 FreeSans 150 0 0 0 VIT_N1
flabel metal3 s 13258 -13777 13258 -13777 2 FreeSans 150 0 0 0 VIT_N2
flabel metal3 s 16327 -8187 16327 -8187 2 FreeSans 3126 0 0 0 VD2
flabel metal3 s -20453 -8943 -20453 -8943 2 FreeSans 150 0 0 0 SUM_P
flabel metal3 s -17229 -8269 -17229 -8269 2 FreeSans 150 0 0 0 SUM_N
flabel metal3 s -19962 1704 -19962 1704 2 FreeSans 3126 0 0 0 VIT_P1
flabel metal3 s -11346 2037 -11346 2037 2 FreeSans 150 0 0 0 VIT_P2
flabel metal3 s -21054 1685 -21054 1685 2 FreeSans 3126 0 0 0 VIT_P1
flabel metal3 s -21101 984 -21101 984 2 FreeSans 3126 0 0 0 VIT_P1
flabel metal3 s -10500 2335 -10500 2335 2 FreeSans 3126 0 0 0 VIT_P1
flabel metal3 s -4637 -3565 -4637 -3565 2 FreeSans 3126 0 0 0 VB4
flabel metal3 s -880 -14106 -880 -14106 2 FreeSans 150 0 0 0 SUM_N
flabel metal3 s 2441 -13789 2441 -13789 2 FreeSans 150 0 0 0 SUM_P
flabel metal3 s 2441 -13789 2441 -13789 2 FreeSans 150 0 0 0 SUM_P
flabel metal3 s 4419 1567 4419 1567 2 FreeSans 150 0 0 0 VD6
flabel metal3 s 630 2205 630 2205 2 FreeSans 150 0 0 0 VD5
flabel metal3 s 5867 7170 5867 7170 2 FreeSans 3126 0 0 0 VCMFB
flabel metal3 s -4577 7055 -4577 7055 2 FreeSans 3126 0 0 0 VCMFB
flabel metal3 s 17372 -12183 17579 -9106 2 FreeSans 150 0 0 0 VO2
port 1 nsew
flabel metal3 s 17475 -10644 17475 -10644 2 FreeSans 150 0 0 0 VO2
flabel metal3 s 8017 -11965 8227 -9117 2 FreeSans 150 0 0 0 VO1
port 2 nsew
flabel metal3 s 17848 -12024 18065 -11121 2 FreeSans 150 0 0 0 VCM
port 3 nsew
flabel metal3 s -26504 -4459 -26264 -1797 2 FreeSans 3126 0 0 0 VI_1B
port 4 nsew
flabel metal3 s -27002 -4415 -26769 -1772 2 FreeSans 3126 0 0 0 VI_1A
port 5 nsew
flabel metal3 s -6065 -4469 -5834 -1805 2 FreeSans 3126 0 0 0 VI_2B
port 6 nsew
flabel metal3 s -5574 -4505 -5323 -1831 2 FreeSans 3126 180 0 0 VI_2A
port 7 nsew
flabel metal3 s 5782 -4511 6030 -2371 2 FreeSans 3126 180 0 0 VB4
port 8 nsew
flabel metal3 s 3193 -12060 3423 -11132 2 FreeSans 3126 0 0 0 VB3
port 9 nsew
flabel metal3 s -3463 -16657 -3232 -15771 2 FreeSans 3126 0 0 0 VB2
port 10 nsew
flabel metal3 s -25746 5703 -25484 8346 2 FreeSans 3126 0 0 0 VB1
port 11 nsew
flabel metal1 s 4784 -17940 8713 -17256 2 FreeSans 3126 0 0 0 AVSS
port 12 nsew
flabel metal1 s -7050 4869 -4249 11281 2 FreeSans 3126 0 0 0 AVDD
port 13 nsew
<< end >>
