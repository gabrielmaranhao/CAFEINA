magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< nwell >>
rect 800 -9284 18380 520
<< pmoshvt >>
rect 1017 68 1217 268
rect 1469 68 1669 268
rect 1727 68 1927 268
rect 1985 68 2185 268
rect 2243 68 2443 268
rect 2695 68 2895 268
rect 2953 68 3153 268
rect 3211 68 3411 268
rect 3663 68 3863 268
rect 3921 68 4121 268
rect 4179 68 4379 268
rect 4437 68 4637 268
rect 4888 68 5088 268
rect 5374 68 5574 268
rect 5826 68 6026 268
rect 6084 68 6284 268
rect 6342 68 6542 268
rect 6600 68 6800 268
rect 7052 68 7252 268
rect 7310 68 7510 268
rect 7568 68 7768 268
rect 8020 68 8220 268
rect 8278 68 8478 268
rect 8536 68 8736 268
rect 8794 68 8994 268
rect 9246 68 9446 268
rect 9734 68 9934 268
rect 10186 68 10386 268
rect 10444 68 10644 268
rect 10702 68 10902 268
rect 10960 68 11160 268
rect 11412 68 11612 268
rect 11670 68 11870 268
rect 11928 68 12128 268
rect 12380 68 12580 268
rect 12638 68 12838 268
rect 12896 68 13096 268
rect 13154 68 13354 268
rect 13606 68 13806 268
rect 14092 68 14292 268
rect 14543 68 14743 268
rect 14801 68 15001 268
rect 15059 68 15259 268
rect 15317 68 15517 268
rect 15769 68 15969 268
rect 16027 68 16227 268
rect 16285 68 16485 268
rect 16737 68 16937 268
rect 16995 68 17195 268
rect 17253 68 17453 268
rect 17511 68 17711 268
rect 17963 68 18163 268
rect 1017 -876 1217 -676
rect 1469 -876 1669 -676
rect 1727 -876 1927 -676
rect 1985 -876 2185 -676
rect 2243 -876 2443 -676
rect 2695 -876 2895 -676
rect 2953 -876 3153 -676
rect 3211 -876 3411 -676
rect 3663 -876 3863 -676
rect 3921 -876 4121 -676
rect 4179 -876 4379 -676
rect 4437 -876 4637 -676
rect 4888 -876 5088 -676
rect 5374 -876 5574 -676
rect 5826 -876 6026 -676
rect 6084 -876 6284 -676
rect 6342 -876 6542 -676
rect 6600 -876 6800 -676
rect 7052 -876 7252 -676
rect 7310 -876 7510 -676
rect 7568 -876 7768 -676
rect 8020 -876 8220 -676
rect 8278 -876 8478 -676
rect 8536 -876 8736 -676
rect 8794 -876 8994 -676
rect 9246 -876 9446 -676
rect 9734 -876 9934 -676
rect 10186 -876 10386 -676
rect 10444 -876 10644 -676
rect 10702 -876 10902 -676
rect 10960 -876 11160 -676
rect 11412 -876 11612 -676
rect 11670 -876 11870 -676
rect 11928 -876 12128 -676
rect 12380 -876 12580 -676
rect 12638 -876 12838 -676
rect 12896 -876 13096 -676
rect 13154 -876 13354 -676
rect 13606 -876 13806 -676
rect 14092 -876 14292 -676
rect 14543 -876 14743 -676
rect 14801 -876 15001 -676
rect 15059 -876 15259 -676
rect 15317 -876 15517 -676
rect 15769 -876 15969 -676
rect 16027 -876 16227 -676
rect 16285 -876 16485 -676
rect 16737 -876 16937 -676
rect 16995 -876 17195 -676
rect 17253 -876 17453 -676
rect 17511 -876 17711 -676
rect 17963 -876 18163 -676
rect 1017 -1567 1217 -1367
rect 1469 -1567 1669 -1367
rect 1727 -1567 1927 -1367
rect 1985 -1567 2185 -1367
rect 2243 -1567 2443 -1367
rect 2695 -1567 2895 -1367
rect 2953 -1567 3153 -1367
rect 3211 -1567 3411 -1367
rect 3663 -1567 3863 -1367
rect 3921 -1567 4121 -1367
rect 4179 -1567 4379 -1367
rect 4437 -1567 4637 -1367
rect 4888 -1567 5088 -1367
rect 5374 -1567 5574 -1367
rect 5826 -1567 6026 -1367
rect 6084 -1567 6284 -1367
rect 6342 -1567 6542 -1367
rect 6600 -1567 6800 -1367
rect 7052 -1567 7252 -1367
rect 7310 -1567 7510 -1367
rect 7568 -1567 7768 -1367
rect 8020 -1567 8220 -1367
rect 8278 -1567 8478 -1367
rect 8536 -1567 8736 -1367
rect 8794 -1567 8994 -1367
rect 9246 -1567 9446 -1367
rect 9734 -1567 9934 -1367
rect 10186 -1567 10386 -1367
rect 10444 -1567 10644 -1367
rect 10702 -1567 10902 -1367
rect 10960 -1567 11160 -1367
rect 11412 -1567 11612 -1367
rect 11670 -1567 11870 -1367
rect 11928 -1567 12128 -1367
rect 12380 -1567 12580 -1367
rect 12638 -1567 12838 -1367
rect 12896 -1567 13096 -1367
rect 13154 -1567 13354 -1367
rect 13606 -1567 13806 -1367
rect 14092 -1567 14292 -1367
rect 14543 -1567 14743 -1367
rect 14801 -1567 15001 -1367
rect 15059 -1567 15259 -1367
rect 15317 -1567 15517 -1367
rect 15769 -1567 15969 -1367
rect 16027 -1567 16227 -1367
rect 16285 -1567 16485 -1367
rect 16737 -1567 16937 -1367
rect 16995 -1567 17195 -1367
rect 17253 -1567 17453 -1367
rect 17511 -1567 17711 -1367
rect 17963 -1567 18163 -1367
rect 1017 -2523 1217 -2323
rect 1469 -2523 1669 -2323
rect 1727 -2523 1927 -2323
rect 1985 -2523 2185 -2323
rect 2243 -2523 2443 -2323
rect 2695 -2523 2895 -2323
rect 2953 -2523 3153 -2323
rect 3211 -2523 3411 -2323
rect 3663 -2523 3863 -2323
rect 3921 -2523 4121 -2323
rect 4179 -2523 4379 -2323
rect 4437 -2523 4637 -2323
rect 4888 -2523 5088 -2323
rect 5374 -2523 5574 -2323
rect 5826 -2523 6026 -2323
rect 6084 -2523 6284 -2323
rect 6342 -2523 6542 -2323
rect 6600 -2523 6800 -2323
rect 7052 -2523 7252 -2323
rect 7310 -2523 7510 -2323
rect 7568 -2523 7768 -2323
rect 8020 -2523 8220 -2323
rect 8278 -2523 8478 -2323
rect 8536 -2523 8736 -2323
rect 8794 -2523 8994 -2323
rect 9246 -2523 9446 -2323
rect 9734 -2523 9934 -2323
rect 10186 -2523 10386 -2323
rect 10444 -2523 10644 -2323
rect 10702 -2523 10902 -2323
rect 10960 -2523 11160 -2323
rect 11412 -2523 11612 -2323
rect 11670 -2523 11870 -2323
rect 11928 -2523 12128 -2323
rect 12380 -2523 12580 -2323
rect 12638 -2523 12838 -2323
rect 12896 -2523 13096 -2323
rect 13154 -2523 13354 -2323
rect 13606 -2523 13806 -2323
rect 14092 -2523 14292 -2323
rect 14543 -2523 14743 -2323
rect 14801 -2523 15001 -2323
rect 15059 -2523 15259 -2323
rect 15317 -2523 15517 -2323
rect 15769 -2523 15969 -2323
rect 16027 -2523 16227 -2323
rect 16285 -2523 16485 -2323
rect 16737 -2523 16937 -2323
rect 16995 -2523 17195 -2323
rect 17253 -2523 17453 -2323
rect 17511 -2523 17711 -2323
rect 17963 -2523 18163 -2323
rect 1017 -3214 1217 -3014
rect 1469 -3214 1669 -3014
rect 1727 -3214 1927 -3014
rect 1985 -3214 2185 -3014
rect 2243 -3214 2443 -3014
rect 2695 -3214 2895 -3014
rect 2953 -3214 3153 -3014
rect 3211 -3214 3411 -3014
rect 3663 -3214 3863 -3014
rect 3921 -3214 4121 -3014
rect 4179 -3214 4379 -3014
rect 4437 -3214 4637 -3014
rect 4888 -3214 5088 -3014
rect 5374 -3214 5574 -3014
rect 5826 -3214 6026 -3014
rect 6084 -3214 6284 -3014
rect 6342 -3214 6542 -3014
rect 6600 -3214 6800 -3014
rect 7052 -3214 7252 -3014
rect 7310 -3214 7510 -3014
rect 7568 -3214 7768 -3014
rect 8020 -3214 8220 -3014
rect 8278 -3214 8478 -3014
rect 8536 -3214 8736 -3014
rect 8794 -3214 8994 -3014
rect 9246 -3214 9446 -3014
rect 9734 -3214 9934 -3014
rect 10186 -3214 10386 -3014
rect 10444 -3214 10644 -3014
rect 10702 -3214 10902 -3014
rect 10960 -3214 11160 -3014
rect 11412 -3214 11612 -3014
rect 11670 -3214 11870 -3014
rect 11928 -3214 12128 -3014
rect 12380 -3214 12580 -3014
rect 12638 -3214 12838 -3014
rect 12896 -3214 13096 -3014
rect 13154 -3214 13354 -3014
rect 13606 -3214 13806 -3014
rect 14092 -3214 14292 -3014
rect 14543 -3214 14743 -3014
rect 14801 -3214 15001 -3014
rect 15059 -3214 15259 -3014
rect 15317 -3214 15517 -3014
rect 15769 -3214 15969 -3014
rect 16027 -3214 16227 -3014
rect 16285 -3214 16485 -3014
rect 16737 -3214 16937 -3014
rect 16995 -3214 17195 -3014
rect 17253 -3214 17453 -3014
rect 17511 -3214 17711 -3014
rect 17963 -3214 18163 -3014
rect 1017 -4204 1217 -4004
rect 1469 -4204 1669 -4004
rect 1727 -4204 1927 -4004
rect 1985 -4204 2185 -4004
rect 2243 -4204 2443 -4004
rect 2695 -4204 2895 -4004
rect 2953 -4204 3153 -4004
rect 3211 -4204 3411 -4004
rect 3663 -4204 3863 -4004
rect 3921 -4204 4121 -4004
rect 4179 -4204 4379 -4004
rect 4437 -4204 4637 -4004
rect 4888 -4204 5088 -4004
rect 5374 -4204 5574 -4004
rect 5826 -4204 6026 -4004
rect 6084 -4204 6284 -4004
rect 6342 -4204 6542 -4004
rect 6600 -4204 6800 -4004
rect 7052 -4204 7252 -4004
rect 7310 -4204 7510 -4004
rect 7568 -4204 7768 -4004
rect 8020 -4204 8220 -4004
rect 8278 -4204 8478 -4004
rect 8536 -4204 8736 -4004
rect 8794 -4204 8994 -4004
rect 9246 -4204 9446 -4004
rect 9734 -4204 9934 -4004
rect 10186 -4204 10386 -4004
rect 10444 -4204 10644 -4004
rect 10702 -4204 10902 -4004
rect 10960 -4204 11160 -4004
rect 11412 -4204 11612 -4004
rect 11670 -4204 11870 -4004
rect 11928 -4204 12128 -4004
rect 12380 -4204 12580 -4004
rect 12638 -4204 12838 -4004
rect 12896 -4204 13096 -4004
rect 13154 -4204 13354 -4004
rect 13606 -4204 13806 -4004
rect 14092 -4204 14292 -4004
rect 14543 -4204 14743 -4004
rect 14801 -4204 15001 -4004
rect 15059 -4204 15259 -4004
rect 15317 -4204 15517 -4004
rect 15769 -4204 15969 -4004
rect 16027 -4204 16227 -4004
rect 16285 -4204 16485 -4004
rect 16737 -4204 16937 -4004
rect 16995 -4204 17195 -4004
rect 17253 -4204 17453 -4004
rect 17511 -4204 17711 -4004
rect 17963 -4204 18163 -4004
rect 1017 -4760 1217 -4560
rect 1469 -4760 1669 -4560
rect 1727 -4760 1927 -4560
rect 1985 -4760 2185 -4560
rect 2243 -4760 2443 -4560
rect 2695 -4760 2895 -4560
rect 2953 -4760 3153 -4560
rect 3211 -4760 3411 -4560
rect 3663 -4760 3863 -4560
rect 3921 -4760 4121 -4560
rect 4179 -4760 4379 -4560
rect 4437 -4760 4637 -4560
rect 4888 -4760 5088 -4560
rect 5374 -4760 5574 -4560
rect 5826 -4760 6026 -4560
rect 6084 -4760 6284 -4560
rect 6342 -4760 6542 -4560
rect 6600 -4760 6800 -4560
rect 7052 -4760 7252 -4560
rect 7310 -4760 7510 -4560
rect 7568 -4760 7768 -4560
rect 8020 -4760 8220 -4560
rect 8278 -4760 8478 -4560
rect 8536 -4760 8736 -4560
rect 8794 -4760 8994 -4560
rect 9246 -4760 9446 -4560
rect 9734 -4760 9934 -4560
rect 10186 -4760 10386 -4560
rect 10444 -4760 10644 -4560
rect 10702 -4760 10902 -4560
rect 10960 -4760 11160 -4560
rect 11412 -4760 11612 -4560
rect 11670 -4760 11870 -4560
rect 11928 -4760 12128 -4560
rect 12380 -4760 12580 -4560
rect 12638 -4760 12838 -4560
rect 12896 -4760 13096 -4560
rect 13154 -4760 13354 -4560
rect 13606 -4760 13806 -4560
rect 14092 -4760 14292 -4560
rect 14543 -4760 14743 -4560
rect 14801 -4760 15001 -4560
rect 15059 -4760 15259 -4560
rect 15317 -4760 15517 -4560
rect 15769 -4760 15969 -4560
rect 16027 -4760 16227 -4560
rect 16285 -4760 16485 -4560
rect 16737 -4760 16937 -4560
rect 16995 -4760 17195 -4560
rect 17253 -4760 17453 -4560
rect 17511 -4760 17711 -4560
rect 17963 -4760 18163 -4560
rect 1017 -5750 1217 -5550
rect 1469 -5750 1669 -5550
rect 1727 -5750 1927 -5550
rect 1985 -5750 2185 -5550
rect 2243 -5750 2443 -5550
rect 2695 -5750 2895 -5550
rect 2953 -5750 3153 -5550
rect 3211 -5750 3411 -5550
rect 3663 -5750 3863 -5550
rect 3921 -5750 4121 -5550
rect 4179 -5750 4379 -5550
rect 4437 -5750 4637 -5550
rect 4888 -5750 5088 -5550
rect 5374 -5750 5574 -5550
rect 5826 -5750 6026 -5550
rect 6084 -5750 6284 -5550
rect 6342 -5750 6542 -5550
rect 6600 -5750 6800 -5550
rect 7052 -5750 7252 -5550
rect 7310 -5750 7510 -5550
rect 7568 -5750 7768 -5550
rect 8020 -5750 8220 -5550
rect 8278 -5750 8478 -5550
rect 8536 -5750 8736 -5550
rect 8794 -5750 8994 -5550
rect 9246 -5750 9446 -5550
rect 9734 -5750 9934 -5550
rect 10186 -5750 10386 -5550
rect 10444 -5750 10644 -5550
rect 10702 -5750 10902 -5550
rect 10960 -5750 11160 -5550
rect 11412 -5750 11612 -5550
rect 11670 -5750 11870 -5550
rect 11928 -5750 12128 -5550
rect 12380 -5750 12580 -5550
rect 12638 -5750 12838 -5550
rect 12896 -5750 13096 -5550
rect 13154 -5750 13354 -5550
rect 13606 -5750 13806 -5550
rect 14092 -5750 14292 -5550
rect 14543 -5750 14743 -5550
rect 14801 -5750 15001 -5550
rect 15059 -5750 15259 -5550
rect 15317 -5750 15517 -5550
rect 15769 -5750 15969 -5550
rect 16027 -5750 16227 -5550
rect 16285 -5750 16485 -5550
rect 16737 -5750 16937 -5550
rect 16995 -5750 17195 -5550
rect 17253 -5750 17453 -5550
rect 17511 -5750 17711 -5550
rect 17963 -5750 18163 -5550
rect 1017 -6440 1217 -6240
rect 1469 -6440 1669 -6240
rect 1727 -6440 1927 -6240
rect 1985 -6440 2185 -6240
rect 2243 -6440 2443 -6240
rect 2695 -6440 2895 -6240
rect 2953 -6440 3153 -6240
rect 3211 -6440 3411 -6240
rect 3663 -6440 3863 -6240
rect 3921 -6440 4121 -6240
rect 4179 -6440 4379 -6240
rect 4437 -6440 4637 -6240
rect 4888 -6440 5088 -6240
rect 5374 -6440 5574 -6240
rect 5826 -6440 6026 -6240
rect 6084 -6440 6284 -6240
rect 6342 -6440 6542 -6240
rect 6600 -6440 6800 -6240
rect 7052 -6440 7252 -6240
rect 7310 -6440 7510 -6240
rect 7568 -6440 7768 -6240
rect 8020 -6440 8220 -6240
rect 8278 -6440 8478 -6240
rect 8536 -6440 8736 -6240
rect 8794 -6440 8994 -6240
rect 9246 -6440 9446 -6240
rect 9734 -6440 9934 -6240
rect 10186 -6440 10386 -6240
rect 10444 -6440 10644 -6240
rect 10702 -6440 10902 -6240
rect 10960 -6440 11160 -6240
rect 11412 -6440 11612 -6240
rect 11670 -6440 11870 -6240
rect 11928 -6440 12128 -6240
rect 12380 -6440 12580 -6240
rect 12638 -6440 12838 -6240
rect 12896 -6440 13096 -6240
rect 13154 -6440 13354 -6240
rect 13606 -6440 13806 -6240
rect 14092 -6440 14292 -6240
rect 14543 -6440 14743 -6240
rect 14801 -6440 15001 -6240
rect 15059 -6440 15259 -6240
rect 15317 -6440 15517 -6240
rect 15769 -6440 15969 -6240
rect 16027 -6440 16227 -6240
rect 16285 -6440 16485 -6240
rect 16737 -6440 16937 -6240
rect 16995 -6440 17195 -6240
rect 17253 -6440 17453 -6240
rect 17511 -6440 17711 -6240
rect 17963 -6440 18163 -6240
rect 1017 -7397 1217 -7197
rect 1469 -7397 1669 -7197
rect 1727 -7397 1927 -7197
rect 1985 -7397 2185 -7197
rect 2243 -7397 2443 -7197
rect 2695 -7397 2895 -7197
rect 2953 -7397 3153 -7197
rect 3211 -7397 3411 -7197
rect 3663 -7397 3863 -7197
rect 3921 -7397 4121 -7197
rect 4179 -7397 4379 -7197
rect 4437 -7397 4637 -7197
rect 4888 -7397 5088 -7197
rect 5374 -7397 5574 -7197
rect 5826 -7397 6026 -7197
rect 6084 -7397 6284 -7197
rect 6342 -7397 6542 -7197
rect 6600 -7397 6800 -7197
rect 7052 -7397 7252 -7197
rect 7310 -7397 7510 -7197
rect 7568 -7397 7768 -7197
rect 8020 -7397 8220 -7197
rect 8278 -7397 8478 -7197
rect 8536 -7397 8736 -7197
rect 8794 -7397 8994 -7197
rect 9246 -7397 9446 -7197
rect 9734 -7397 9934 -7197
rect 10186 -7397 10386 -7197
rect 10444 -7397 10644 -7197
rect 10702 -7397 10902 -7197
rect 10960 -7397 11160 -7197
rect 11412 -7397 11612 -7197
rect 11670 -7397 11870 -7197
rect 11928 -7397 12128 -7197
rect 12380 -7397 12580 -7197
rect 12638 -7397 12838 -7197
rect 12896 -7397 13096 -7197
rect 13154 -7397 13354 -7197
rect 13606 -7397 13806 -7197
rect 14092 -7397 14292 -7197
rect 14543 -7397 14743 -7197
rect 14801 -7397 15001 -7197
rect 15059 -7397 15259 -7197
rect 15317 -7397 15517 -7197
rect 15769 -7397 15969 -7197
rect 16027 -7397 16227 -7197
rect 16285 -7397 16485 -7197
rect 16737 -7397 16937 -7197
rect 16995 -7397 17195 -7197
rect 17253 -7397 17453 -7197
rect 17511 -7397 17711 -7197
rect 17963 -7397 18163 -7197
rect 1017 -8087 1217 -7887
rect 1469 -8087 1669 -7887
rect 1727 -8087 1927 -7887
rect 1985 -8087 2185 -7887
rect 2243 -8087 2443 -7887
rect 2695 -8087 2895 -7887
rect 2953 -8087 3153 -7887
rect 3211 -8087 3411 -7887
rect 3663 -8087 3863 -7887
rect 3921 -8087 4121 -7887
rect 4179 -8087 4379 -7887
rect 4437 -8087 4637 -7887
rect 4888 -8087 5088 -7887
rect 5374 -8087 5574 -7887
rect 5826 -8087 6026 -7887
rect 6084 -8087 6284 -7887
rect 6342 -8087 6542 -7887
rect 6600 -8087 6800 -7887
rect 7052 -8087 7252 -7887
rect 7310 -8087 7510 -7887
rect 7568 -8087 7768 -7887
rect 8020 -8087 8220 -7887
rect 8278 -8087 8478 -7887
rect 8536 -8087 8736 -7887
rect 8794 -8087 8994 -7887
rect 9246 -8087 9446 -7887
rect 9734 -8087 9934 -7887
rect 10186 -8087 10386 -7887
rect 10444 -8087 10644 -7887
rect 10702 -8087 10902 -7887
rect 10960 -8087 11160 -7887
rect 11412 -8087 11612 -7887
rect 11670 -8087 11870 -7887
rect 11928 -8087 12128 -7887
rect 12380 -8087 12580 -7887
rect 12638 -8087 12838 -7887
rect 12896 -8087 13096 -7887
rect 13154 -8087 13354 -7887
rect 13606 -8087 13806 -7887
rect 14092 -8087 14292 -7887
rect 14543 -8087 14743 -7887
rect 14801 -8087 15001 -7887
rect 15059 -8087 15259 -7887
rect 15317 -8087 15517 -7887
rect 15769 -8087 15969 -7887
rect 16027 -8087 16227 -7887
rect 16285 -8087 16485 -7887
rect 16737 -8087 16937 -7887
rect 16995 -8087 17195 -7887
rect 17253 -8087 17453 -7887
rect 17511 -8087 17711 -7887
rect 17963 -8087 18163 -7887
rect 1017 -9031 1217 -8831
rect 1469 -9031 1669 -8831
rect 1727 -9031 1927 -8831
rect 1985 -9031 2185 -8831
rect 2243 -9031 2443 -8831
rect 2695 -9031 2895 -8831
rect 2953 -9031 3153 -8831
rect 3211 -9031 3411 -8831
rect 3663 -9031 3863 -8831
rect 3921 -9031 4121 -8831
rect 4179 -9031 4379 -8831
rect 4437 -9031 4637 -8831
rect 4888 -9031 5088 -8831
rect 5374 -9031 5574 -8831
rect 5826 -9031 6026 -8831
rect 6084 -9031 6284 -8831
rect 6342 -9031 6542 -8831
rect 6600 -9031 6800 -8831
rect 7052 -9031 7252 -8831
rect 7310 -9031 7510 -8831
rect 7568 -9031 7768 -8831
rect 8020 -9031 8220 -8831
rect 8278 -9031 8478 -8831
rect 8536 -9031 8736 -8831
rect 8794 -9031 8994 -8831
rect 9246 -9031 9446 -8831
rect 9734 -9031 9934 -8831
rect 10186 -9031 10386 -8831
rect 10444 -9031 10644 -8831
rect 10702 -9031 10902 -8831
rect 10960 -9031 11160 -8831
rect 11412 -9031 11612 -8831
rect 11670 -9031 11870 -8831
rect 11928 -9031 12128 -8831
rect 12380 -9031 12580 -8831
rect 12638 -9031 12838 -8831
rect 12896 -9031 13096 -8831
rect 13154 -9031 13354 -8831
rect 13606 -9031 13806 -8831
rect 14092 -9031 14292 -8831
rect 14543 -9031 14743 -8831
rect 14801 -9031 15001 -8831
rect 15059 -9031 15259 -8831
rect 15317 -9031 15517 -8831
rect 15769 -9031 15969 -8831
rect 16027 -9031 16227 -8831
rect 16285 -9031 16485 -8831
rect 16737 -9031 16937 -8831
rect 16995 -9031 17195 -8831
rect 17253 -9031 17453 -8831
rect 17511 -9031 17711 -8831
rect 17963 -9031 18163 -8831
<< pdiff >>
rect 959 253 1017 268
rect 959 219 971 253
rect 1005 219 1017 253
rect 959 185 1017 219
rect 959 151 971 185
rect 1005 151 1017 185
rect 959 117 1017 151
rect 959 83 971 117
rect 1005 83 1017 117
rect 959 68 1017 83
rect 1217 253 1275 268
rect 1217 219 1229 253
rect 1263 219 1275 253
rect 1217 185 1275 219
rect 1217 151 1229 185
rect 1263 151 1275 185
rect 1217 117 1275 151
rect 1217 83 1229 117
rect 1263 83 1275 117
rect 1217 68 1275 83
rect 1411 253 1469 268
rect 1411 219 1423 253
rect 1457 219 1469 253
rect 1411 185 1469 219
rect 1411 151 1423 185
rect 1457 151 1469 185
rect 1411 117 1469 151
rect 1411 83 1423 117
rect 1457 83 1469 117
rect 1411 68 1469 83
rect 1669 253 1727 268
rect 1669 219 1681 253
rect 1715 219 1727 253
rect 1669 185 1727 219
rect 1669 151 1681 185
rect 1715 151 1727 185
rect 1669 117 1727 151
rect 1669 83 1681 117
rect 1715 83 1727 117
rect 1669 68 1727 83
rect 1927 253 1985 268
rect 1927 219 1939 253
rect 1973 219 1985 253
rect 1927 185 1985 219
rect 1927 151 1939 185
rect 1973 151 1985 185
rect 1927 117 1985 151
rect 1927 83 1939 117
rect 1973 83 1985 117
rect 1927 68 1985 83
rect 2185 253 2243 268
rect 2185 219 2197 253
rect 2231 219 2243 253
rect 2185 185 2243 219
rect 2185 151 2197 185
rect 2231 151 2243 185
rect 2185 117 2243 151
rect 2185 83 2197 117
rect 2231 83 2243 117
rect 2185 68 2243 83
rect 2443 253 2501 268
rect 2443 219 2455 253
rect 2489 219 2501 253
rect 2443 185 2501 219
rect 2443 151 2455 185
rect 2489 151 2501 185
rect 2443 117 2501 151
rect 2443 83 2455 117
rect 2489 83 2501 117
rect 2443 68 2501 83
rect 2637 253 2695 268
rect 2637 219 2649 253
rect 2683 219 2695 253
rect 2637 185 2695 219
rect 2637 151 2649 185
rect 2683 151 2695 185
rect 2637 117 2695 151
rect 2637 83 2649 117
rect 2683 83 2695 117
rect 2637 68 2695 83
rect 2895 253 2953 268
rect 2895 219 2907 253
rect 2941 219 2953 253
rect 2895 185 2953 219
rect 2895 151 2907 185
rect 2941 151 2953 185
rect 2895 117 2953 151
rect 2895 83 2907 117
rect 2941 83 2953 117
rect 2895 68 2953 83
rect 3153 253 3211 268
rect 3153 219 3165 253
rect 3199 219 3211 253
rect 3153 185 3211 219
rect 3153 151 3165 185
rect 3199 151 3211 185
rect 3153 117 3211 151
rect 3153 83 3165 117
rect 3199 83 3211 117
rect 3153 68 3211 83
rect 3411 253 3469 268
rect 3411 219 3423 253
rect 3457 219 3469 253
rect 3411 185 3469 219
rect 3411 151 3423 185
rect 3457 151 3469 185
rect 3411 117 3469 151
rect 3411 83 3423 117
rect 3457 83 3469 117
rect 3411 68 3469 83
rect 3605 253 3663 268
rect 3605 219 3617 253
rect 3651 219 3663 253
rect 3605 185 3663 219
rect 3605 151 3617 185
rect 3651 151 3663 185
rect 3605 117 3663 151
rect 3605 83 3617 117
rect 3651 83 3663 117
rect 3605 68 3663 83
rect 3863 253 3921 268
rect 3863 219 3875 253
rect 3909 219 3921 253
rect 3863 185 3921 219
rect 3863 151 3875 185
rect 3909 151 3921 185
rect 3863 117 3921 151
rect 3863 83 3875 117
rect 3909 83 3921 117
rect 3863 68 3921 83
rect 4121 253 4179 268
rect 4121 219 4133 253
rect 4167 219 4179 253
rect 4121 185 4179 219
rect 4121 151 4133 185
rect 4167 151 4179 185
rect 4121 117 4179 151
rect 4121 83 4133 117
rect 4167 83 4179 117
rect 4121 68 4179 83
rect 4379 253 4437 268
rect 4379 219 4391 253
rect 4425 219 4437 253
rect 4379 185 4437 219
rect 4379 151 4391 185
rect 4425 151 4437 185
rect 4379 117 4437 151
rect 4379 83 4391 117
rect 4425 83 4437 117
rect 4379 68 4437 83
rect 4637 253 4695 268
rect 4637 219 4649 253
rect 4683 219 4695 253
rect 4637 185 4695 219
rect 4637 151 4649 185
rect 4683 151 4695 185
rect 4637 117 4695 151
rect 4637 83 4649 117
rect 4683 83 4695 117
rect 4637 68 4695 83
rect 4830 253 4888 268
rect 4830 219 4842 253
rect 4876 219 4888 253
rect 4830 185 4888 219
rect 4830 151 4842 185
rect 4876 151 4888 185
rect 4830 117 4888 151
rect 4830 83 4842 117
rect 4876 83 4888 117
rect 4830 68 4888 83
rect 5088 253 5146 268
rect 5088 219 5100 253
rect 5134 219 5146 253
rect 5088 185 5146 219
rect 5088 151 5100 185
rect 5134 151 5146 185
rect 5088 117 5146 151
rect 5088 83 5100 117
rect 5134 83 5146 117
rect 5088 68 5146 83
rect 5316 253 5374 268
rect 5316 219 5328 253
rect 5362 219 5374 253
rect 5316 185 5374 219
rect 5316 151 5328 185
rect 5362 151 5374 185
rect 5316 117 5374 151
rect 5316 83 5328 117
rect 5362 83 5374 117
rect 5316 68 5374 83
rect 5574 253 5632 268
rect 5574 219 5586 253
rect 5620 219 5632 253
rect 5574 185 5632 219
rect 5574 151 5586 185
rect 5620 151 5632 185
rect 5574 117 5632 151
rect 5574 83 5586 117
rect 5620 83 5632 117
rect 5574 68 5632 83
rect 5768 253 5826 268
rect 5768 219 5780 253
rect 5814 219 5826 253
rect 5768 185 5826 219
rect 5768 151 5780 185
rect 5814 151 5826 185
rect 5768 117 5826 151
rect 5768 83 5780 117
rect 5814 83 5826 117
rect 5768 68 5826 83
rect 6026 253 6084 268
rect 6026 219 6038 253
rect 6072 219 6084 253
rect 6026 185 6084 219
rect 6026 151 6038 185
rect 6072 151 6084 185
rect 6026 117 6084 151
rect 6026 83 6038 117
rect 6072 83 6084 117
rect 6026 68 6084 83
rect 6284 253 6342 268
rect 6284 219 6296 253
rect 6330 219 6342 253
rect 6284 185 6342 219
rect 6284 151 6296 185
rect 6330 151 6342 185
rect 6284 117 6342 151
rect 6284 83 6296 117
rect 6330 83 6342 117
rect 6284 68 6342 83
rect 6542 253 6600 268
rect 6542 219 6554 253
rect 6588 219 6600 253
rect 6542 185 6600 219
rect 6542 151 6554 185
rect 6588 151 6600 185
rect 6542 117 6600 151
rect 6542 83 6554 117
rect 6588 83 6600 117
rect 6542 68 6600 83
rect 6800 253 6858 268
rect 6800 219 6812 253
rect 6846 219 6858 253
rect 6800 185 6858 219
rect 6800 151 6812 185
rect 6846 151 6858 185
rect 6800 117 6858 151
rect 6800 83 6812 117
rect 6846 83 6858 117
rect 6800 68 6858 83
rect 6994 253 7052 268
rect 6994 219 7006 253
rect 7040 219 7052 253
rect 6994 185 7052 219
rect 6994 151 7006 185
rect 7040 151 7052 185
rect 6994 117 7052 151
rect 6994 83 7006 117
rect 7040 83 7052 117
rect 6994 68 7052 83
rect 7252 253 7310 268
rect 7252 219 7264 253
rect 7298 219 7310 253
rect 7252 185 7310 219
rect 7252 151 7264 185
rect 7298 151 7310 185
rect 7252 117 7310 151
rect 7252 83 7264 117
rect 7298 83 7310 117
rect 7252 68 7310 83
rect 7510 253 7568 268
rect 7510 219 7522 253
rect 7556 219 7568 253
rect 7510 185 7568 219
rect 7510 151 7522 185
rect 7556 151 7568 185
rect 7510 117 7568 151
rect 7510 83 7522 117
rect 7556 83 7568 117
rect 7510 68 7568 83
rect 7768 253 7826 268
rect 7768 219 7780 253
rect 7814 219 7826 253
rect 7768 185 7826 219
rect 7768 151 7780 185
rect 7814 151 7826 185
rect 7768 117 7826 151
rect 7768 83 7780 117
rect 7814 83 7826 117
rect 7768 68 7826 83
rect 7962 253 8020 268
rect 7962 219 7974 253
rect 8008 219 8020 253
rect 7962 185 8020 219
rect 7962 151 7974 185
rect 8008 151 8020 185
rect 7962 117 8020 151
rect 7962 83 7974 117
rect 8008 83 8020 117
rect 7962 68 8020 83
rect 8220 253 8278 268
rect 8220 219 8232 253
rect 8266 219 8278 253
rect 8220 185 8278 219
rect 8220 151 8232 185
rect 8266 151 8278 185
rect 8220 117 8278 151
rect 8220 83 8232 117
rect 8266 83 8278 117
rect 8220 68 8278 83
rect 8478 253 8536 268
rect 8478 219 8490 253
rect 8524 219 8536 253
rect 8478 185 8536 219
rect 8478 151 8490 185
rect 8524 151 8536 185
rect 8478 117 8536 151
rect 8478 83 8490 117
rect 8524 83 8536 117
rect 8478 68 8536 83
rect 8736 253 8794 268
rect 8736 219 8748 253
rect 8782 219 8794 253
rect 8736 185 8794 219
rect 8736 151 8748 185
rect 8782 151 8794 185
rect 8736 117 8794 151
rect 8736 83 8748 117
rect 8782 83 8794 117
rect 8736 68 8794 83
rect 8994 253 9052 268
rect 8994 219 9006 253
rect 9040 219 9052 253
rect 8994 185 9052 219
rect 8994 151 9006 185
rect 9040 151 9052 185
rect 8994 117 9052 151
rect 8994 83 9006 117
rect 9040 83 9052 117
rect 8994 68 9052 83
rect 9188 253 9246 268
rect 9188 219 9200 253
rect 9234 219 9246 253
rect 9188 185 9246 219
rect 9188 151 9200 185
rect 9234 151 9246 185
rect 9188 117 9246 151
rect 9188 83 9200 117
rect 9234 83 9246 117
rect 9188 68 9246 83
rect 9446 253 9504 268
rect 9446 219 9458 253
rect 9492 219 9504 253
rect 9446 185 9504 219
rect 9446 151 9458 185
rect 9492 151 9504 185
rect 9446 117 9504 151
rect 9446 83 9458 117
rect 9492 83 9504 117
rect 9446 68 9504 83
rect 9676 253 9734 268
rect 9676 219 9688 253
rect 9722 219 9734 253
rect 9676 185 9734 219
rect 9676 151 9688 185
rect 9722 151 9734 185
rect 9676 117 9734 151
rect 9676 83 9688 117
rect 9722 83 9734 117
rect 9676 68 9734 83
rect 9934 253 9992 268
rect 9934 219 9946 253
rect 9980 219 9992 253
rect 9934 185 9992 219
rect 9934 151 9946 185
rect 9980 151 9992 185
rect 9934 117 9992 151
rect 9934 83 9946 117
rect 9980 83 9992 117
rect 9934 68 9992 83
rect 10128 253 10186 268
rect 10128 219 10140 253
rect 10174 219 10186 253
rect 10128 185 10186 219
rect 10128 151 10140 185
rect 10174 151 10186 185
rect 10128 117 10186 151
rect 10128 83 10140 117
rect 10174 83 10186 117
rect 10128 68 10186 83
rect 10386 253 10444 268
rect 10386 219 10398 253
rect 10432 219 10444 253
rect 10386 185 10444 219
rect 10386 151 10398 185
rect 10432 151 10444 185
rect 10386 117 10444 151
rect 10386 83 10398 117
rect 10432 83 10444 117
rect 10386 68 10444 83
rect 10644 253 10702 268
rect 10644 219 10656 253
rect 10690 219 10702 253
rect 10644 185 10702 219
rect 10644 151 10656 185
rect 10690 151 10702 185
rect 10644 117 10702 151
rect 10644 83 10656 117
rect 10690 83 10702 117
rect 10644 68 10702 83
rect 10902 253 10960 268
rect 10902 219 10914 253
rect 10948 219 10960 253
rect 10902 185 10960 219
rect 10902 151 10914 185
rect 10948 151 10960 185
rect 10902 117 10960 151
rect 10902 83 10914 117
rect 10948 83 10960 117
rect 10902 68 10960 83
rect 11160 253 11218 268
rect 11160 219 11172 253
rect 11206 219 11218 253
rect 11160 185 11218 219
rect 11160 151 11172 185
rect 11206 151 11218 185
rect 11160 117 11218 151
rect 11160 83 11172 117
rect 11206 83 11218 117
rect 11160 68 11218 83
rect 11354 253 11412 268
rect 11354 219 11366 253
rect 11400 219 11412 253
rect 11354 185 11412 219
rect 11354 151 11366 185
rect 11400 151 11412 185
rect 11354 117 11412 151
rect 11354 83 11366 117
rect 11400 83 11412 117
rect 11354 68 11412 83
rect 11612 253 11670 268
rect 11612 219 11624 253
rect 11658 219 11670 253
rect 11612 185 11670 219
rect 11612 151 11624 185
rect 11658 151 11670 185
rect 11612 117 11670 151
rect 11612 83 11624 117
rect 11658 83 11670 117
rect 11612 68 11670 83
rect 11870 253 11928 268
rect 11870 219 11882 253
rect 11916 219 11928 253
rect 11870 185 11928 219
rect 11870 151 11882 185
rect 11916 151 11928 185
rect 11870 117 11928 151
rect 11870 83 11882 117
rect 11916 83 11928 117
rect 11870 68 11928 83
rect 12128 253 12186 268
rect 12128 219 12140 253
rect 12174 219 12186 253
rect 12128 185 12186 219
rect 12128 151 12140 185
rect 12174 151 12186 185
rect 12128 117 12186 151
rect 12128 83 12140 117
rect 12174 83 12186 117
rect 12128 68 12186 83
rect 12322 253 12380 268
rect 12322 219 12334 253
rect 12368 219 12380 253
rect 12322 185 12380 219
rect 12322 151 12334 185
rect 12368 151 12380 185
rect 12322 117 12380 151
rect 12322 83 12334 117
rect 12368 83 12380 117
rect 12322 68 12380 83
rect 12580 253 12638 268
rect 12580 219 12592 253
rect 12626 219 12638 253
rect 12580 185 12638 219
rect 12580 151 12592 185
rect 12626 151 12638 185
rect 12580 117 12638 151
rect 12580 83 12592 117
rect 12626 83 12638 117
rect 12580 68 12638 83
rect 12838 253 12896 268
rect 12838 219 12850 253
rect 12884 219 12896 253
rect 12838 185 12896 219
rect 12838 151 12850 185
rect 12884 151 12896 185
rect 12838 117 12896 151
rect 12838 83 12850 117
rect 12884 83 12896 117
rect 12838 68 12896 83
rect 13096 253 13154 268
rect 13096 219 13108 253
rect 13142 219 13154 253
rect 13096 185 13154 219
rect 13096 151 13108 185
rect 13142 151 13154 185
rect 13096 117 13154 151
rect 13096 83 13108 117
rect 13142 83 13154 117
rect 13096 68 13154 83
rect 13354 253 13412 268
rect 13354 219 13366 253
rect 13400 219 13412 253
rect 13354 185 13412 219
rect 13354 151 13366 185
rect 13400 151 13412 185
rect 13354 117 13412 151
rect 13354 83 13366 117
rect 13400 83 13412 117
rect 13354 68 13412 83
rect 13548 253 13606 268
rect 13548 219 13560 253
rect 13594 219 13606 253
rect 13548 185 13606 219
rect 13548 151 13560 185
rect 13594 151 13606 185
rect 13548 117 13606 151
rect 13548 83 13560 117
rect 13594 83 13606 117
rect 13548 68 13606 83
rect 13806 253 13864 268
rect 13806 219 13818 253
rect 13852 219 13864 253
rect 13806 185 13864 219
rect 13806 151 13818 185
rect 13852 151 13864 185
rect 13806 117 13864 151
rect 13806 83 13818 117
rect 13852 83 13864 117
rect 13806 68 13864 83
rect 14034 253 14092 268
rect 14034 219 14046 253
rect 14080 219 14092 253
rect 14034 185 14092 219
rect 14034 151 14046 185
rect 14080 151 14092 185
rect 14034 117 14092 151
rect 14034 83 14046 117
rect 14080 83 14092 117
rect 14034 68 14092 83
rect 14292 253 14350 268
rect 14292 219 14304 253
rect 14338 219 14350 253
rect 14292 185 14350 219
rect 14292 151 14304 185
rect 14338 151 14350 185
rect 14292 117 14350 151
rect 14292 83 14304 117
rect 14338 83 14350 117
rect 14292 68 14350 83
rect 14485 253 14543 268
rect 14485 219 14497 253
rect 14531 219 14543 253
rect 14485 185 14543 219
rect 14485 151 14497 185
rect 14531 151 14543 185
rect 14485 117 14543 151
rect 14485 83 14497 117
rect 14531 83 14543 117
rect 14485 68 14543 83
rect 14743 253 14801 268
rect 14743 219 14755 253
rect 14789 219 14801 253
rect 14743 185 14801 219
rect 14743 151 14755 185
rect 14789 151 14801 185
rect 14743 117 14801 151
rect 14743 83 14755 117
rect 14789 83 14801 117
rect 14743 68 14801 83
rect 15001 253 15059 268
rect 15001 219 15013 253
rect 15047 219 15059 253
rect 15001 185 15059 219
rect 15001 151 15013 185
rect 15047 151 15059 185
rect 15001 117 15059 151
rect 15001 83 15013 117
rect 15047 83 15059 117
rect 15001 68 15059 83
rect 15259 253 15317 268
rect 15259 219 15271 253
rect 15305 219 15317 253
rect 15259 185 15317 219
rect 15259 151 15271 185
rect 15305 151 15317 185
rect 15259 117 15317 151
rect 15259 83 15271 117
rect 15305 83 15317 117
rect 15259 68 15317 83
rect 15517 253 15575 268
rect 15517 219 15529 253
rect 15563 219 15575 253
rect 15517 185 15575 219
rect 15517 151 15529 185
rect 15563 151 15575 185
rect 15517 117 15575 151
rect 15517 83 15529 117
rect 15563 83 15575 117
rect 15517 68 15575 83
rect 15711 253 15769 268
rect 15711 219 15723 253
rect 15757 219 15769 253
rect 15711 185 15769 219
rect 15711 151 15723 185
rect 15757 151 15769 185
rect 15711 117 15769 151
rect 15711 83 15723 117
rect 15757 83 15769 117
rect 15711 68 15769 83
rect 15969 253 16027 268
rect 15969 219 15981 253
rect 16015 219 16027 253
rect 15969 185 16027 219
rect 15969 151 15981 185
rect 16015 151 16027 185
rect 15969 117 16027 151
rect 15969 83 15981 117
rect 16015 83 16027 117
rect 15969 68 16027 83
rect 16227 253 16285 268
rect 16227 219 16239 253
rect 16273 219 16285 253
rect 16227 185 16285 219
rect 16227 151 16239 185
rect 16273 151 16285 185
rect 16227 117 16285 151
rect 16227 83 16239 117
rect 16273 83 16285 117
rect 16227 68 16285 83
rect 16485 253 16543 268
rect 16485 219 16497 253
rect 16531 219 16543 253
rect 16485 185 16543 219
rect 16485 151 16497 185
rect 16531 151 16543 185
rect 16485 117 16543 151
rect 16485 83 16497 117
rect 16531 83 16543 117
rect 16485 68 16543 83
rect 16679 253 16737 268
rect 16679 219 16691 253
rect 16725 219 16737 253
rect 16679 185 16737 219
rect 16679 151 16691 185
rect 16725 151 16737 185
rect 16679 117 16737 151
rect 16679 83 16691 117
rect 16725 83 16737 117
rect 16679 68 16737 83
rect 16937 253 16995 268
rect 16937 219 16949 253
rect 16983 219 16995 253
rect 16937 185 16995 219
rect 16937 151 16949 185
rect 16983 151 16995 185
rect 16937 117 16995 151
rect 16937 83 16949 117
rect 16983 83 16995 117
rect 16937 68 16995 83
rect 17195 253 17253 268
rect 17195 219 17207 253
rect 17241 219 17253 253
rect 17195 185 17253 219
rect 17195 151 17207 185
rect 17241 151 17253 185
rect 17195 117 17253 151
rect 17195 83 17207 117
rect 17241 83 17253 117
rect 17195 68 17253 83
rect 17453 253 17511 268
rect 17453 219 17465 253
rect 17499 219 17511 253
rect 17453 185 17511 219
rect 17453 151 17465 185
rect 17499 151 17511 185
rect 17453 117 17511 151
rect 17453 83 17465 117
rect 17499 83 17511 117
rect 17453 68 17511 83
rect 17711 253 17769 268
rect 17711 219 17723 253
rect 17757 219 17769 253
rect 17711 185 17769 219
rect 17711 151 17723 185
rect 17757 151 17769 185
rect 17711 117 17769 151
rect 17711 83 17723 117
rect 17757 83 17769 117
rect 17711 68 17769 83
rect 17905 253 17963 268
rect 17905 219 17917 253
rect 17951 219 17963 253
rect 17905 185 17963 219
rect 17905 151 17917 185
rect 17951 151 17963 185
rect 17905 117 17963 151
rect 17905 83 17917 117
rect 17951 83 17963 117
rect 17905 68 17963 83
rect 18163 253 18221 268
rect 18163 219 18175 253
rect 18209 219 18221 253
rect 18163 185 18221 219
rect 18163 151 18175 185
rect 18209 151 18221 185
rect 18163 117 18221 151
rect 18163 83 18175 117
rect 18209 83 18221 117
rect 18163 68 18221 83
rect 959 -691 1017 -676
rect 959 -725 971 -691
rect 1005 -725 1017 -691
rect 959 -759 1017 -725
rect 959 -793 971 -759
rect 1005 -793 1017 -759
rect 959 -827 1017 -793
rect 959 -861 971 -827
rect 1005 -861 1017 -827
rect 959 -876 1017 -861
rect 1217 -691 1275 -676
rect 1217 -725 1229 -691
rect 1263 -725 1275 -691
rect 1217 -759 1275 -725
rect 1217 -793 1229 -759
rect 1263 -793 1275 -759
rect 1217 -827 1275 -793
rect 1217 -861 1229 -827
rect 1263 -861 1275 -827
rect 1217 -876 1275 -861
rect 1411 -691 1469 -676
rect 1411 -725 1423 -691
rect 1457 -725 1469 -691
rect 1411 -759 1469 -725
rect 1411 -793 1423 -759
rect 1457 -793 1469 -759
rect 1411 -827 1469 -793
rect 1411 -861 1423 -827
rect 1457 -861 1469 -827
rect 1411 -876 1469 -861
rect 1669 -691 1727 -676
rect 1669 -725 1681 -691
rect 1715 -725 1727 -691
rect 1669 -759 1727 -725
rect 1669 -793 1681 -759
rect 1715 -793 1727 -759
rect 1669 -827 1727 -793
rect 1669 -861 1681 -827
rect 1715 -861 1727 -827
rect 1669 -876 1727 -861
rect 1927 -691 1985 -676
rect 1927 -725 1939 -691
rect 1973 -725 1985 -691
rect 1927 -759 1985 -725
rect 1927 -793 1939 -759
rect 1973 -793 1985 -759
rect 1927 -827 1985 -793
rect 1927 -861 1939 -827
rect 1973 -861 1985 -827
rect 1927 -876 1985 -861
rect 2185 -691 2243 -676
rect 2185 -725 2197 -691
rect 2231 -725 2243 -691
rect 2185 -759 2243 -725
rect 2185 -793 2197 -759
rect 2231 -793 2243 -759
rect 2185 -827 2243 -793
rect 2185 -861 2197 -827
rect 2231 -861 2243 -827
rect 2185 -876 2243 -861
rect 2443 -691 2501 -676
rect 2443 -725 2455 -691
rect 2489 -725 2501 -691
rect 2443 -759 2501 -725
rect 2443 -793 2455 -759
rect 2489 -793 2501 -759
rect 2443 -827 2501 -793
rect 2443 -861 2455 -827
rect 2489 -861 2501 -827
rect 2443 -876 2501 -861
rect 2637 -691 2695 -676
rect 2637 -725 2649 -691
rect 2683 -725 2695 -691
rect 2637 -759 2695 -725
rect 2637 -793 2649 -759
rect 2683 -793 2695 -759
rect 2637 -827 2695 -793
rect 2637 -861 2649 -827
rect 2683 -861 2695 -827
rect 2637 -876 2695 -861
rect 2895 -691 2953 -676
rect 2895 -725 2907 -691
rect 2941 -725 2953 -691
rect 2895 -759 2953 -725
rect 2895 -793 2907 -759
rect 2941 -793 2953 -759
rect 2895 -827 2953 -793
rect 2895 -861 2907 -827
rect 2941 -861 2953 -827
rect 2895 -876 2953 -861
rect 3153 -691 3211 -676
rect 3153 -725 3165 -691
rect 3199 -725 3211 -691
rect 3153 -759 3211 -725
rect 3153 -793 3165 -759
rect 3199 -793 3211 -759
rect 3153 -827 3211 -793
rect 3153 -861 3165 -827
rect 3199 -861 3211 -827
rect 3153 -876 3211 -861
rect 3411 -691 3469 -676
rect 3411 -725 3423 -691
rect 3457 -725 3469 -691
rect 3411 -759 3469 -725
rect 3411 -793 3423 -759
rect 3457 -793 3469 -759
rect 3411 -827 3469 -793
rect 3411 -861 3423 -827
rect 3457 -861 3469 -827
rect 3411 -876 3469 -861
rect 3605 -691 3663 -676
rect 3605 -725 3617 -691
rect 3651 -725 3663 -691
rect 3605 -759 3663 -725
rect 3605 -793 3617 -759
rect 3651 -793 3663 -759
rect 3605 -827 3663 -793
rect 3605 -861 3617 -827
rect 3651 -861 3663 -827
rect 3605 -876 3663 -861
rect 3863 -691 3921 -676
rect 3863 -725 3875 -691
rect 3909 -725 3921 -691
rect 3863 -759 3921 -725
rect 3863 -793 3875 -759
rect 3909 -793 3921 -759
rect 3863 -827 3921 -793
rect 3863 -861 3875 -827
rect 3909 -861 3921 -827
rect 3863 -876 3921 -861
rect 4121 -691 4179 -676
rect 4121 -725 4133 -691
rect 4167 -725 4179 -691
rect 4121 -759 4179 -725
rect 4121 -793 4133 -759
rect 4167 -793 4179 -759
rect 4121 -827 4179 -793
rect 4121 -861 4133 -827
rect 4167 -861 4179 -827
rect 4121 -876 4179 -861
rect 4379 -691 4437 -676
rect 4379 -725 4391 -691
rect 4425 -725 4437 -691
rect 4379 -759 4437 -725
rect 4379 -793 4391 -759
rect 4425 -793 4437 -759
rect 4379 -827 4437 -793
rect 4379 -861 4391 -827
rect 4425 -861 4437 -827
rect 4379 -876 4437 -861
rect 4637 -691 4695 -676
rect 4637 -725 4649 -691
rect 4683 -725 4695 -691
rect 4637 -759 4695 -725
rect 4637 -793 4649 -759
rect 4683 -793 4695 -759
rect 4637 -827 4695 -793
rect 4637 -861 4649 -827
rect 4683 -861 4695 -827
rect 4637 -876 4695 -861
rect 4830 -691 4888 -676
rect 4830 -725 4842 -691
rect 4876 -725 4888 -691
rect 4830 -759 4888 -725
rect 4830 -793 4842 -759
rect 4876 -793 4888 -759
rect 4830 -827 4888 -793
rect 4830 -861 4842 -827
rect 4876 -861 4888 -827
rect 4830 -876 4888 -861
rect 5088 -691 5146 -676
rect 5088 -725 5100 -691
rect 5134 -725 5146 -691
rect 5088 -759 5146 -725
rect 5088 -793 5100 -759
rect 5134 -793 5146 -759
rect 5088 -827 5146 -793
rect 5088 -861 5100 -827
rect 5134 -861 5146 -827
rect 5088 -876 5146 -861
rect 5316 -691 5374 -676
rect 5316 -725 5328 -691
rect 5362 -725 5374 -691
rect 5316 -759 5374 -725
rect 5316 -793 5328 -759
rect 5362 -793 5374 -759
rect 5316 -827 5374 -793
rect 5316 -861 5328 -827
rect 5362 -861 5374 -827
rect 5316 -876 5374 -861
rect 5574 -691 5632 -676
rect 5574 -725 5586 -691
rect 5620 -725 5632 -691
rect 5574 -759 5632 -725
rect 5574 -793 5586 -759
rect 5620 -793 5632 -759
rect 5574 -827 5632 -793
rect 5574 -861 5586 -827
rect 5620 -861 5632 -827
rect 5574 -876 5632 -861
rect 5768 -691 5826 -676
rect 5768 -725 5780 -691
rect 5814 -725 5826 -691
rect 5768 -759 5826 -725
rect 5768 -793 5780 -759
rect 5814 -793 5826 -759
rect 5768 -827 5826 -793
rect 5768 -861 5780 -827
rect 5814 -861 5826 -827
rect 5768 -876 5826 -861
rect 6026 -691 6084 -676
rect 6026 -725 6038 -691
rect 6072 -725 6084 -691
rect 6026 -759 6084 -725
rect 6026 -793 6038 -759
rect 6072 -793 6084 -759
rect 6026 -827 6084 -793
rect 6026 -861 6038 -827
rect 6072 -861 6084 -827
rect 6026 -876 6084 -861
rect 6284 -691 6342 -676
rect 6284 -725 6296 -691
rect 6330 -725 6342 -691
rect 6284 -759 6342 -725
rect 6284 -793 6296 -759
rect 6330 -793 6342 -759
rect 6284 -827 6342 -793
rect 6284 -861 6296 -827
rect 6330 -861 6342 -827
rect 6284 -876 6342 -861
rect 6542 -691 6600 -676
rect 6542 -725 6554 -691
rect 6588 -725 6600 -691
rect 6542 -759 6600 -725
rect 6542 -793 6554 -759
rect 6588 -793 6600 -759
rect 6542 -827 6600 -793
rect 6542 -861 6554 -827
rect 6588 -861 6600 -827
rect 6542 -876 6600 -861
rect 6800 -691 6858 -676
rect 6800 -725 6812 -691
rect 6846 -725 6858 -691
rect 6800 -759 6858 -725
rect 6800 -793 6812 -759
rect 6846 -793 6858 -759
rect 6800 -827 6858 -793
rect 6800 -861 6812 -827
rect 6846 -861 6858 -827
rect 6800 -876 6858 -861
rect 6994 -691 7052 -676
rect 6994 -725 7006 -691
rect 7040 -725 7052 -691
rect 6994 -759 7052 -725
rect 6994 -793 7006 -759
rect 7040 -793 7052 -759
rect 6994 -827 7052 -793
rect 6994 -861 7006 -827
rect 7040 -861 7052 -827
rect 6994 -876 7052 -861
rect 7252 -691 7310 -676
rect 7252 -725 7264 -691
rect 7298 -725 7310 -691
rect 7252 -759 7310 -725
rect 7252 -793 7264 -759
rect 7298 -793 7310 -759
rect 7252 -827 7310 -793
rect 7252 -861 7264 -827
rect 7298 -861 7310 -827
rect 7252 -876 7310 -861
rect 7510 -691 7568 -676
rect 7510 -725 7522 -691
rect 7556 -725 7568 -691
rect 7510 -759 7568 -725
rect 7510 -793 7522 -759
rect 7556 -793 7568 -759
rect 7510 -827 7568 -793
rect 7510 -861 7522 -827
rect 7556 -861 7568 -827
rect 7510 -876 7568 -861
rect 7768 -691 7826 -676
rect 7768 -725 7780 -691
rect 7814 -725 7826 -691
rect 7768 -759 7826 -725
rect 7768 -793 7780 -759
rect 7814 -793 7826 -759
rect 7768 -827 7826 -793
rect 7768 -861 7780 -827
rect 7814 -861 7826 -827
rect 7768 -876 7826 -861
rect 7962 -691 8020 -676
rect 7962 -725 7974 -691
rect 8008 -725 8020 -691
rect 7962 -759 8020 -725
rect 7962 -793 7974 -759
rect 8008 -793 8020 -759
rect 7962 -827 8020 -793
rect 7962 -861 7974 -827
rect 8008 -861 8020 -827
rect 7962 -876 8020 -861
rect 8220 -691 8278 -676
rect 8220 -725 8232 -691
rect 8266 -725 8278 -691
rect 8220 -759 8278 -725
rect 8220 -793 8232 -759
rect 8266 -793 8278 -759
rect 8220 -827 8278 -793
rect 8220 -861 8232 -827
rect 8266 -861 8278 -827
rect 8220 -876 8278 -861
rect 8478 -691 8536 -676
rect 8478 -725 8490 -691
rect 8524 -725 8536 -691
rect 8478 -759 8536 -725
rect 8478 -793 8490 -759
rect 8524 -793 8536 -759
rect 8478 -827 8536 -793
rect 8478 -861 8490 -827
rect 8524 -861 8536 -827
rect 8478 -876 8536 -861
rect 8736 -691 8794 -676
rect 8736 -725 8748 -691
rect 8782 -725 8794 -691
rect 8736 -759 8794 -725
rect 8736 -793 8748 -759
rect 8782 -793 8794 -759
rect 8736 -827 8794 -793
rect 8736 -861 8748 -827
rect 8782 -861 8794 -827
rect 8736 -876 8794 -861
rect 8994 -691 9052 -676
rect 8994 -725 9006 -691
rect 9040 -725 9052 -691
rect 8994 -759 9052 -725
rect 8994 -793 9006 -759
rect 9040 -793 9052 -759
rect 8994 -827 9052 -793
rect 8994 -861 9006 -827
rect 9040 -861 9052 -827
rect 8994 -876 9052 -861
rect 9188 -691 9246 -676
rect 9188 -725 9200 -691
rect 9234 -725 9246 -691
rect 9188 -759 9246 -725
rect 9188 -793 9200 -759
rect 9234 -793 9246 -759
rect 9188 -827 9246 -793
rect 9188 -861 9200 -827
rect 9234 -861 9246 -827
rect 9188 -876 9246 -861
rect 9446 -691 9504 -676
rect 9446 -725 9458 -691
rect 9492 -725 9504 -691
rect 9446 -759 9504 -725
rect 9446 -793 9458 -759
rect 9492 -793 9504 -759
rect 9446 -827 9504 -793
rect 9446 -861 9458 -827
rect 9492 -861 9504 -827
rect 9446 -876 9504 -861
rect 9676 -691 9734 -676
rect 9676 -725 9688 -691
rect 9722 -725 9734 -691
rect 9676 -759 9734 -725
rect 9676 -793 9688 -759
rect 9722 -793 9734 -759
rect 9676 -827 9734 -793
rect 9676 -861 9688 -827
rect 9722 -861 9734 -827
rect 9676 -876 9734 -861
rect 9934 -691 9992 -676
rect 9934 -725 9946 -691
rect 9980 -725 9992 -691
rect 9934 -759 9992 -725
rect 9934 -793 9946 -759
rect 9980 -793 9992 -759
rect 9934 -827 9992 -793
rect 9934 -861 9946 -827
rect 9980 -861 9992 -827
rect 9934 -876 9992 -861
rect 10128 -691 10186 -676
rect 10128 -725 10140 -691
rect 10174 -725 10186 -691
rect 10128 -759 10186 -725
rect 10128 -793 10140 -759
rect 10174 -793 10186 -759
rect 10128 -827 10186 -793
rect 10128 -861 10140 -827
rect 10174 -861 10186 -827
rect 10128 -876 10186 -861
rect 10386 -691 10444 -676
rect 10386 -725 10398 -691
rect 10432 -725 10444 -691
rect 10386 -759 10444 -725
rect 10386 -793 10398 -759
rect 10432 -793 10444 -759
rect 10386 -827 10444 -793
rect 10386 -861 10398 -827
rect 10432 -861 10444 -827
rect 10386 -876 10444 -861
rect 10644 -691 10702 -676
rect 10644 -725 10656 -691
rect 10690 -725 10702 -691
rect 10644 -759 10702 -725
rect 10644 -793 10656 -759
rect 10690 -793 10702 -759
rect 10644 -827 10702 -793
rect 10644 -861 10656 -827
rect 10690 -861 10702 -827
rect 10644 -876 10702 -861
rect 10902 -691 10960 -676
rect 10902 -725 10914 -691
rect 10948 -725 10960 -691
rect 10902 -759 10960 -725
rect 10902 -793 10914 -759
rect 10948 -793 10960 -759
rect 10902 -827 10960 -793
rect 10902 -861 10914 -827
rect 10948 -861 10960 -827
rect 10902 -876 10960 -861
rect 11160 -691 11218 -676
rect 11160 -725 11172 -691
rect 11206 -725 11218 -691
rect 11160 -759 11218 -725
rect 11160 -793 11172 -759
rect 11206 -793 11218 -759
rect 11160 -827 11218 -793
rect 11160 -861 11172 -827
rect 11206 -861 11218 -827
rect 11160 -876 11218 -861
rect 11354 -691 11412 -676
rect 11354 -725 11366 -691
rect 11400 -725 11412 -691
rect 11354 -759 11412 -725
rect 11354 -793 11366 -759
rect 11400 -793 11412 -759
rect 11354 -827 11412 -793
rect 11354 -861 11366 -827
rect 11400 -861 11412 -827
rect 11354 -876 11412 -861
rect 11612 -691 11670 -676
rect 11612 -725 11624 -691
rect 11658 -725 11670 -691
rect 11612 -759 11670 -725
rect 11612 -793 11624 -759
rect 11658 -793 11670 -759
rect 11612 -827 11670 -793
rect 11612 -861 11624 -827
rect 11658 -861 11670 -827
rect 11612 -876 11670 -861
rect 11870 -691 11928 -676
rect 11870 -725 11882 -691
rect 11916 -725 11928 -691
rect 11870 -759 11928 -725
rect 11870 -793 11882 -759
rect 11916 -793 11928 -759
rect 11870 -827 11928 -793
rect 11870 -861 11882 -827
rect 11916 -861 11928 -827
rect 11870 -876 11928 -861
rect 12128 -691 12186 -676
rect 12128 -725 12140 -691
rect 12174 -725 12186 -691
rect 12128 -759 12186 -725
rect 12128 -793 12140 -759
rect 12174 -793 12186 -759
rect 12128 -827 12186 -793
rect 12128 -861 12140 -827
rect 12174 -861 12186 -827
rect 12128 -876 12186 -861
rect 12322 -691 12380 -676
rect 12322 -725 12334 -691
rect 12368 -725 12380 -691
rect 12322 -759 12380 -725
rect 12322 -793 12334 -759
rect 12368 -793 12380 -759
rect 12322 -827 12380 -793
rect 12322 -861 12334 -827
rect 12368 -861 12380 -827
rect 12322 -876 12380 -861
rect 12580 -691 12638 -676
rect 12580 -725 12592 -691
rect 12626 -725 12638 -691
rect 12580 -759 12638 -725
rect 12580 -793 12592 -759
rect 12626 -793 12638 -759
rect 12580 -827 12638 -793
rect 12580 -861 12592 -827
rect 12626 -861 12638 -827
rect 12580 -876 12638 -861
rect 12838 -691 12896 -676
rect 12838 -725 12850 -691
rect 12884 -725 12896 -691
rect 12838 -759 12896 -725
rect 12838 -793 12850 -759
rect 12884 -793 12896 -759
rect 12838 -827 12896 -793
rect 12838 -861 12850 -827
rect 12884 -861 12896 -827
rect 12838 -876 12896 -861
rect 13096 -691 13154 -676
rect 13096 -725 13108 -691
rect 13142 -725 13154 -691
rect 13096 -759 13154 -725
rect 13096 -793 13108 -759
rect 13142 -793 13154 -759
rect 13096 -827 13154 -793
rect 13096 -861 13108 -827
rect 13142 -861 13154 -827
rect 13096 -876 13154 -861
rect 13354 -691 13412 -676
rect 13354 -725 13366 -691
rect 13400 -725 13412 -691
rect 13354 -759 13412 -725
rect 13354 -793 13366 -759
rect 13400 -793 13412 -759
rect 13354 -827 13412 -793
rect 13354 -861 13366 -827
rect 13400 -861 13412 -827
rect 13354 -876 13412 -861
rect 13548 -691 13606 -676
rect 13548 -725 13560 -691
rect 13594 -725 13606 -691
rect 13548 -759 13606 -725
rect 13548 -793 13560 -759
rect 13594 -793 13606 -759
rect 13548 -827 13606 -793
rect 13548 -861 13560 -827
rect 13594 -861 13606 -827
rect 13548 -876 13606 -861
rect 13806 -691 13864 -676
rect 13806 -725 13818 -691
rect 13852 -725 13864 -691
rect 13806 -759 13864 -725
rect 13806 -793 13818 -759
rect 13852 -793 13864 -759
rect 13806 -827 13864 -793
rect 13806 -861 13818 -827
rect 13852 -861 13864 -827
rect 13806 -876 13864 -861
rect 14034 -691 14092 -676
rect 14034 -725 14046 -691
rect 14080 -725 14092 -691
rect 14034 -759 14092 -725
rect 14034 -793 14046 -759
rect 14080 -793 14092 -759
rect 14034 -827 14092 -793
rect 14034 -861 14046 -827
rect 14080 -861 14092 -827
rect 14034 -876 14092 -861
rect 14292 -691 14350 -676
rect 14292 -725 14304 -691
rect 14338 -725 14350 -691
rect 14292 -759 14350 -725
rect 14292 -793 14304 -759
rect 14338 -793 14350 -759
rect 14292 -827 14350 -793
rect 14292 -861 14304 -827
rect 14338 -861 14350 -827
rect 14292 -876 14350 -861
rect 14485 -691 14543 -676
rect 14485 -725 14497 -691
rect 14531 -725 14543 -691
rect 14485 -759 14543 -725
rect 14485 -793 14497 -759
rect 14531 -793 14543 -759
rect 14485 -827 14543 -793
rect 14485 -861 14497 -827
rect 14531 -861 14543 -827
rect 14485 -876 14543 -861
rect 14743 -691 14801 -676
rect 14743 -725 14755 -691
rect 14789 -725 14801 -691
rect 14743 -759 14801 -725
rect 14743 -793 14755 -759
rect 14789 -793 14801 -759
rect 14743 -827 14801 -793
rect 14743 -861 14755 -827
rect 14789 -861 14801 -827
rect 14743 -876 14801 -861
rect 15001 -691 15059 -676
rect 15001 -725 15013 -691
rect 15047 -725 15059 -691
rect 15001 -759 15059 -725
rect 15001 -793 15013 -759
rect 15047 -793 15059 -759
rect 15001 -827 15059 -793
rect 15001 -861 15013 -827
rect 15047 -861 15059 -827
rect 15001 -876 15059 -861
rect 15259 -691 15317 -676
rect 15259 -725 15271 -691
rect 15305 -725 15317 -691
rect 15259 -759 15317 -725
rect 15259 -793 15271 -759
rect 15305 -793 15317 -759
rect 15259 -827 15317 -793
rect 15259 -861 15271 -827
rect 15305 -861 15317 -827
rect 15259 -876 15317 -861
rect 15517 -691 15575 -676
rect 15517 -725 15529 -691
rect 15563 -725 15575 -691
rect 15517 -759 15575 -725
rect 15517 -793 15529 -759
rect 15563 -793 15575 -759
rect 15517 -827 15575 -793
rect 15517 -861 15529 -827
rect 15563 -861 15575 -827
rect 15517 -876 15575 -861
rect 15711 -691 15769 -676
rect 15711 -725 15723 -691
rect 15757 -725 15769 -691
rect 15711 -759 15769 -725
rect 15711 -793 15723 -759
rect 15757 -793 15769 -759
rect 15711 -827 15769 -793
rect 15711 -861 15723 -827
rect 15757 -861 15769 -827
rect 15711 -876 15769 -861
rect 15969 -691 16027 -676
rect 15969 -725 15981 -691
rect 16015 -725 16027 -691
rect 15969 -759 16027 -725
rect 15969 -793 15981 -759
rect 16015 -793 16027 -759
rect 15969 -827 16027 -793
rect 15969 -861 15981 -827
rect 16015 -861 16027 -827
rect 15969 -876 16027 -861
rect 16227 -691 16285 -676
rect 16227 -725 16239 -691
rect 16273 -725 16285 -691
rect 16227 -759 16285 -725
rect 16227 -793 16239 -759
rect 16273 -793 16285 -759
rect 16227 -827 16285 -793
rect 16227 -861 16239 -827
rect 16273 -861 16285 -827
rect 16227 -876 16285 -861
rect 16485 -691 16543 -676
rect 16485 -725 16497 -691
rect 16531 -725 16543 -691
rect 16485 -759 16543 -725
rect 16485 -793 16497 -759
rect 16531 -793 16543 -759
rect 16485 -827 16543 -793
rect 16485 -861 16497 -827
rect 16531 -861 16543 -827
rect 16485 -876 16543 -861
rect 16679 -691 16737 -676
rect 16679 -725 16691 -691
rect 16725 -725 16737 -691
rect 16679 -759 16737 -725
rect 16679 -793 16691 -759
rect 16725 -793 16737 -759
rect 16679 -827 16737 -793
rect 16679 -861 16691 -827
rect 16725 -861 16737 -827
rect 16679 -876 16737 -861
rect 16937 -691 16995 -676
rect 16937 -725 16949 -691
rect 16983 -725 16995 -691
rect 16937 -759 16995 -725
rect 16937 -793 16949 -759
rect 16983 -793 16995 -759
rect 16937 -827 16995 -793
rect 16937 -861 16949 -827
rect 16983 -861 16995 -827
rect 16937 -876 16995 -861
rect 17195 -691 17253 -676
rect 17195 -725 17207 -691
rect 17241 -725 17253 -691
rect 17195 -759 17253 -725
rect 17195 -793 17207 -759
rect 17241 -793 17253 -759
rect 17195 -827 17253 -793
rect 17195 -861 17207 -827
rect 17241 -861 17253 -827
rect 17195 -876 17253 -861
rect 17453 -691 17511 -676
rect 17453 -725 17465 -691
rect 17499 -725 17511 -691
rect 17453 -759 17511 -725
rect 17453 -793 17465 -759
rect 17499 -793 17511 -759
rect 17453 -827 17511 -793
rect 17453 -861 17465 -827
rect 17499 -861 17511 -827
rect 17453 -876 17511 -861
rect 17711 -691 17769 -676
rect 17711 -725 17723 -691
rect 17757 -725 17769 -691
rect 17711 -759 17769 -725
rect 17711 -793 17723 -759
rect 17757 -793 17769 -759
rect 17711 -827 17769 -793
rect 17711 -861 17723 -827
rect 17757 -861 17769 -827
rect 17711 -876 17769 -861
rect 17905 -691 17963 -676
rect 17905 -725 17917 -691
rect 17951 -725 17963 -691
rect 17905 -759 17963 -725
rect 17905 -793 17917 -759
rect 17951 -793 17963 -759
rect 17905 -827 17963 -793
rect 17905 -861 17917 -827
rect 17951 -861 17963 -827
rect 17905 -876 17963 -861
rect 18163 -691 18221 -676
rect 18163 -725 18175 -691
rect 18209 -725 18221 -691
rect 18163 -759 18221 -725
rect 18163 -793 18175 -759
rect 18209 -793 18221 -759
rect 18163 -827 18221 -793
rect 18163 -861 18175 -827
rect 18209 -861 18221 -827
rect 18163 -876 18221 -861
rect 959 -1382 1017 -1367
rect 959 -1416 971 -1382
rect 1005 -1416 1017 -1382
rect 959 -1450 1017 -1416
rect 959 -1484 971 -1450
rect 1005 -1484 1017 -1450
rect 959 -1518 1017 -1484
rect 959 -1552 971 -1518
rect 1005 -1552 1017 -1518
rect 959 -1567 1017 -1552
rect 1217 -1382 1275 -1367
rect 1217 -1416 1229 -1382
rect 1263 -1416 1275 -1382
rect 1217 -1450 1275 -1416
rect 1217 -1484 1229 -1450
rect 1263 -1484 1275 -1450
rect 1217 -1518 1275 -1484
rect 1217 -1552 1229 -1518
rect 1263 -1552 1275 -1518
rect 1217 -1567 1275 -1552
rect 1411 -1382 1469 -1367
rect 1411 -1416 1423 -1382
rect 1457 -1416 1469 -1382
rect 1411 -1450 1469 -1416
rect 1411 -1484 1423 -1450
rect 1457 -1484 1469 -1450
rect 1411 -1518 1469 -1484
rect 1411 -1552 1423 -1518
rect 1457 -1552 1469 -1518
rect 1411 -1567 1469 -1552
rect 1669 -1382 1727 -1367
rect 1669 -1416 1681 -1382
rect 1715 -1416 1727 -1382
rect 1669 -1450 1727 -1416
rect 1669 -1484 1681 -1450
rect 1715 -1484 1727 -1450
rect 1669 -1518 1727 -1484
rect 1669 -1552 1681 -1518
rect 1715 -1552 1727 -1518
rect 1669 -1567 1727 -1552
rect 1927 -1382 1985 -1367
rect 1927 -1416 1939 -1382
rect 1973 -1416 1985 -1382
rect 1927 -1450 1985 -1416
rect 1927 -1484 1939 -1450
rect 1973 -1484 1985 -1450
rect 1927 -1518 1985 -1484
rect 1927 -1552 1939 -1518
rect 1973 -1552 1985 -1518
rect 1927 -1567 1985 -1552
rect 2185 -1382 2243 -1367
rect 2185 -1416 2197 -1382
rect 2231 -1416 2243 -1382
rect 2185 -1450 2243 -1416
rect 2185 -1484 2197 -1450
rect 2231 -1484 2243 -1450
rect 2185 -1518 2243 -1484
rect 2185 -1552 2197 -1518
rect 2231 -1552 2243 -1518
rect 2185 -1567 2243 -1552
rect 2443 -1382 2501 -1367
rect 2443 -1416 2455 -1382
rect 2489 -1416 2501 -1382
rect 2443 -1450 2501 -1416
rect 2443 -1484 2455 -1450
rect 2489 -1484 2501 -1450
rect 2443 -1518 2501 -1484
rect 2443 -1552 2455 -1518
rect 2489 -1552 2501 -1518
rect 2443 -1567 2501 -1552
rect 2637 -1382 2695 -1367
rect 2637 -1416 2649 -1382
rect 2683 -1416 2695 -1382
rect 2637 -1450 2695 -1416
rect 2637 -1484 2649 -1450
rect 2683 -1484 2695 -1450
rect 2637 -1518 2695 -1484
rect 2637 -1552 2649 -1518
rect 2683 -1552 2695 -1518
rect 2637 -1567 2695 -1552
rect 2895 -1382 2953 -1367
rect 2895 -1416 2907 -1382
rect 2941 -1416 2953 -1382
rect 2895 -1450 2953 -1416
rect 2895 -1484 2907 -1450
rect 2941 -1484 2953 -1450
rect 2895 -1518 2953 -1484
rect 2895 -1552 2907 -1518
rect 2941 -1552 2953 -1518
rect 2895 -1567 2953 -1552
rect 3153 -1382 3211 -1367
rect 3153 -1416 3165 -1382
rect 3199 -1416 3211 -1382
rect 3153 -1450 3211 -1416
rect 3153 -1484 3165 -1450
rect 3199 -1484 3211 -1450
rect 3153 -1518 3211 -1484
rect 3153 -1552 3165 -1518
rect 3199 -1552 3211 -1518
rect 3153 -1567 3211 -1552
rect 3411 -1382 3469 -1367
rect 3411 -1416 3423 -1382
rect 3457 -1416 3469 -1382
rect 3411 -1450 3469 -1416
rect 3411 -1484 3423 -1450
rect 3457 -1484 3469 -1450
rect 3411 -1518 3469 -1484
rect 3411 -1552 3423 -1518
rect 3457 -1552 3469 -1518
rect 3411 -1567 3469 -1552
rect 3605 -1382 3663 -1367
rect 3605 -1416 3617 -1382
rect 3651 -1416 3663 -1382
rect 3605 -1450 3663 -1416
rect 3605 -1484 3617 -1450
rect 3651 -1484 3663 -1450
rect 3605 -1518 3663 -1484
rect 3605 -1552 3617 -1518
rect 3651 -1552 3663 -1518
rect 3605 -1567 3663 -1552
rect 3863 -1382 3921 -1367
rect 3863 -1416 3875 -1382
rect 3909 -1416 3921 -1382
rect 3863 -1450 3921 -1416
rect 3863 -1484 3875 -1450
rect 3909 -1484 3921 -1450
rect 3863 -1518 3921 -1484
rect 3863 -1552 3875 -1518
rect 3909 -1552 3921 -1518
rect 3863 -1567 3921 -1552
rect 4121 -1382 4179 -1367
rect 4121 -1416 4133 -1382
rect 4167 -1416 4179 -1382
rect 4121 -1450 4179 -1416
rect 4121 -1484 4133 -1450
rect 4167 -1484 4179 -1450
rect 4121 -1518 4179 -1484
rect 4121 -1552 4133 -1518
rect 4167 -1552 4179 -1518
rect 4121 -1567 4179 -1552
rect 4379 -1382 4437 -1367
rect 4379 -1416 4391 -1382
rect 4425 -1416 4437 -1382
rect 4379 -1450 4437 -1416
rect 4379 -1484 4391 -1450
rect 4425 -1484 4437 -1450
rect 4379 -1518 4437 -1484
rect 4379 -1552 4391 -1518
rect 4425 -1552 4437 -1518
rect 4379 -1567 4437 -1552
rect 4637 -1382 4695 -1367
rect 4637 -1416 4649 -1382
rect 4683 -1416 4695 -1382
rect 4637 -1450 4695 -1416
rect 4637 -1484 4649 -1450
rect 4683 -1484 4695 -1450
rect 4637 -1518 4695 -1484
rect 4637 -1552 4649 -1518
rect 4683 -1552 4695 -1518
rect 4637 -1567 4695 -1552
rect 4830 -1382 4888 -1367
rect 4830 -1416 4842 -1382
rect 4876 -1416 4888 -1382
rect 4830 -1450 4888 -1416
rect 4830 -1484 4842 -1450
rect 4876 -1484 4888 -1450
rect 4830 -1518 4888 -1484
rect 4830 -1552 4842 -1518
rect 4876 -1552 4888 -1518
rect 4830 -1567 4888 -1552
rect 5088 -1382 5146 -1367
rect 5088 -1416 5100 -1382
rect 5134 -1416 5146 -1382
rect 5088 -1450 5146 -1416
rect 5088 -1484 5100 -1450
rect 5134 -1484 5146 -1450
rect 5088 -1518 5146 -1484
rect 5088 -1552 5100 -1518
rect 5134 -1552 5146 -1518
rect 5088 -1567 5146 -1552
rect 5316 -1382 5374 -1367
rect 5316 -1416 5328 -1382
rect 5362 -1416 5374 -1382
rect 5316 -1450 5374 -1416
rect 5316 -1484 5328 -1450
rect 5362 -1484 5374 -1450
rect 5316 -1518 5374 -1484
rect 5316 -1552 5328 -1518
rect 5362 -1552 5374 -1518
rect 5316 -1567 5374 -1552
rect 5574 -1382 5632 -1367
rect 5574 -1416 5586 -1382
rect 5620 -1416 5632 -1382
rect 5574 -1450 5632 -1416
rect 5574 -1484 5586 -1450
rect 5620 -1484 5632 -1450
rect 5574 -1518 5632 -1484
rect 5574 -1552 5586 -1518
rect 5620 -1552 5632 -1518
rect 5574 -1567 5632 -1552
rect 5768 -1382 5826 -1367
rect 5768 -1416 5780 -1382
rect 5814 -1416 5826 -1382
rect 5768 -1450 5826 -1416
rect 5768 -1484 5780 -1450
rect 5814 -1484 5826 -1450
rect 5768 -1518 5826 -1484
rect 5768 -1552 5780 -1518
rect 5814 -1552 5826 -1518
rect 5768 -1567 5826 -1552
rect 6026 -1382 6084 -1367
rect 6026 -1416 6038 -1382
rect 6072 -1416 6084 -1382
rect 6026 -1450 6084 -1416
rect 6026 -1484 6038 -1450
rect 6072 -1484 6084 -1450
rect 6026 -1518 6084 -1484
rect 6026 -1552 6038 -1518
rect 6072 -1552 6084 -1518
rect 6026 -1567 6084 -1552
rect 6284 -1382 6342 -1367
rect 6284 -1416 6296 -1382
rect 6330 -1416 6342 -1382
rect 6284 -1450 6342 -1416
rect 6284 -1484 6296 -1450
rect 6330 -1484 6342 -1450
rect 6284 -1518 6342 -1484
rect 6284 -1552 6296 -1518
rect 6330 -1552 6342 -1518
rect 6284 -1567 6342 -1552
rect 6542 -1382 6600 -1367
rect 6542 -1416 6554 -1382
rect 6588 -1416 6600 -1382
rect 6542 -1450 6600 -1416
rect 6542 -1484 6554 -1450
rect 6588 -1484 6600 -1450
rect 6542 -1518 6600 -1484
rect 6542 -1552 6554 -1518
rect 6588 -1552 6600 -1518
rect 6542 -1567 6600 -1552
rect 6800 -1382 6858 -1367
rect 6800 -1416 6812 -1382
rect 6846 -1416 6858 -1382
rect 6800 -1450 6858 -1416
rect 6800 -1484 6812 -1450
rect 6846 -1484 6858 -1450
rect 6800 -1518 6858 -1484
rect 6800 -1552 6812 -1518
rect 6846 -1552 6858 -1518
rect 6800 -1567 6858 -1552
rect 6994 -1382 7052 -1367
rect 6994 -1416 7006 -1382
rect 7040 -1416 7052 -1382
rect 6994 -1450 7052 -1416
rect 6994 -1484 7006 -1450
rect 7040 -1484 7052 -1450
rect 6994 -1518 7052 -1484
rect 6994 -1552 7006 -1518
rect 7040 -1552 7052 -1518
rect 6994 -1567 7052 -1552
rect 7252 -1382 7310 -1367
rect 7252 -1416 7264 -1382
rect 7298 -1416 7310 -1382
rect 7252 -1450 7310 -1416
rect 7252 -1484 7264 -1450
rect 7298 -1484 7310 -1450
rect 7252 -1518 7310 -1484
rect 7252 -1552 7264 -1518
rect 7298 -1552 7310 -1518
rect 7252 -1567 7310 -1552
rect 7510 -1382 7568 -1367
rect 7510 -1416 7522 -1382
rect 7556 -1416 7568 -1382
rect 7510 -1450 7568 -1416
rect 7510 -1484 7522 -1450
rect 7556 -1484 7568 -1450
rect 7510 -1518 7568 -1484
rect 7510 -1552 7522 -1518
rect 7556 -1552 7568 -1518
rect 7510 -1567 7568 -1552
rect 7768 -1382 7826 -1367
rect 7768 -1416 7780 -1382
rect 7814 -1416 7826 -1382
rect 7768 -1450 7826 -1416
rect 7768 -1484 7780 -1450
rect 7814 -1484 7826 -1450
rect 7768 -1518 7826 -1484
rect 7768 -1552 7780 -1518
rect 7814 -1552 7826 -1518
rect 7768 -1567 7826 -1552
rect 7962 -1382 8020 -1367
rect 7962 -1416 7974 -1382
rect 8008 -1416 8020 -1382
rect 7962 -1450 8020 -1416
rect 7962 -1484 7974 -1450
rect 8008 -1484 8020 -1450
rect 7962 -1518 8020 -1484
rect 7962 -1552 7974 -1518
rect 8008 -1552 8020 -1518
rect 7962 -1567 8020 -1552
rect 8220 -1382 8278 -1367
rect 8220 -1416 8232 -1382
rect 8266 -1416 8278 -1382
rect 8220 -1450 8278 -1416
rect 8220 -1484 8232 -1450
rect 8266 -1484 8278 -1450
rect 8220 -1518 8278 -1484
rect 8220 -1552 8232 -1518
rect 8266 -1552 8278 -1518
rect 8220 -1567 8278 -1552
rect 8478 -1382 8536 -1367
rect 8478 -1416 8490 -1382
rect 8524 -1416 8536 -1382
rect 8478 -1450 8536 -1416
rect 8478 -1484 8490 -1450
rect 8524 -1484 8536 -1450
rect 8478 -1518 8536 -1484
rect 8478 -1552 8490 -1518
rect 8524 -1552 8536 -1518
rect 8478 -1567 8536 -1552
rect 8736 -1382 8794 -1367
rect 8736 -1416 8748 -1382
rect 8782 -1416 8794 -1382
rect 8736 -1450 8794 -1416
rect 8736 -1484 8748 -1450
rect 8782 -1484 8794 -1450
rect 8736 -1518 8794 -1484
rect 8736 -1552 8748 -1518
rect 8782 -1552 8794 -1518
rect 8736 -1567 8794 -1552
rect 8994 -1382 9052 -1367
rect 8994 -1416 9006 -1382
rect 9040 -1416 9052 -1382
rect 8994 -1450 9052 -1416
rect 8994 -1484 9006 -1450
rect 9040 -1484 9052 -1450
rect 8994 -1518 9052 -1484
rect 8994 -1552 9006 -1518
rect 9040 -1552 9052 -1518
rect 8994 -1567 9052 -1552
rect 9188 -1382 9246 -1367
rect 9188 -1416 9200 -1382
rect 9234 -1416 9246 -1382
rect 9188 -1450 9246 -1416
rect 9188 -1484 9200 -1450
rect 9234 -1484 9246 -1450
rect 9188 -1518 9246 -1484
rect 9188 -1552 9200 -1518
rect 9234 -1552 9246 -1518
rect 9188 -1567 9246 -1552
rect 9446 -1382 9504 -1367
rect 9446 -1416 9458 -1382
rect 9492 -1416 9504 -1382
rect 9446 -1450 9504 -1416
rect 9446 -1484 9458 -1450
rect 9492 -1484 9504 -1450
rect 9446 -1518 9504 -1484
rect 9446 -1552 9458 -1518
rect 9492 -1552 9504 -1518
rect 9446 -1567 9504 -1552
rect 9676 -1382 9734 -1367
rect 9676 -1416 9688 -1382
rect 9722 -1416 9734 -1382
rect 9676 -1450 9734 -1416
rect 9676 -1484 9688 -1450
rect 9722 -1484 9734 -1450
rect 9676 -1518 9734 -1484
rect 9676 -1552 9688 -1518
rect 9722 -1552 9734 -1518
rect 9676 -1567 9734 -1552
rect 9934 -1382 9992 -1367
rect 9934 -1416 9946 -1382
rect 9980 -1416 9992 -1382
rect 9934 -1450 9992 -1416
rect 9934 -1484 9946 -1450
rect 9980 -1484 9992 -1450
rect 9934 -1518 9992 -1484
rect 9934 -1552 9946 -1518
rect 9980 -1552 9992 -1518
rect 9934 -1567 9992 -1552
rect 10128 -1382 10186 -1367
rect 10128 -1416 10140 -1382
rect 10174 -1416 10186 -1382
rect 10128 -1450 10186 -1416
rect 10128 -1484 10140 -1450
rect 10174 -1484 10186 -1450
rect 10128 -1518 10186 -1484
rect 10128 -1552 10140 -1518
rect 10174 -1552 10186 -1518
rect 10128 -1567 10186 -1552
rect 10386 -1382 10444 -1367
rect 10386 -1416 10398 -1382
rect 10432 -1416 10444 -1382
rect 10386 -1450 10444 -1416
rect 10386 -1484 10398 -1450
rect 10432 -1484 10444 -1450
rect 10386 -1518 10444 -1484
rect 10386 -1552 10398 -1518
rect 10432 -1552 10444 -1518
rect 10386 -1567 10444 -1552
rect 10644 -1382 10702 -1367
rect 10644 -1416 10656 -1382
rect 10690 -1416 10702 -1382
rect 10644 -1450 10702 -1416
rect 10644 -1484 10656 -1450
rect 10690 -1484 10702 -1450
rect 10644 -1518 10702 -1484
rect 10644 -1552 10656 -1518
rect 10690 -1552 10702 -1518
rect 10644 -1567 10702 -1552
rect 10902 -1382 10960 -1367
rect 10902 -1416 10914 -1382
rect 10948 -1416 10960 -1382
rect 10902 -1450 10960 -1416
rect 10902 -1484 10914 -1450
rect 10948 -1484 10960 -1450
rect 10902 -1518 10960 -1484
rect 10902 -1552 10914 -1518
rect 10948 -1552 10960 -1518
rect 10902 -1567 10960 -1552
rect 11160 -1382 11218 -1367
rect 11160 -1416 11172 -1382
rect 11206 -1416 11218 -1382
rect 11160 -1450 11218 -1416
rect 11160 -1484 11172 -1450
rect 11206 -1484 11218 -1450
rect 11160 -1518 11218 -1484
rect 11160 -1552 11172 -1518
rect 11206 -1552 11218 -1518
rect 11160 -1567 11218 -1552
rect 11354 -1382 11412 -1367
rect 11354 -1416 11366 -1382
rect 11400 -1416 11412 -1382
rect 11354 -1450 11412 -1416
rect 11354 -1484 11366 -1450
rect 11400 -1484 11412 -1450
rect 11354 -1518 11412 -1484
rect 11354 -1552 11366 -1518
rect 11400 -1552 11412 -1518
rect 11354 -1567 11412 -1552
rect 11612 -1382 11670 -1367
rect 11612 -1416 11624 -1382
rect 11658 -1416 11670 -1382
rect 11612 -1450 11670 -1416
rect 11612 -1484 11624 -1450
rect 11658 -1484 11670 -1450
rect 11612 -1518 11670 -1484
rect 11612 -1552 11624 -1518
rect 11658 -1552 11670 -1518
rect 11612 -1567 11670 -1552
rect 11870 -1382 11928 -1367
rect 11870 -1416 11882 -1382
rect 11916 -1416 11928 -1382
rect 11870 -1450 11928 -1416
rect 11870 -1484 11882 -1450
rect 11916 -1484 11928 -1450
rect 11870 -1518 11928 -1484
rect 11870 -1552 11882 -1518
rect 11916 -1552 11928 -1518
rect 11870 -1567 11928 -1552
rect 12128 -1382 12186 -1367
rect 12128 -1416 12140 -1382
rect 12174 -1416 12186 -1382
rect 12128 -1450 12186 -1416
rect 12128 -1484 12140 -1450
rect 12174 -1484 12186 -1450
rect 12128 -1518 12186 -1484
rect 12128 -1552 12140 -1518
rect 12174 -1552 12186 -1518
rect 12128 -1567 12186 -1552
rect 12322 -1382 12380 -1367
rect 12322 -1416 12334 -1382
rect 12368 -1416 12380 -1382
rect 12322 -1450 12380 -1416
rect 12322 -1484 12334 -1450
rect 12368 -1484 12380 -1450
rect 12322 -1518 12380 -1484
rect 12322 -1552 12334 -1518
rect 12368 -1552 12380 -1518
rect 12322 -1567 12380 -1552
rect 12580 -1382 12638 -1367
rect 12580 -1416 12592 -1382
rect 12626 -1416 12638 -1382
rect 12580 -1450 12638 -1416
rect 12580 -1484 12592 -1450
rect 12626 -1484 12638 -1450
rect 12580 -1518 12638 -1484
rect 12580 -1552 12592 -1518
rect 12626 -1552 12638 -1518
rect 12580 -1567 12638 -1552
rect 12838 -1382 12896 -1367
rect 12838 -1416 12850 -1382
rect 12884 -1416 12896 -1382
rect 12838 -1450 12896 -1416
rect 12838 -1484 12850 -1450
rect 12884 -1484 12896 -1450
rect 12838 -1518 12896 -1484
rect 12838 -1552 12850 -1518
rect 12884 -1552 12896 -1518
rect 12838 -1567 12896 -1552
rect 13096 -1382 13154 -1367
rect 13096 -1416 13108 -1382
rect 13142 -1416 13154 -1382
rect 13096 -1450 13154 -1416
rect 13096 -1484 13108 -1450
rect 13142 -1484 13154 -1450
rect 13096 -1518 13154 -1484
rect 13096 -1552 13108 -1518
rect 13142 -1552 13154 -1518
rect 13096 -1567 13154 -1552
rect 13354 -1382 13412 -1367
rect 13354 -1416 13366 -1382
rect 13400 -1416 13412 -1382
rect 13354 -1450 13412 -1416
rect 13354 -1484 13366 -1450
rect 13400 -1484 13412 -1450
rect 13354 -1518 13412 -1484
rect 13354 -1552 13366 -1518
rect 13400 -1552 13412 -1518
rect 13354 -1567 13412 -1552
rect 13548 -1382 13606 -1367
rect 13548 -1416 13560 -1382
rect 13594 -1416 13606 -1382
rect 13548 -1450 13606 -1416
rect 13548 -1484 13560 -1450
rect 13594 -1484 13606 -1450
rect 13548 -1518 13606 -1484
rect 13548 -1552 13560 -1518
rect 13594 -1552 13606 -1518
rect 13548 -1567 13606 -1552
rect 13806 -1382 13864 -1367
rect 13806 -1416 13818 -1382
rect 13852 -1416 13864 -1382
rect 13806 -1450 13864 -1416
rect 13806 -1484 13818 -1450
rect 13852 -1484 13864 -1450
rect 13806 -1518 13864 -1484
rect 13806 -1552 13818 -1518
rect 13852 -1552 13864 -1518
rect 13806 -1567 13864 -1552
rect 14034 -1382 14092 -1367
rect 14034 -1416 14046 -1382
rect 14080 -1416 14092 -1382
rect 14034 -1450 14092 -1416
rect 14034 -1484 14046 -1450
rect 14080 -1484 14092 -1450
rect 14034 -1518 14092 -1484
rect 14034 -1552 14046 -1518
rect 14080 -1552 14092 -1518
rect 14034 -1567 14092 -1552
rect 14292 -1382 14350 -1367
rect 14292 -1416 14304 -1382
rect 14338 -1416 14350 -1382
rect 14292 -1450 14350 -1416
rect 14292 -1484 14304 -1450
rect 14338 -1484 14350 -1450
rect 14292 -1518 14350 -1484
rect 14292 -1552 14304 -1518
rect 14338 -1552 14350 -1518
rect 14292 -1567 14350 -1552
rect 14485 -1382 14543 -1367
rect 14485 -1416 14497 -1382
rect 14531 -1416 14543 -1382
rect 14485 -1450 14543 -1416
rect 14485 -1484 14497 -1450
rect 14531 -1484 14543 -1450
rect 14485 -1518 14543 -1484
rect 14485 -1552 14497 -1518
rect 14531 -1552 14543 -1518
rect 14485 -1567 14543 -1552
rect 14743 -1382 14801 -1367
rect 14743 -1416 14755 -1382
rect 14789 -1416 14801 -1382
rect 14743 -1450 14801 -1416
rect 14743 -1484 14755 -1450
rect 14789 -1484 14801 -1450
rect 14743 -1518 14801 -1484
rect 14743 -1552 14755 -1518
rect 14789 -1552 14801 -1518
rect 14743 -1567 14801 -1552
rect 15001 -1382 15059 -1367
rect 15001 -1416 15013 -1382
rect 15047 -1416 15059 -1382
rect 15001 -1450 15059 -1416
rect 15001 -1484 15013 -1450
rect 15047 -1484 15059 -1450
rect 15001 -1518 15059 -1484
rect 15001 -1552 15013 -1518
rect 15047 -1552 15059 -1518
rect 15001 -1567 15059 -1552
rect 15259 -1382 15317 -1367
rect 15259 -1416 15271 -1382
rect 15305 -1416 15317 -1382
rect 15259 -1450 15317 -1416
rect 15259 -1484 15271 -1450
rect 15305 -1484 15317 -1450
rect 15259 -1518 15317 -1484
rect 15259 -1552 15271 -1518
rect 15305 -1552 15317 -1518
rect 15259 -1567 15317 -1552
rect 15517 -1382 15575 -1367
rect 15517 -1416 15529 -1382
rect 15563 -1416 15575 -1382
rect 15517 -1450 15575 -1416
rect 15517 -1484 15529 -1450
rect 15563 -1484 15575 -1450
rect 15517 -1518 15575 -1484
rect 15517 -1552 15529 -1518
rect 15563 -1552 15575 -1518
rect 15517 -1567 15575 -1552
rect 15711 -1382 15769 -1367
rect 15711 -1416 15723 -1382
rect 15757 -1416 15769 -1382
rect 15711 -1450 15769 -1416
rect 15711 -1484 15723 -1450
rect 15757 -1484 15769 -1450
rect 15711 -1518 15769 -1484
rect 15711 -1552 15723 -1518
rect 15757 -1552 15769 -1518
rect 15711 -1567 15769 -1552
rect 15969 -1382 16027 -1367
rect 15969 -1416 15981 -1382
rect 16015 -1416 16027 -1382
rect 15969 -1450 16027 -1416
rect 15969 -1484 15981 -1450
rect 16015 -1484 16027 -1450
rect 15969 -1518 16027 -1484
rect 15969 -1552 15981 -1518
rect 16015 -1552 16027 -1518
rect 15969 -1567 16027 -1552
rect 16227 -1382 16285 -1367
rect 16227 -1416 16239 -1382
rect 16273 -1416 16285 -1382
rect 16227 -1450 16285 -1416
rect 16227 -1484 16239 -1450
rect 16273 -1484 16285 -1450
rect 16227 -1518 16285 -1484
rect 16227 -1552 16239 -1518
rect 16273 -1552 16285 -1518
rect 16227 -1567 16285 -1552
rect 16485 -1382 16543 -1367
rect 16485 -1416 16497 -1382
rect 16531 -1416 16543 -1382
rect 16485 -1450 16543 -1416
rect 16485 -1484 16497 -1450
rect 16531 -1484 16543 -1450
rect 16485 -1518 16543 -1484
rect 16485 -1552 16497 -1518
rect 16531 -1552 16543 -1518
rect 16485 -1567 16543 -1552
rect 16679 -1382 16737 -1367
rect 16679 -1416 16691 -1382
rect 16725 -1416 16737 -1382
rect 16679 -1450 16737 -1416
rect 16679 -1484 16691 -1450
rect 16725 -1484 16737 -1450
rect 16679 -1518 16737 -1484
rect 16679 -1552 16691 -1518
rect 16725 -1552 16737 -1518
rect 16679 -1567 16737 -1552
rect 16937 -1382 16995 -1367
rect 16937 -1416 16949 -1382
rect 16983 -1416 16995 -1382
rect 16937 -1450 16995 -1416
rect 16937 -1484 16949 -1450
rect 16983 -1484 16995 -1450
rect 16937 -1518 16995 -1484
rect 16937 -1552 16949 -1518
rect 16983 -1552 16995 -1518
rect 16937 -1567 16995 -1552
rect 17195 -1382 17253 -1367
rect 17195 -1416 17207 -1382
rect 17241 -1416 17253 -1382
rect 17195 -1450 17253 -1416
rect 17195 -1484 17207 -1450
rect 17241 -1484 17253 -1450
rect 17195 -1518 17253 -1484
rect 17195 -1552 17207 -1518
rect 17241 -1552 17253 -1518
rect 17195 -1567 17253 -1552
rect 17453 -1382 17511 -1367
rect 17453 -1416 17465 -1382
rect 17499 -1416 17511 -1382
rect 17453 -1450 17511 -1416
rect 17453 -1484 17465 -1450
rect 17499 -1484 17511 -1450
rect 17453 -1518 17511 -1484
rect 17453 -1552 17465 -1518
rect 17499 -1552 17511 -1518
rect 17453 -1567 17511 -1552
rect 17711 -1382 17769 -1367
rect 17711 -1416 17723 -1382
rect 17757 -1416 17769 -1382
rect 17711 -1450 17769 -1416
rect 17711 -1484 17723 -1450
rect 17757 -1484 17769 -1450
rect 17711 -1518 17769 -1484
rect 17711 -1552 17723 -1518
rect 17757 -1552 17769 -1518
rect 17711 -1567 17769 -1552
rect 17905 -1382 17963 -1367
rect 17905 -1416 17917 -1382
rect 17951 -1416 17963 -1382
rect 17905 -1450 17963 -1416
rect 17905 -1484 17917 -1450
rect 17951 -1484 17963 -1450
rect 17905 -1518 17963 -1484
rect 17905 -1552 17917 -1518
rect 17951 -1552 17963 -1518
rect 17905 -1567 17963 -1552
rect 18163 -1382 18221 -1367
rect 18163 -1416 18175 -1382
rect 18209 -1416 18221 -1382
rect 18163 -1450 18221 -1416
rect 18163 -1484 18175 -1450
rect 18209 -1484 18221 -1450
rect 18163 -1518 18221 -1484
rect 18163 -1552 18175 -1518
rect 18209 -1552 18221 -1518
rect 18163 -1567 18221 -1552
rect 959 -2338 1017 -2323
rect 959 -2372 971 -2338
rect 1005 -2372 1017 -2338
rect 959 -2406 1017 -2372
rect 959 -2440 971 -2406
rect 1005 -2440 1017 -2406
rect 959 -2474 1017 -2440
rect 959 -2508 971 -2474
rect 1005 -2508 1017 -2474
rect 959 -2523 1017 -2508
rect 1217 -2338 1275 -2323
rect 1217 -2372 1229 -2338
rect 1263 -2372 1275 -2338
rect 1217 -2406 1275 -2372
rect 1217 -2440 1229 -2406
rect 1263 -2440 1275 -2406
rect 1217 -2474 1275 -2440
rect 1217 -2508 1229 -2474
rect 1263 -2508 1275 -2474
rect 1217 -2523 1275 -2508
rect 1411 -2338 1469 -2323
rect 1411 -2372 1423 -2338
rect 1457 -2372 1469 -2338
rect 1411 -2406 1469 -2372
rect 1411 -2440 1423 -2406
rect 1457 -2440 1469 -2406
rect 1411 -2474 1469 -2440
rect 1411 -2508 1423 -2474
rect 1457 -2508 1469 -2474
rect 1411 -2523 1469 -2508
rect 1669 -2338 1727 -2323
rect 1669 -2372 1681 -2338
rect 1715 -2372 1727 -2338
rect 1669 -2406 1727 -2372
rect 1669 -2440 1681 -2406
rect 1715 -2440 1727 -2406
rect 1669 -2474 1727 -2440
rect 1669 -2508 1681 -2474
rect 1715 -2508 1727 -2474
rect 1669 -2523 1727 -2508
rect 1927 -2338 1985 -2323
rect 1927 -2372 1939 -2338
rect 1973 -2372 1985 -2338
rect 1927 -2406 1985 -2372
rect 1927 -2440 1939 -2406
rect 1973 -2440 1985 -2406
rect 1927 -2474 1985 -2440
rect 1927 -2508 1939 -2474
rect 1973 -2508 1985 -2474
rect 1927 -2523 1985 -2508
rect 2185 -2338 2243 -2323
rect 2185 -2372 2197 -2338
rect 2231 -2372 2243 -2338
rect 2185 -2406 2243 -2372
rect 2185 -2440 2197 -2406
rect 2231 -2440 2243 -2406
rect 2185 -2474 2243 -2440
rect 2185 -2508 2197 -2474
rect 2231 -2508 2243 -2474
rect 2185 -2523 2243 -2508
rect 2443 -2338 2501 -2323
rect 2443 -2372 2455 -2338
rect 2489 -2372 2501 -2338
rect 2443 -2406 2501 -2372
rect 2443 -2440 2455 -2406
rect 2489 -2440 2501 -2406
rect 2443 -2474 2501 -2440
rect 2443 -2508 2455 -2474
rect 2489 -2508 2501 -2474
rect 2443 -2523 2501 -2508
rect 2637 -2338 2695 -2323
rect 2637 -2372 2649 -2338
rect 2683 -2372 2695 -2338
rect 2637 -2406 2695 -2372
rect 2637 -2440 2649 -2406
rect 2683 -2440 2695 -2406
rect 2637 -2474 2695 -2440
rect 2637 -2508 2649 -2474
rect 2683 -2508 2695 -2474
rect 2637 -2523 2695 -2508
rect 2895 -2338 2953 -2323
rect 2895 -2372 2907 -2338
rect 2941 -2372 2953 -2338
rect 2895 -2406 2953 -2372
rect 2895 -2440 2907 -2406
rect 2941 -2440 2953 -2406
rect 2895 -2474 2953 -2440
rect 2895 -2508 2907 -2474
rect 2941 -2508 2953 -2474
rect 2895 -2523 2953 -2508
rect 3153 -2338 3211 -2323
rect 3153 -2372 3165 -2338
rect 3199 -2372 3211 -2338
rect 3153 -2406 3211 -2372
rect 3153 -2440 3165 -2406
rect 3199 -2440 3211 -2406
rect 3153 -2474 3211 -2440
rect 3153 -2508 3165 -2474
rect 3199 -2508 3211 -2474
rect 3153 -2523 3211 -2508
rect 3411 -2338 3469 -2323
rect 3411 -2372 3423 -2338
rect 3457 -2372 3469 -2338
rect 3411 -2406 3469 -2372
rect 3411 -2440 3423 -2406
rect 3457 -2440 3469 -2406
rect 3411 -2474 3469 -2440
rect 3411 -2508 3423 -2474
rect 3457 -2508 3469 -2474
rect 3411 -2523 3469 -2508
rect 3605 -2338 3663 -2323
rect 3605 -2372 3617 -2338
rect 3651 -2372 3663 -2338
rect 3605 -2406 3663 -2372
rect 3605 -2440 3617 -2406
rect 3651 -2440 3663 -2406
rect 3605 -2474 3663 -2440
rect 3605 -2508 3617 -2474
rect 3651 -2508 3663 -2474
rect 3605 -2523 3663 -2508
rect 3863 -2338 3921 -2323
rect 3863 -2372 3875 -2338
rect 3909 -2372 3921 -2338
rect 3863 -2406 3921 -2372
rect 3863 -2440 3875 -2406
rect 3909 -2440 3921 -2406
rect 3863 -2474 3921 -2440
rect 3863 -2508 3875 -2474
rect 3909 -2508 3921 -2474
rect 3863 -2523 3921 -2508
rect 4121 -2338 4179 -2323
rect 4121 -2372 4133 -2338
rect 4167 -2372 4179 -2338
rect 4121 -2406 4179 -2372
rect 4121 -2440 4133 -2406
rect 4167 -2440 4179 -2406
rect 4121 -2474 4179 -2440
rect 4121 -2508 4133 -2474
rect 4167 -2508 4179 -2474
rect 4121 -2523 4179 -2508
rect 4379 -2338 4437 -2323
rect 4379 -2372 4391 -2338
rect 4425 -2372 4437 -2338
rect 4379 -2406 4437 -2372
rect 4379 -2440 4391 -2406
rect 4425 -2440 4437 -2406
rect 4379 -2474 4437 -2440
rect 4379 -2508 4391 -2474
rect 4425 -2508 4437 -2474
rect 4379 -2523 4437 -2508
rect 4637 -2338 4695 -2323
rect 4637 -2372 4649 -2338
rect 4683 -2372 4695 -2338
rect 4637 -2406 4695 -2372
rect 4637 -2440 4649 -2406
rect 4683 -2440 4695 -2406
rect 4637 -2474 4695 -2440
rect 4637 -2508 4649 -2474
rect 4683 -2508 4695 -2474
rect 4637 -2523 4695 -2508
rect 4830 -2338 4888 -2323
rect 4830 -2372 4842 -2338
rect 4876 -2372 4888 -2338
rect 4830 -2406 4888 -2372
rect 4830 -2440 4842 -2406
rect 4876 -2440 4888 -2406
rect 4830 -2474 4888 -2440
rect 4830 -2508 4842 -2474
rect 4876 -2508 4888 -2474
rect 4830 -2523 4888 -2508
rect 5088 -2338 5146 -2323
rect 5088 -2372 5100 -2338
rect 5134 -2372 5146 -2338
rect 5088 -2406 5146 -2372
rect 5088 -2440 5100 -2406
rect 5134 -2440 5146 -2406
rect 5088 -2474 5146 -2440
rect 5088 -2508 5100 -2474
rect 5134 -2508 5146 -2474
rect 5088 -2523 5146 -2508
rect 5316 -2338 5374 -2323
rect 5316 -2372 5328 -2338
rect 5362 -2372 5374 -2338
rect 5316 -2406 5374 -2372
rect 5316 -2440 5328 -2406
rect 5362 -2440 5374 -2406
rect 5316 -2474 5374 -2440
rect 5316 -2508 5328 -2474
rect 5362 -2508 5374 -2474
rect 5316 -2523 5374 -2508
rect 5574 -2338 5632 -2323
rect 5574 -2372 5586 -2338
rect 5620 -2372 5632 -2338
rect 5574 -2406 5632 -2372
rect 5574 -2440 5586 -2406
rect 5620 -2440 5632 -2406
rect 5574 -2474 5632 -2440
rect 5574 -2508 5586 -2474
rect 5620 -2508 5632 -2474
rect 5574 -2523 5632 -2508
rect 5768 -2338 5826 -2323
rect 5768 -2372 5780 -2338
rect 5814 -2372 5826 -2338
rect 5768 -2406 5826 -2372
rect 5768 -2440 5780 -2406
rect 5814 -2440 5826 -2406
rect 5768 -2474 5826 -2440
rect 5768 -2508 5780 -2474
rect 5814 -2508 5826 -2474
rect 5768 -2523 5826 -2508
rect 6026 -2338 6084 -2323
rect 6026 -2372 6038 -2338
rect 6072 -2372 6084 -2338
rect 6026 -2406 6084 -2372
rect 6026 -2440 6038 -2406
rect 6072 -2440 6084 -2406
rect 6026 -2474 6084 -2440
rect 6026 -2508 6038 -2474
rect 6072 -2508 6084 -2474
rect 6026 -2523 6084 -2508
rect 6284 -2338 6342 -2323
rect 6284 -2372 6296 -2338
rect 6330 -2372 6342 -2338
rect 6284 -2406 6342 -2372
rect 6284 -2440 6296 -2406
rect 6330 -2440 6342 -2406
rect 6284 -2474 6342 -2440
rect 6284 -2508 6296 -2474
rect 6330 -2508 6342 -2474
rect 6284 -2523 6342 -2508
rect 6542 -2338 6600 -2323
rect 6542 -2372 6554 -2338
rect 6588 -2372 6600 -2338
rect 6542 -2406 6600 -2372
rect 6542 -2440 6554 -2406
rect 6588 -2440 6600 -2406
rect 6542 -2474 6600 -2440
rect 6542 -2508 6554 -2474
rect 6588 -2508 6600 -2474
rect 6542 -2523 6600 -2508
rect 6800 -2338 6858 -2323
rect 6800 -2372 6812 -2338
rect 6846 -2372 6858 -2338
rect 6800 -2406 6858 -2372
rect 6800 -2440 6812 -2406
rect 6846 -2440 6858 -2406
rect 6800 -2474 6858 -2440
rect 6800 -2508 6812 -2474
rect 6846 -2508 6858 -2474
rect 6800 -2523 6858 -2508
rect 6994 -2338 7052 -2323
rect 6994 -2372 7006 -2338
rect 7040 -2372 7052 -2338
rect 6994 -2406 7052 -2372
rect 6994 -2440 7006 -2406
rect 7040 -2440 7052 -2406
rect 6994 -2474 7052 -2440
rect 6994 -2508 7006 -2474
rect 7040 -2508 7052 -2474
rect 6994 -2523 7052 -2508
rect 7252 -2338 7310 -2323
rect 7252 -2372 7264 -2338
rect 7298 -2372 7310 -2338
rect 7252 -2406 7310 -2372
rect 7252 -2440 7264 -2406
rect 7298 -2440 7310 -2406
rect 7252 -2474 7310 -2440
rect 7252 -2508 7264 -2474
rect 7298 -2508 7310 -2474
rect 7252 -2523 7310 -2508
rect 7510 -2338 7568 -2323
rect 7510 -2372 7522 -2338
rect 7556 -2372 7568 -2338
rect 7510 -2406 7568 -2372
rect 7510 -2440 7522 -2406
rect 7556 -2440 7568 -2406
rect 7510 -2474 7568 -2440
rect 7510 -2508 7522 -2474
rect 7556 -2508 7568 -2474
rect 7510 -2523 7568 -2508
rect 7768 -2338 7826 -2323
rect 7768 -2372 7780 -2338
rect 7814 -2372 7826 -2338
rect 7768 -2406 7826 -2372
rect 7768 -2440 7780 -2406
rect 7814 -2440 7826 -2406
rect 7768 -2474 7826 -2440
rect 7768 -2508 7780 -2474
rect 7814 -2508 7826 -2474
rect 7768 -2523 7826 -2508
rect 7962 -2338 8020 -2323
rect 7962 -2372 7974 -2338
rect 8008 -2372 8020 -2338
rect 7962 -2406 8020 -2372
rect 7962 -2440 7974 -2406
rect 8008 -2440 8020 -2406
rect 7962 -2474 8020 -2440
rect 7962 -2508 7974 -2474
rect 8008 -2508 8020 -2474
rect 7962 -2523 8020 -2508
rect 8220 -2338 8278 -2323
rect 8220 -2372 8232 -2338
rect 8266 -2372 8278 -2338
rect 8220 -2406 8278 -2372
rect 8220 -2440 8232 -2406
rect 8266 -2440 8278 -2406
rect 8220 -2474 8278 -2440
rect 8220 -2508 8232 -2474
rect 8266 -2508 8278 -2474
rect 8220 -2523 8278 -2508
rect 8478 -2338 8536 -2323
rect 8478 -2372 8490 -2338
rect 8524 -2372 8536 -2338
rect 8478 -2406 8536 -2372
rect 8478 -2440 8490 -2406
rect 8524 -2440 8536 -2406
rect 8478 -2474 8536 -2440
rect 8478 -2508 8490 -2474
rect 8524 -2508 8536 -2474
rect 8478 -2523 8536 -2508
rect 8736 -2338 8794 -2323
rect 8736 -2372 8748 -2338
rect 8782 -2372 8794 -2338
rect 8736 -2406 8794 -2372
rect 8736 -2440 8748 -2406
rect 8782 -2440 8794 -2406
rect 8736 -2474 8794 -2440
rect 8736 -2508 8748 -2474
rect 8782 -2508 8794 -2474
rect 8736 -2523 8794 -2508
rect 8994 -2338 9052 -2323
rect 8994 -2372 9006 -2338
rect 9040 -2372 9052 -2338
rect 8994 -2406 9052 -2372
rect 8994 -2440 9006 -2406
rect 9040 -2440 9052 -2406
rect 8994 -2474 9052 -2440
rect 8994 -2508 9006 -2474
rect 9040 -2508 9052 -2474
rect 8994 -2523 9052 -2508
rect 9188 -2338 9246 -2323
rect 9188 -2372 9200 -2338
rect 9234 -2372 9246 -2338
rect 9188 -2406 9246 -2372
rect 9188 -2440 9200 -2406
rect 9234 -2440 9246 -2406
rect 9188 -2474 9246 -2440
rect 9188 -2508 9200 -2474
rect 9234 -2508 9246 -2474
rect 9188 -2523 9246 -2508
rect 9446 -2338 9504 -2323
rect 9446 -2372 9458 -2338
rect 9492 -2372 9504 -2338
rect 9446 -2406 9504 -2372
rect 9446 -2440 9458 -2406
rect 9492 -2440 9504 -2406
rect 9446 -2474 9504 -2440
rect 9446 -2508 9458 -2474
rect 9492 -2508 9504 -2474
rect 9446 -2523 9504 -2508
rect 9676 -2338 9734 -2323
rect 9676 -2372 9688 -2338
rect 9722 -2372 9734 -2338
rect 9676 -2406 9734 -2372
rect 9676 -2440 9688 -2406
rect 9722 -2440 9734 -2406
rect 9676 -2474 9734 -2440
rect 9676 -2508 9688 -2474
rect 9722 -2508 9734 -2474
rect 9676 -2523 9734 -2508
rect 9934 -2338 9992 -2323
rect 9934 -2372 9946 -2338
rect 9980 -2372 9992 -2338
rect 9934 -2406 9992 -2372
rect 9934 -2440 9946 -2406
rect 9980 -2440 9992 -2406
rect 9934 -2474 9992 -2440
rect 9934 -2508 9946 -2474
rect 9980 -2508 9992 -2474
rect 9934 -2523 9992 -2508
rect 10128 -2338 10186 -2323
rect 10128 -2372 10140 -2338
rect 10174 -2372 10186 -2338
rect 10128 -2406 10186 -2372
rect 10128 -2440 10140 -2406
rect 10174 -2440 10186 -2406
rect 10128 -2474 10186 -2440
rect 10128 -2508 10140 -2474
rect 10174 -2508 10186 -2474
rect 10128 -2523 10186 -2508
rect 10386 -2338 10444 -2323
rect 10386 -2372 10398 -2338
rect 10432 -2372 10444 -2338
rect 10386 -2406 10444 -2372
rect 10386 -2440 10398 -2406
rect 10432 -2440 10444 -2406
rect 10386 -2474 10444 -2440
rect 10386 -2508 10398 -2474
rect 10432 -2508 10444 -2474
rect 10386 -2523 10444 -2508
rect 10644 -2338 10702 -2323
rect 10644 -2372 10656 -2338
rect 10690 -2372 10702 -2338
rect 10644 -2406 10702 -2372
rect 10644 -2440 10656 -2406
rect 10690 -2440 10702 -2406
rect 10644 -2474 10702 -2440
rect 10644 -2508 10656 -2474
rect 10690 -2508 10702 -2474
rect 10644 -2523 10702 -2508
rect 10902 -2338 10960 -2323
rect 10902 -2372 10914 -2338
rect 10948 -2372 10960 -2338
rect 10902 -2406 10960 -2372
rect 10902 -2440 10914 -2406
rect 10948 -2440 10960 -2406
rect 10902 -2474 10960 -2440
rect 10902 -2508 10914 -2474
rect 10948 -2508 10960 -2474
rect 10902 -2523 10960 -2508
rect 11160 -2338 11218 -2323
rect 11160 -2372 11172 -2338
rect 11206 -2372 11218 -2338
rect 11160 -2406 11218 -2372
rect 11160 -2440 11172 -2406
rect 11206 -2440 11218 -2406
rect 11160 -2474 11218 -2440
rect 11160 -2508 11172 -2474
rect 11206 -2508 11218 -2474
rect 11160 -2523 11218 -2508
rect 11354 -2338 11412 -2323
rect 11354 -2372 11366 -2338
rect 11400 -2372 11412 -2338
rect 11354 -2406 11412 -2372
rect 11354 -2440 11366 -2406
rect 11400 -2440 11412 -2406
rect 11354 -2474 11412 -2440
rect 11354 -2508 11366 -2474
rect 11400 -2508 11412 -2474
rect 11354 -2523 11412 -2508
rect 11612 -2338 11670 -2323
rect 11612 -2372 11624 -2338
rect 11658 -2372 11670 -2338
rect 11612 -2406 11670 -2372
rect 11612 -2440 11624 -2406
rect 11658 -2440 11670 -2406
rect 11612 -2474 11670 -2440
rect 11612 -2508 11624 -2474
rect 11658 -2508 11670 -2474
rect 11612 -2523 11670 -2508
rect 11870 -2338 11928 -2323
rect 11870 -2372 11882 -2338
rect 11916 -2372 11928 -2338
rect 11870 -2406 11928 -2372
rect 11870 -2440 11882 -2406
rect 11916 -2440 11928 -2406
rect 11870 -2474 11928 -2440
rect 11870 -2508 11882 -2474
rect 11916 -2508 11928 -2474
rect 11870 -2523 11928 -2508
rect 12128 -2338 12186 -2323
rect 12128 -2372 12140 -2338
rect 12174 -2372 12186 -2338
rect 12128 -2406 12186 -2372
rect 12128 -2440 12140 -2406
rect 12174 -2440 12186 -2406
rect 12128 -2474 12186 -2440
rect 12128 -2508 12140 -2474
rect 12174 -2508 12186 -2474
rect 12128 -2523 12186 -2508
rect 12322 -2338 12380 -2323
rect 12322 -2372 12334 -2338
rect 12368 -2372 12380 -2338
rect 12322 -2406 12380 -2372
rect 12322 -2440 12334 -2406
rect 12368 -2440 12380 -2406
rect 12322 -2474 12380 -2440
rect 12322 -2508 12334 -2474
rect 12368 -2508 12380 -2474
rect 12322 -2523 12380 -2508
rect 12580 -2338 12638 -2323
rect 12580 -2372 12592 -2338
rect 12626 -2372 12638 -2338
rect 12580 -2406 12638 -2372
rect 12580 -2440 12592 -2406
rect 12626 -2440 12638 -2406
rect 12580 -2474 12638 -2440
rect 12580 -2508 12592 -2474
rect 12626 -2508 12638 -2474
rect 12580 -2523 12638 -2508
rect 12838 -2338 12896 -2323
rect 12838 -2372 12850 -2338
rect 12884 -2372 12896 -2338
rect 12838 -2406 12896 -2372
rect 12838 -2440 12850 -2406
rect 12884 -2440 12896 -2406
rect 12838 -2474 12896 -2440
rect 12838 -2508 12850 -2474
rect 12884 -2508 12896 -2474
rect 12838 -2523 12896 -2508
rect 13096 -2338 13154 -2323
rect 13096 -2372 13108 -2338
rect 13142 -2372 13154 -2338
rect 13096 -2406 13154 -2372
rect 13096 -2440 13108 -2406
rect 13142 -2440 13154 -2406
rect 13096 -2474 13154 -2440
rect 13096 -2508 13108 -2474
rect 13142 -2508 13154 -2474
rect 13096 -2523 13154 -2508
rect 13354 -2338 13412 -2323
rect 13354 -2372 13366 -2338
rect 13400 -2372 13412 -2338
rect 13354 -2406 13412 -2372
rect 13354 -2440 13366 -2406
rect 13400 -2440 13412 -2406
rect 13354 -2474 13412 -2440
rect 13354 -2508 13366 -2474
rect 13400 -2508 13412 -2474
rect 13354 -2523 13412 -2508
rect 13548 -2338 13606 -2323
rect 13548 -2372 13560 -2338
rect 13594 -2372 13606 -2338
rect 13548 -2406 13606 -2372
rect 13548 -2440 13560 -2406
rect 13594 -2440 13606 -2406
rect 13548 -2474 13606 -2440
rect 13548 -2508 13560 -2474
rect 13594 -2508 13606 -2474
rect 13548 -2523 13606 -2508
rect 13806 -2338 13864 -2323
rect 13806 -2372 13818 -2338
rect 13852 -2372 13864 -2338
rect 13806 -2406 13864 -2372
rect 13806 -2440 13818 -2406
rect 13852 -2440 13864 -2406
rect 13806 -2474 13864 -2440
rect 13806 -2508 13818 -2474
rect 13852 -2508 13864 -2474
rect 13806 -2523 13864 -2508
rect 14034 -2338 14092 -2323
rect 14034 -2372 14046 -2338
rect 14080 -2372 14092 -2338
rect 14034 -2406 14092 -2372
rect 14034 -2440 14046 -2406
rect 14080 -2440 14092 -2406
rect 14034 -2474 14092 -2440
rect 14034 -2508 14046 -2474
rect 14080 -2508 14092 -2474
rect 14034 -2523 14092 -2508
rect 14292 -2338 14350 -2323
rect 14292 -2372 14304 -2338
rect 14338 -2372 14350 -2338
rect 14292 -2406 14350 -2372
rect 14292 -2440 14304 -2406
rect 14338 -2440 14350 -2406
rect 14292 -2474 14350 -2440
rect 14292 -2508 14304 -2474
rect 14338 -2508 14350 -2474
rect 14292 -2523 14350 -2508
rect 14485 -2338 14543 -2323
rect 14485 -2372 14497 -2338
rect 14531 -2372 14543 -2338
rect 14485 -2406 14543 -2372
rect 14485 -2440 14497 -2406
rect 14531 -2440 14543 -2406
rect 14485 -2474 14543 -2440
rect 14485 -2508 14497 -2474
rect 14531 -2508 14543 -2474
rect 14485 -2523 14543 -2508
rect 14743 -2338 14801 -2323
rect 14743 -2372 14755 -2338
rect 14789 -2372 14801 -2338
rect 14743 -2406 14801 -2372
rect 14743 -2440 14755 -2406
rect 14789 -2440 14801 -2406
rect 14743 -2474 14801 -2440
rect 14743 -2508 14755 -2474
rect 14789 -2508 14801 -2474
rect 14743 -2523 14801 -2508
rect 15001 -2338 15059 -2323
rect 15001 -2372 15013 -2338
rect 15047 -2372 15059 -2338
rect 15001 -2406 15059 -2372
rect 15001 -2440 15013 -2406
rect 15047 -2440 15059 -2406
rect 15001 -2474 15059 -2440
rect 15001 -2508 15013 -2474
rect 15047 -2508 15059 -2474
rect 15001 -2523 15059 -2508
rect 15259 -2338 15317 -2323
rect 15259 -2372 15271 -2338
rect 15305 -2372 15317 -2338
rect 15259 -2406 15317 -2372
rect 15259 -2440 15271 -2406
rect 15305 -2440 15317 -2406
rect 15259 -2474 15317 -2440
rect 15259 -2508 15271 -2474
rect 15305 -2508 15317 -2474
rect 15259 -2523 15317 -2508
rect 15517 -2338 15575 -2323
rect 15517 -2372 15529 -2338
rect 15563 -2372 15575 -2338
rect 15517 -2406 15575 -2372
rect 15517 -2440 15529 -2406
rect 15563 -2440 15575 -2406
rect 15517 -2474 15575 -2440
rect 15517 -2508 15529 -2474
rect 15563 -2508 15575 -2474
rect 15517 -2523 15575 -2508
rect 15711 -2338 15769 -2323
rect 15711 -2372 15723 -2338
rect 15757 -2372 15769 -2338
rect 15711 -2406 15769 -2372
rect 15711 -2440 15723 -2406
rect 15757 -2440 15769 -2406
rect 15711 -2474 15769 -2440
rect 15711 -2508 15723 -2474
rect 15757 -2508 15769 -2474
rect 15711 -2523 15769 -2508
rect 15969 -2338 16027 -2323
rect 15969 -2372 15981 -2338
rect 16015 -2372 16027 -2338
rect 15969 -2406 16027 -2372
rect 15969 -2440 15981 -2406
rect 16015 -2440 16027 -2406
rect 15969 -2474 16027 -2440
rect 15969 -2508 15981 -2474
rect 16015 -2508 16027 -2474
rect 15969 -2523 16027 -2508
rect 16227 -2338 16285 -2323
rect 16227 -2372 16239 -2338
rect 16273 -2372 16285 -2338
rect 16227 -2406 16285 -2372
rect 16227 -2440 16239 -2406
rect 16273 -2440 16285 -2406
rect 16227 -2474 16285 -2440
rect 16227 -2508 16239 -2474
rect 16273 -2508 16285 -2474
rect 16227 -2523 16285 -2508
rect 16485 -2338 16543 -2323
rect 16485 -2372 16497 -2338
rect 16531 -2372 16543 -2338
rect 16485 -2406 16543 -2372
rect 16485 -2440 16497 -2406
rect 16531 -2440 16543 -2406
rect 16485 -2474 16543 -2440
rect 16485 -2508 16497 -2474
rect 16531 -2508 16543 -2474
rect 16485 -2523 16543 -2508
rect 16679 -2338 16737 -2323
rect 16679 -2372 16691 -2338
rect 16725 -2372 16737 -2338
rect 16679 -2406 16737 -2372
rect 16679 -2440 16691 -2406
rect 16725 -2440 16737 -2406
rect 16679 -2474 16737 -2440
rect 16679 -2508 16691 -2474
rect 16725 -2508 16737 -2474
rect 16679 -2523 16737 -2508
rect 16937 -2338 16995 -2323
rect 16937 -2372 16949 -2338
rect 16983 -2372 16995 -2338
rect 16937 -2406 16995 -2372
rect 16937 -2440 16949 -2406
rect 16983 -2440 16995 -2406
rect 16937 -2474 16995 -2440
rect 16937 -2508 16949 -2474
rect 16983 -2508 16995 -2474
rect 16937 -2523 16995 -2508
rect 17195 -2338 17253 -2323
rect 17195 -2372 17207 -2338
rect 17241 -2372 17253 -2338
rect 17195 -2406 17253 -2372
rect 17195 -2440 17207 -2406
rect 17241 -2440 17253 -2406
rect 17195 -2474 17253 -2440
rect 17195 -2508 17207 -2474
rect 17241 -2508 17253 -2474
rect 17195 -2523 17253 -2508
rect 17453 -2338 17511 -2323
rect 17453 -2372 17465 -2338
rect 17499 -2372 17511 -2338
rect 17453 -2406 17511 -2372
rect 17453 -2440 17465 -2406
rect 17499 -2440 17511 -2406
rect 17453 -2474 17511 -2440
rect 17453 -2508 17465 -2474
rect 17499 -2508 17511 -2474
rect 17453 -2523 17511 -2508
rect 17711 -2338 17769 -2323
rect 17711 -2372 17723 -2338
rect 17757 -2372 17769 -2338
rect 17711 -2406 17769 -2372
rect 17711 -2440 17723 -2406
rect 17757 -2440 17769 -2406
rect 17711 -2474 17769 -2440
rect 17711 -2508 17723 -2474
rect 17757 -2508 17769 -2474
rect 17711 -2523 17769 -2508
rect 17905 -2338 17963 -2323
rect 17905 -2372 17917 -2338
rect 17951 -2372 17963 -2338
rect 17905 -2406 17963 -2372
rect 17905 -2440 17917 -2406
rect 17951 -2440 17963 -2406
rect 17905 -2474 17963 -2440
rect 17905 -2508 17917 -2474
rect 17951 -2508 17963 -2474
rect 17905 -2523 17963 -2508
rect 18163 -2338 18221 -2323
rect 18163 -2372 18175 -2338
rect 18209 -2372 18221 -2338
rect 18163 -2406 18221 -2372
rect 18163 -2440 18175 -2406
rect 18209 -2440 18221 -2406
rect 18163 -2474 18221 -2440
rect 18163 -2508 18175 -2474
rect 18209 -2508 18221 -2474
rect 18163 -2523 18221 -2508
rect 959 -3029 1017 -3014
rect 959 -3063 971 -3029
rect 1005 -3063 1017 -3029
rect 959 -3097 1017 -3063
rect 959 -3131 971 -3097
rect 1005 -3131 1017 -3097
rect 959 -3165 1017 -3131
rect 959 -3199 971 -3165
rect 1005 -3199 1017 -3165
rect 959 -3214 1017 -3199
rect 1217 -3029 1275 -3014
rect 1217 -3063 1229 -3029
rect 1263 -3063 1275 -3029
rect 1217 -3097 1275 -3063
rect 1217 -3131 1229 -3097
rect 1263 -3131 1275 -3097
rect 1217 -3165 1275 -3131
rect 1217 -3199 1229 -3165
rect 1263 -3199 1275 -3165
rect 1217 -3214 1275 -3199
rect 1411 -3029 1469 -3014
rect 1411 -3063 1423 -3029
rect 1457 -3063 1469 -3029
rect 1411 -3097 1469 -3063
rect 1411 -3131 1423 -3097
rect 1457 -3131 1469 -3097
rect 1411 -3165 1469 -3131
rect 1411 -3199 1423 -3165
rect 1457 -3199 1469 -3165
rect 1411 -3214 1469 -3199
rect 1669 -3029 1727 -3014
rect 1669 -3063 1681 -3029
rect 1715 -3063 1727 -3029
rect 1669 -3097 1727 -3063
rect 1669 -3131 1681 -3097
rect 1715 -3131 1727 -3097
rect 1669 -3165 1727 -3131
rect 1669 -3199 1681 -3165
rect 1715 -3199 1727 -3165
rect 1669 -3214 1727 -3199
rect 1927 -3029 1985 -3014
rect 1927 -3063 1939 -3029
rect 1973 -3063 1985 -3029
rect 1927 -3097 1985 -3063
rect 1927 -3131 1939 -3097
rect 1973 -3131 1985 -3097
rect 1927 -3165 1985 -3131
rect 1927 -3199 1939 -3165
rect 1973 -3199 1985 -3165
rect 1927 -3214 1985 -3199
rect 2185 -3029 2243 -3014
rect 2185 -3063 2197 -3029
rect 2231 -3063 2243 -3029
rect 2185 -3097 2243 -3063
rect 2185 -3131 2197 -3097
rect 2231 -3131 2243 -3097
rect 2185 -3165 2243 -3131
rect 2185 -3199 2197 -3165
rect 2231 -3199 2243 -3165
rect 2185 -3214 2243 -3199
rect 2443 -3029 2501 -3014
rect 2443 -3063 2455 -3029
rect 2489 -3063 2501 -3029
rect 2443 -3097 2501 -3063
rect 2443 -3131 2455 -3097
rect 2489 -3131 2501 -3097
rect 2443 -3165 2501 -3131
rect 2443 -3199 2455 -3165
rect 2489 -3199 2501 -3165
rect 2443 -3214 2501 -3199
rect 2637 -3029 2695 -3014
rect 2637 -3063 2649 -3029
rect 2683 -3063 2695 -3029
rect 2637 -3097 2695 -3063
rect 2637 -3131 2649 -3097
rect 2683 -3131 2695 -3097
rect 2637 -3165 2695 -3131
rect 2637 -3199 2649 -3165
rect 2683 -3199 2695 -3165
rect 2637 -3214 2695 -3199
rect 2895 -3029 2953 -3014
rect 2895 -3063 2907 -3029
rect 2941 -3063 2953 -3029
rect 2895 -3097 2953 -3063
rect 2895 -3131 2907 -3097
rect 2941 -3131 2953 -3097
rect 2895 -3165 2953 -3131
rect 2895 -3199 2907 -3165
rect 2941 -3199 2953 -3165
rect 2895 -3214 2953 -3199
rect 3153 -3029 3211 -3014
rect 3153 -3063 3165 -3029
rect 3199 -3063 3211 -3029
rect 3153 -3097 3211 -3063
rect 3153 -3131 3165 -3097
rect 3199 -3131 3211 -3097
rect 3153 -3165 3211 -3131
rect 3153 -3199 3165 -3165
rect 3199 -3199 3211 -3165
rect 3153 -3214 3211 -3199
rect 3411 -3029 3469 -3014
rect 3411 -3063 3423 -3029
rect 3457 -3063 3469 -3029
rect 3411 -3097 3469 -3063
rect 3411 -3131 3423 -3097
rect 3457 -3131 3469 -3097
rect 3411 -3165 3469 -3131
rect 3411 -3199 3423 -3165
rect 3457 -3199 3469 -3165
rect 3411 -3214 3469 -3199
rect 3605 -3029 3663 -3014
rect 3605 -3063 3617 -3029
rect 3651 -3063 3663 -3029
rect 3605 -3097 3663 -3063
rect 3605 -3131 3617 -3097
rect 3651 -3131 3663 -3097
rect 3605 -3165 3663 -3131
rect 3605 -3199 3617 -3165
rect 3651 -3199 3663 -3165
rect 3605 -3214 3663 -3199
rect 3863 -3029 3921 -3014
rect 3863 -3063 3875 -3029
rect 3909 -3063 3921 -3029
rect 3863 -3097 3921 -3063
rect 3863 -3131 3875 -3097
rect 3909 -3131 3921 -3097
rect 3863 -3165 3921 -3131
rect 3863 -3199 3875 -3165
rect 3909 -3199 3921 -3165
rect 3863 -3214 3921 -3199
rect 4121 -3029 4179 -3014
rect 4121 -3063 4133 -3029
rect 4167 -3063 4179 -3029
rect 4121 -3097 4179 -3063
rect 4121 -3131 4133 -3097
rect 4167 -3131 4179 -3097
rect 4121 -3165 4179 -3131
rect 4121 -3199 4133 -3165
rect 4167 -3199 4179 -3165
rect 4121 -3214 4179 -3199
rect 4379 -3029 4437 -3014
rect 4379 -3063 4391 -3029
rect 4425 -3063 4437 -3029
rect 4379 -3097 4437 -3063
rect 4379 -3131 4391 -3097
rect 4425 -3131 4437 -3097
rect 4379 -3165 4437 -3131
rect 4379 -3199 4391 -3165
rect 4425 -3199 4437 -3165
rect 4379 -3214 4437 -3199
rect 4637 -3029 4695 -3014
rect 4637 -3063 4649 -3029
rect 4683 -3063 4695 -3029
rect 4637 -3097 4695 -3063
rect 4637 -3131 4649 -3097
rect 4683 -3131 4695 -3097
rect 4637 -3165 4695 -3131
rect 4637 -3199 4649 -3165
rect 4683 -3199 4695 -3165
rect 4637 -3214 4695 -3199
rect 4830 -3029 4888 -3014
rect 4830 -3063 4842 -3029
rect 4876 -3063 4888 -3029
rect 4830 -3097 4888 -3063
rect 4830 -3131 4842 -3097
rect 4876 -3131 4888 -3097
rect 4830 -3165 4888 -3131
rect 4830 -3199 4842 -3165
rect 4876 -3199 4888 -3165
rect 4830 -3214 4888 -3199
rect 5088 -3029 5146 -3014
rect 5088 -3063 5100 -3029
rect 5134 -3063 5146 -3029
rect 5088 -3097 5146 -3063
rect 5088 -3131 5100 -3097
rect 5134 -3131 5146 -3097
rect 5088 -3165 5146 -3131
rect 5088 -3199 5100 -3165
rect 5134 -3199 5146 -3165
rect 5088 -3214 5146 -3199
rect 5316 -3029 5374 -3014
rect 5316 -3063 5328 -3029
rect 5362 -3063 5374 -3029
rect 5316 -3097 5374 -3063
rect 5316 -3131 5328 -3097
rect 5362 -3131 5374 -3097
rect 5316 -3165 5374 -3131
rect 5316 -3199 5328 -3165
rect 5362 -3199 5374 -3165
rect 5316 -3214 5374 -3199
rect 5574 -3029 5632 -3014
rect 5574 -3063 5586 -3029
rect 5620 -3063 5632 -3029
rect 5574 -3097 5632 -3063
rect 5574 -3131 5586 -3097
rect 5620 -3131 5632 -3097
rect 5574 -3165 5632 -3131
rect 5574 -3199 5586 -3165
rect 5620 -3199 5632 -3165
rect 5574 -3214 5632 -3199
rect 5768 -3029 5826 -3014
rect 5768 -3063 5780 -3029
rect 5814 -3063 5826 -3029
rect 5768 -3097 5826 -3063
rect 5768 -3131 5780 -3097
rect 5814 -3131 5826 -3097
rect 5768 -3165 5826 -3131
rect 5768 -3199 5780 -3165
rect 5814 -3199 5826 -3165
rect 5768 -3214 5826 -3199
rect 6026 -3029 6084 -3014
rect 6026 -3063 6038 -3029
rect 6072 -3063 6084 -3029
rect 6026 -3097 6084 -3063
rect 6026 -3131 6038 -3097
rect 6072 -3131 6084 -3097
rect 6026 -3165 6084 -3131
rect 6026 -3199 6038 -3165
rect 6072 -3199 6084 -3165
rect 6026 -3214 6084 -3199
rect 6284 -3029 6342 -3014
rect 6284 -3063 6296 -3029
rect 6330 -3063 6342 -3029
rect 6284 -3097 6342 -3063
rect 6284 -3131 6296 -3097
rect 6330 -3131 6342 -3097
rect 6284 -3165 6342 -3131
rect 6284 -3199 6296 -3165
rect 6330 -3199 6342 -3165
rect 6284 -3214 6342 -3199
rect 6542 -3029 6600 -3014
rect 6542 -3063 6554 -3029
rect 6588 -3063 6600 -3029
rect 6542 -3097 6600 -3063
rect 6542 -3131 6554 -3097
rect 6588 -3131 6600 -3097
rect 6542 -3165 6600 -3131
rect 6542 -3199 6554 -3165
rect 6588 -3199 6600 -3165
rect 6542 -3214 6600 -3199
rect 6800 -3029 6858 -3014
rect 6800 -3063 6812 -3029
rect 6846 -3063 6858 -3029
rect 6800 -3097 6858 -3063
rect 6800 -3131 6812 -3097
rect 6846 -3131 6858 -3097
rect 6800 -3165 6858 -3131
rect 6800 -3199 6812 -3165
rect 6846 -3199 6858 -3165
rect 6800 -3214 6858 -3199
rect 6994 -3029 7052 -3014
rect 6994 -3063 7006 -3029
rect 7040 -3063 7052 -3029
rect 6994 -3097 7052 -3063
rect 6994 -3131 7006 -3097
rect 7040 -3131 7052 -3097
rect 6994 -3165 7052 -3131
rect 6994 -3199 7006 -3165
rect 7040 -3199 7052 -3165
rect 6994 -3214 7052 -3199
rect 7252 -3029 7310 -3014
rect 7252 -3063 7264 -3029
rect 7298 -3063 7310 -3029
rect 7252 -3097 7310 -3063
rect 7252 -3131 7264 -3097
rect 7298 -3131 7310 -3097
rect 7252 -3165 7310 -3131
rect 7252 -3199 7264 -3165
rect 7298 -3199 7310 -3165
rect 7252 -3214 7310 -3199
rect 7510 -3029 7568 -3014
rect 7510 -3063 7522 -3029
rect 7556 -3063 7568 -3029
rect 7510 -3097 7568 -3063
rect 7510 -3131 7522 -3097
rect 7556 -3131 7568 -3097
rect 7510 -3165 7568 -3131
rect 7510 -3199 7522 -3165
rect 7556 -3199 7568 -3165
rect 7510 -3214 7568 -3199
rect 7768 -3029 7826 -3014
rect 7768 -3063 7780 -3029
rect 7814 -3063 7826 -3029
rect 7768 -3097 7826 -3063
rect 7768 -3131 7780 -3097
rect 7814 -3131 7826 -3097
rect 7768 -3165 7826 -3131
rect 7768 -3199 7780 -3165
rect 7814 -3199 7826 -3165
rect 7768 -3214 7826 -3199
rect 7962 -3029 8020 -3014
rect 7962 -3063 7974 -3029
rect 8008 -3063 8020 -3029
rect 7962 -3097 8020 -3063
rect 7962 -3131 7974 -3097
rect 8008 -3131 8020 -3097
rect 7962 -3165 8020 -3131
rect 7962 -3199 7974 -3165
rect 8008 -3199 8020 -3165
rect 7962 -3214 8020 -3199
rect 8220 -3029 8278 -3014
rect 8220 -3063 8232 -3029
rect 8266 -3063 8278 -3029
rect 8220 -3097 8278 -3063
rect 8220 -3131 8232 -3097
rect 8266 -3131 8278 -3097
rect 8220 -3165 8278 -3131
rect 8220 -3199 8232 -3165
rect 8266 -3199 8278 -3165
rect 8220 -3214 8278 -3199
rect 8478 -3029 8536 -3014
rect 8478 -3063 8490 -3029
rect 8524 -3063 8536 -3029
rect 8478 -3097 8536 -3063
rect 8478 -3131 8490 -3097
rect 8524 -3131 8536 -3097
rect 8478 -3165 8536 -3131
rect 8478 -3199 8490 -3165
rect 8524 -3199 8536 -3165
rect 8478 -3214 8536 -3199
rect 8736 -3029 8794 -3014
rect 8736 -3063 8748 -3029
rect 8782 -3063 8794 -3029
rect 8736 -3097 8794 -3063
rect 8736 -3131 8748 -3097
rect 8782 -3131 8794 -3097
rect 8736 -3165 8794 -3131
rect 8736 -3199 8748 -3165
rect 8782 -3199 8794 -3165
rect 8736 -3214 8794 -3199
rect 8994 -3029 9052 -3014
rect 8994 -3063 9006 -3029
rect 9040 -3063 9052 -3029
rect 8994 -3097 9052 -3063
rect 8994 -3131 9006 -3097
rect 9040 -3131 9052 -3097
rect 8994 -3165 9052 -3131
rect 8994 -3199 9006 -3165
rect 9040 -3199 9052 -3165
rect 8994 -3214 9052 -3199
rect 9188 -3029 9246 -3014
rect 9188 -3063 9200 -3029
rect 9234 -3063 9246 -3029
rect 9188 -3097 9246 -3063
rect 9188 -3131 9200 -3097
rect 9234 -3131 9246 -3097
rect 9188 -3165 9246 -3131
rect 9188 -3199 9200 -3165
rect 9234 -3199 9246 -3165
rect 9188 -3214 9246 -3199
rect 9446 -3029 9504 -3014
rect 9446 -3063 9458 -3029
rect 9492 -3063 9504 -3029
rect 9446 -3097 9504 -3063
rect 9446 -3131 9458 -3097
rect 9492 -3131 9504 -3097
rect 9446 -3165 9504 -3131
rect 9446 -3199 9458 -3165
rect 9492 -3199 9504 -3165
rect 9446 -3214 9504 -3199
rect 9676 -3029 9734 -3014
rect 9676 -3063 9688 -3029
rect 9722 -3063 9734 -3029
rect 9676 -3097 9734 -3063
rect 9676 -3131 9688 -3097
rect 9722 -3131 9734 -3097
rect 9676 -3165 9734 -3131
rect 9676 -3199 9688 -3165
rect 9722 -3199 9734 -3165
rect 9676 -3214 9734 -3199
rect 9934 -3029 9992 -3014
rect 9934 -3063 9946 -3029
rect 9980 -3063 9992 -3029
rect 9934 -3097 9992 -3063
rect 9934 -3131 9946 -3097
rect 9980 -3131 9992 -3097
rect 9934 -3165 9992 -3131
rect 9934 -3199 9946 -3165
rect 9980 -3199 9992 -3165
rect 9934 -3214 9992 -3199
rect 10128 -3029 10186 -3014
rect 10128 -3063 10140 -3029
rect 10174 -3063 10186 -3029
rect 10128 -3097 10186 -3063
rect 10128 -3131 10140 -3097
rect 10174 -3131 10186 -3097
rect 10128 -3165 10186 -3131
rect 10128 -3199 10140 -3165
rect 10174 -3199 10186 -3165
rect 10128 -3214 10186 -3199
rect 10386 -3029 10444 -3014
rect 10386 -3063 10398 -3029
rect 10432 -3063 10444 -3029
rect 10386 -3097 10444 -3063
rect 10386 -3131 10398 -3097
rect 10432 -3131 10444 -3097
rect 10386 -3165 10444 -3131
rect 10386 -3199 10398 -3165
rect 10432 -3199 10444 -3165
rect 10386 -3214 10444 -3199
rect 10644 -3029 10702 -3014
rect 10644 -3063 10656 -3029
rect 10690 -3063 10702 -3029
rect 10644 -3097 10702 -3063
rect 10644 -3131 10656 -3097
rect 10690 -3131 10702 -3097
rect 10644 -3165 10702 -3131
rect 10644 -3199 10656 -3165
rect 10690 -3199 10702 -3165
rect 10644 -3214 10702 -3199
rect 10902 -3029 10960 -3014
rect 10902 -3063 10914 -3029
rect 10948 -3063 10960 -3029
rect 10902 -3097 10960 -3063
rect 10902 -3131 10914 -3097
rect 10948 -3131 10960 -3097
rect 10902 -3165 10960 -3131
rect 10902 -3199 10914 -3165
rect 10948 -3199 10960 -3165
rect 10902 -3214 10960 -3199
rect 11160 -3029 11218 -3014
rect 11160 -3063 11172 -3029
rect 11206 -3063 11218 -3029
rect 11160 -3097 11218 -3063
rect 11160 -3131 11172 -3097
rect 11206 -3131 11218 -3097
rect 11160 -3165 11218 -3131
rect 11160 -3199 11172 -3165
rect 11206 -3199 11218 -3165
rect 11160 -3214 11218 -3199
rect 11354 -3029 11412 -3014
rect 11354 -3063 11366 -3029
rect 11400 -3063 11412 -3029
rect 11354 -3097 11412 -3063
rect 11354 -3131 11366 -3097
rect 11400 -3131 11412 -3097
rect 11354 -3165 11412 -3131
rect 11354 -3199 11366 -3165
rect 11400 -3199 11412 -3165
rect 11354 -3214 11412 -3199
rect 11612 -3029 11670 -3014
rect 11612 -3063 11624 -3029
rect 11658 -3063 11670 -3029
rect 11612 -3097 11670 -3063
rect 11612 -3131 11624 -3097
rect 11658 -3131 11670 -3097
rect 11612 -3165 11670 -3131
rect 11612 -3199 11624 -3165
rect 11658 -3199 11670 -3165
rect 11612 -3214 11670 -3199
rect 11870 -3029 11928 -3014
rect 11870 -3063 11882 -3029
rect 11916 -3063 11928 -3029
rect 11870 -3097 11928 -3063
rect 11870 -3131 11882 -3097
rect 11916 -3131 11928 -3097
rect 11870 -3165 11928 -3131
rect 11870 -3199 11882 -3165
rect 11916 -3199 11928 -3165
rect 11870 -3214 11928 -3199
rect 12128 -3029 12186 -3014
rect 12128 -3063 12140 -3029
rect 12174 -3063 12186 -3029
rect 12128 -3097 12186 -3063
rect 12128 -3131 12140 -3097
rect 12174 -3131 12186 -3097
rect 12128 -3165 12186 -3131
rect 12128 -3199 12140 -3165
rect 12174 -3199 12186 -3165
rect 12128 -3214 12186 -3199
rect 12322 -3029 12380 -3014
rect 12322 -3063 12334 -3029
rect 12368 -3063 12380 -3029
rect 12322 -3097 12380 -3063
rect 12322 -3131 12334 -3097
rect 12368 -3131 12380 -3097
rect 12322 -3165 12380 -3131
rect 12322 -3199 12334 -3165
rect 12368 -3199 12380 -3165
rect 12322 -3214 12380 -3199
rect 12580 -3029 12638 -3014
rect 12580 -3063 12592 -3029
rect 12626 -3063 12638 -3029
rect 12580 -3097 12638 -3063
rect 12580 -3131 12592 -3097
rect 12626 -3131 12638 -3097
rect 12580 -3165 12638 -3131
rect 12580 -3199 12592 -3165
rect 12626 -3199 12638 -3165
rect 12580 -3214 12638 -3199
rect 12838 -3029 12896 -3014
rect 12838 -3063 12850 -3029
rect 12884 -3063 12896 -3029
rect 12838 -3097 12896 -3063
rect 12838 -3131 12850 -3097
rect 12884 -3131 12896 -3097
rect 12838 -3165 12896 -3131
rect 12838 -3199 12850 -3165
rect 12884 -3199 12896 -3165
rect 12838 -3214 12896 -3199
rect 13096 -3029 13154 -3014
rect 13096 -3063 13108 -3029
rect 13142 -3063 13154 -3029
rect 13096 -3097 13154 -3063
rect 13096 -3131 13108 -3097
rect 13142 -3131 13154 -3097
rect 13096 -3165 13154 -3131
rect 13096 -3199 13108 -3165
rect 13142 -3199 13154 -3165
rect 13096 -3214 13154 -3199
rect 13354 -3029 13412 -3014
rect 13354 -3063 13366 -3029
rect 13400 -3063 13412 -3029
rect 13354 -3097 13412 -3063
rect 13354 -3131 13366 -3097
rect 13400 -3131 13412 -3097
rect 13354 -3165 13412 -3131
rect 13354 -3199 13366 -3165
rect 13400 -3199 13412 -3165
rect 13354 -3214 13412 -3199
rect 13548 -3029 13606 -3014
rect 13548 -3063 13560 -3029
rect 13594 -3063 13606 -3029
rect 13548 -3097 13606 -3063
rect 13548 -3131 13560 -3097
rect 13594 -3131 13606 -3097
rect 13548 -3165 13606 -3131
rect 13548 -3199 13560 -3165
rect 13594 -3199 13606 -3165
rect 13548 -3214 13606 -3199
rect 13806 -3029 13864 -3014
rect 13806 -3063 13818 -3029
rect 13852 -3063 13864 -3029
rect 13806 -3097 13864 -3063
rect 13806 -3131 13818 -3097
rect 13852 -3131 13864 -3097
rect 13806 -3165 13864 -3131
rect 13806 -3199 13818 -3165
rect 13852 -3199 13864 -3165
rect 13806 -3214 13864 -3199
rect 14034 -3029 14092 -3014
rect 14034 -3063 14046 -3029
rect 14080 -3063 14092 -3029
rect 14034 -3097 14092 -3063
rect 14034 -3131 14046 -3097
rect 14080 -3131 14092 -3097
rect 14034 -3165 14092 -3131
rect 14034 -3199 14046 -3165
rect 14080 -3199 14092 -3165
rect 14034 -3214 14092 -3199
rect 14292 -3029 14350 -3014
rect 14292 -3063 14304 -3029
rect 14338 -3063 14350 -3029
rect 14292 -3097 14350 -3063
rect 14292 -3131 14304 -3097
rect 14338 -3131 14350 -3097
rect 14292 -3165 14350 -3131
rect 14292 -3199 14304 -3165
rect 14338 -3199 14350 -3165
rect 14292 -3214 14350 -3199
rect 14485 -3029 14543 -3014
rect 14485 -3063 14497 -3029
rect 14531 -3063 14543 -3029
rect 14485 -3097 14543 -3063
rect 14485 -3131 14497 -3097
rect 14531 -3131 14543 -3097
rect 14485 -3165 14543 -3131
rect 14485 -3199 14497 -3165
rect 14531 -3199 14543 -3165
rect 14485 -3214 14543 -3199
rect 14743 -3029 14801 -3014
rect 14743 -3063 14755 -3029
rect 14789 -3063 14801 -3029
rect 14743 -3097 14801 -3063
rect 14743 -3131 14755 -3097
rect 14789 -3131 14801 -3097
rect 14743 -3165 14801 -3131
rect 14743 -3199 14755 -3165
rect 14789 -3199 14801 -3165
rect 14743 -3214 14801 -3199
rect 15001 -3029 15059 -3014
rect 15001 -3063 15013 -3029
rect 15047 -3063 15059 -3029
rect 15001 -3097 15059 -3063
rect 15001 -3131 15013 -3097
rect 15047 -3131 15059 -3097
rect 15001 -3165 15059 -3131
rect 15001 -3199 15013 -3165
rect 15047 -3199 15059 -3165
rect 15001 -3214 15059 -3199
rect 15259 -3029 15317 -3014
rect 15259 -3063 15271 -3029
rect 15305 -3063 15317 -3029
rect 15259 -3097 15317 -3063
rect 15259 -3131 15271 -3097
rect 15305 -3131 15317 -3097
rect 15259 -3165 15317 -3131
rect 15259 -3199 15271 -3165
rect 15305 -3199 15317 -3165
rect 15259 -3214 15317 -3199
rect 15517 -3029 15575 -3014
rect 15517 -3063 15529 -3029
rect 15563 -3063 15575 -3029
rect 15517 -3097 15575 -3063
rect 15517 -3131 15529 -3097
rect 15563 -3131 15575 -3097
rect 15517 -3165 15575 -3131
rect 15517 -3199 15529 -3165
rect 15563 -3199 15575 -3165
rect 15517 -3214 15575 -3199
rect 15711 -3029 15769 -3014
rect 15711 -3063 15723 -3029
rect 15757 -3063 15769 -3029
rect 15711 -3097 15769 -3063
rect 15711 -3131 15723 -3097
rect 15757 -3131 15769 -3097
rect 15711 -3165 15769 -3131
rect 15711 -3199 15723 -3165
rect 15757 -3199 15769 -3165
rect 15711 -3214 15769 -3199
rect 15969 -3029 16027 -3014
rect 15969 -3063 15981 -3029
rect 16015 -3063 16027 -3029
rect 15969 -3097 16027 -3063
rect 15969 -3131 15981 -3097
rect 16015 -3131 16027 -3097
rect 15969 -3165 16027 -3131
rect 15969 -3199 15981 -3165
rect 16015 -3199 16027 -3165
rect 15969 -3214 16027 -3199
rect 16227 -3029 16285 -3014
rect 16227 -3063 16239 -3029
rect 16273 -3063 16285 -3029
rect 16227 -3097 16285 -3063
rect 16227 -3131 16239 -3097
rect 16273 -3131 16285 -3097
rect 16227 -3165 16285 -3131
rect 16227 -3199 16239 -3165
rect 16273 -3199 16285 -3165
rect 16227 -3214 16285 -3199
rect 16485 -3029 16543 -3014
rect 16485 -3063 16497 -3029
rect 16531 -3063 16543 -3029
rect 16485 -3097 16543 -3063
rect 16485 -3131 16497 -3097
rect 16531 -3131 16543 -3097
rect 16485 -3165 16543 -3131
rect 16485 -3199 16497 -3165
rect 16531 -3199 16543 -3165
rect 16485 -3214 16543 -3199
rect 16679 -3029 16737 -3014
rect 16679 -3063 16691 -3029
rect 16725 -3063 16737 -3029
rect 16679 -3097 16737 -3063
rect 16679 -3131 16691 -3097
rect 16725 -3131 16737 -3097
rect 16679 -3165 16737 -3131
rect 16679 -3199 16691 -3165
rect 16725 -3199 16737 -3165
rect 16679 -3214 16737 -3199
rect 16937 -3029 16995 -3014
rect 16937 -3063 16949 -3029
rect 16983 -3063 16995 -3029
rect 16937 -3097 16995 -3063
rect 16937 -3131 16949 -3097
rect 16983 -3131 16995 -3097
rect 16937 -3165 16995 -3131
rect 16937 -3199 16949 -3165
rect 16983 -3199 16995 -3165
rect 16937 -3214 16995 -3199
rect 17195 -3029 17253 -3014
rect 17195 -3063 17207 -3029
rect 17241 -3063 17253 -3029
rect 17195 -3097 17253 -3063
rect 17195 -3131 17207 -3097
rect 17241 -3131 17253 -3097
rect 17195 -3165 17253 -3131
rect 17195 -3199 17207 -3165
rect 17241 -3199 17253 -3165
rect 17195 -3214 17253 -3199
rect 17453 -3029 17511 -3014
rect 17453 -3063 17465 -3029
rect 17499 -3063 17511 -3029
rect 17453 -3097 17511 -3063
rect 17453 -3131 17465 -3097
rect 17499 -3131 17511 -3097
rect 17453 -3165 17511 -3131
rect 17453 -3199 17465 -3165
rect 17499 -3199 17511 -3165
rect 17453 -3214 17511 -3199
rect 17711 -3029 17769 -3014
rect 17711 -3063 17723 -3029
rect 17757 -3063 17769 -3029
rect 17711 -3097 17769 -3063
rect 17711 -3131 17723 -3097
rect 17757 -3131 17769 -3097
rect 17711 -3165 17769 -3131
rect 17711 -3199 17723 -3165
rect 17757 -3199 17769 -3165
rect 17711 -3214 17769 -3199
rect 17905 -3029 17963 -3014
rect 17905 -3063 17917 -3029
rect 17951 -3063 17963 -3029
rect 17905 -3097 17963 -3063
rect 17905 -3131 17917 -3097
rect 17951 -3131 17963 -3097
rect 17905 -3165 17963 -3131
rect 17905 -3199 17917 -3165
rect 17951 -3199 17963 -3165
rect 17905 -3214 17963 -3199
rect 18163 -3029 18221 -3014
rect 18163 -3063 18175 -3029
rect 18209 -3063 18221 -3029
rect 18163 -3097 18221 -3063
rect 18163 -3131 18175 -3097
rect 18209 -3131 18221 -3097
rect 18163 -3165 18221 -3131
rect 18163 -3199 18175 -3165
rect 18209 -3199 18221 -3165
rect 18163 -3214 18221 -3199
rect 959 -4019 1017 -4004
rect 959 -4053 971 -4019
rect 1005 -4053 1017 -4019
rect 959 -4087 1017 -4053
rect 959 -4121 971 -4087
rect 1005 -4121 1017 -4087
rect 959 -4155 1017 -4121
rect 959 -4189 971 -4155
rect 1005 -4189 1017 -4155
rect 959 -4204 1017 -4189
rect 1217 -4019 1275 -4004
rect 1217 -4053 1229 -4019
rect 1263 -4053 1275 -4019
rect 1217 -4087 1275 -4053
rect 1217 -4121 1229 -4087
rect 1263 -4121 1275 -4087
rect 1217 -4155 1275 -4121
rect 1217 -4189 1229 -4155
rect 1263 -4189 1275 -4155
rect 1217 -4204 1275 -4189
rect 1411 -4019 1469 -4004
rect 1411 -4053 1423 -4019
rect 1457 -4053 1469 -4019
rect 1411 -4087 1469 -4053
rect 1411 -4121 1423 -4087
rect 1457 -4121 1469 -4087
rect 1411 -4155 1469 -4121
rect 1411 -4189 1423 -4155
rect 1457 -4189 1469 -4155
rect 1411 -4204 1469 -4189
rect 1669 -4019 1727 -4004
rect 1669 -4053 1681 -4019
rect 1715 -4053 1727 -4019
rect 1669 -4087 1727 -4053
rect 1669 -4121 1681 -4087
rect 1715 -4121 1727 -4087
rect 1669 -4155 1727 -4121
rect 1669 -4189 1681 -4155
rect 1715 -4189 1727 -4155
rect 1669 -4204 1727 -4189
rect 1927 -4019 1985 -4004
rect 1927 -4053 1939 -4019
rect 1973 -4053 1985 -4019
rect 1927 -4087 1985 -4053
rect 1927 -4121 1939 -4087
rect 1973 -4121 1985 -4087
rect 1927 -4155 1985 -4121
rect 1927 -4189 1939 -4155
rect 1973 -4189 1985 -4155
rect 1927 -4204 1985 -4189
rect 2185 -4019 2243 -4004
rect 2185 -4053 2197 -4019
rect 2231 -4053 2243 -4019
rect 2185 -4087 2243 -4053
rect 2185 -4121 2197 -4087
rect 2231 -4121 2243 -4087
rect 2185 -4155 2243 -4121
rect 2185 -4189 2197 -4155
rect 2231 -4189 2243 -4155
rect 2185 -4204 2243 -4189
rect 2443 -4019 2501 -4004
rect 2443 -4053 2455 -4019
rect 2489 -4053 2501 -4019
rect 2443 -4087 2501 -4053
rect 2443 -4121 2455 -4087
rect 2489 -4121 2501 -4087
rect 2443 -4155 2501 -4121
rect 2443 -4189 2455 -4155
rect 2489 -4189 2501 -4155
rect 2443 -4204 2501 -4189
rect 2637 -4019 2695 -4004
rect 2637 -4053 2649 -4019
rect 2683 -4053 2695 -4019
rect 2637 -4087 2695 -4053
rect 2637 -4121 2649 -4087
rect 2683 -4121 2695 -4087
rect 2637 -4155 2695 -4121
rect 2637 -4189 2649 -4155
rect 2683 -4189 2695 -4155
rect 2637 -4204 2695 -4189
rect 2895 -4019 2953 -4004
rect 2895 -4053 2907 -4019
rect 2941 -4053 2953 -4019
rect 2895 -4087 2953 -4053
rect 2895 -4121 2907 -4087
rect 2941 -4121 2953 -4087
rect 2895 -4155 2953 -4121
rect 2895 -4189 2907 -4155
rect 2941 -4189 2953 -4155
rect 2895 -4204 2953 -4189
rect 3153 -4019 3211 -4004
rect 3153 -4053 3165 -4019
rect 3199 -4053 3211 -4019
rect 3153 -4087 3211 -4053
rect 3153 -4121 3165 -4087
rect 3199 -4121 3211 -4087
rect 3153 -4155 3211 -4121
rect 3153 -4189 3165 -4155
rect 3199 -4189 3211 -4155
rect 3153 -4204 3211 -4189
rect 3411 -4019 3469 -4004
rect 3411 -4053 3423 -4019
rect 3457 -4053 3469 -4019
rect 3411 -4087 3469 -4053
rect 3411 -4121 3423 -4087
rect 3457 -4121 3469 -4087
rect 3411 -4155 3469 -4121
rect 3411 -4189 3423 -4155
rect 3457 -4189 3469 -4155
rect 3411 -4204 3469 -4189
rect 3605 -4019 3663 -4004
rect 3605 -4053 3617 -4019
rect 3651 -4053 3663 -4019
rect 3605 -4087 3663 -4053
rect 3605 -4121 3617 -4087
rect 3651 -4121 3663 -4087
rect 3605 -4155 3663 -4121
rect 3605 -4189 3617 -4155
rect 3651 -4189 3663 -4155
rect 3605 -4204 3663 -4189
rect 3863 -4019 3921 -4004
rect 3863 -4053 3875 -4019
rect 3909 -4053 3921 -4019
rect 3863 -4087 3921 -4053
rect 3863 -4121 3875 -4087
rect 3909 -4121 3921 -4087
rect 3863 -4155 3921 -4121
rect 3863 -4189 3875 -4155
rect 3909 -4189 3921 -4155
rect 3863 -4204 3921 -4189
rect 4121 -4019 4179 -4004
rect 4121 -4053 4133 -4019
rect 4167 -4053 4179 -4019
rect 4121 -4087 4179 -4053
rect 4121 -4121 4133 -4087
rect 4167 -4121 4179 -4087
rect 4121 -4155 4179 -4121
rect 4121 -4189 4133 -4155
rect 4167 -4189 4179 -4155
rect 4121 -4204 4179 -4189
rect 4379 -4019 4437 -4004
rect 4379 -4053 4391 -4019
rect 4425 -4053 4437 -4019
rect 4379 -4087 4437 -4053
rect 4379 -4121 4391 -4087
rect 4425 -4121 4437 -4087
rect 4379 -4155 4437 -4121
rect 4379 -4189 4391 -4155
rect 4425 -4189 4437 -4155
rect 4379 -4204 4437 -4189
rect 4637 -4019 4695 -4004
rect 4637 -4053 4649 -4019
rect 4683 -4053 4695 -4019
rect 4637 -4087 4695 -4053
rect 4637 -4121 4649 -4087
rect 4683 -4121 4695 -4087
rect 4637 -4155 4695 -4121
rect 4637 -4189 4649 -4155
rect 4683 -4189 4695 -4155
rect 4637 -4204 4695 -4189
rect 4830 -4019 4888 -4004
rect 4830 -4053 4842 -4019
rect 4876 -4053 4888 -4019
rect 4830 -4087 4888 -4053
rect 4830 -4121 4842 -4087
rect 4876 -4121 4888 -4087
rect 4830 -4155 4888 -4121
rect 4830 -4189 4842 -4155
rect 4876 -4189 4888 -4155
rect 4830 -4204 4888 -4189
rect 5088 -4019 5146 -4004
rect 5088 -4053 5100 -4019
rect 5134 -4053 5146 -4019
rect 5088 -4087 5146 -4053
rect 5088 -4121 5100 -4087
rect 5134 -4121 5146 -4087
rect 5088 -4155 5146 -4121
rect 5088 -4189 5100 -4155
rect 5134 -4189 5146 -4155
rect 5088 -4204 5146 -4189
rect 5316 -4019 5374 -4004
rect 5316 -4053 5328 -4019
rect 5362 -4053 5374 -4019
rect 5316 -4087 5374 -4053
rect 5316 -4121 5328 -4087
rect 5362 -4121 5374 -4087
rect 5316 -4155 5374 -4121
rect 5316 -4189 5328 -4155
rect 5362 -4189 5374 -4155
rect 5316 -4204 5374 -4189
rect 5574 -4019 5632 -4004
rect 5574 -4053 5586 -4019
rect 5620 -4053 5632 -4019
rect 5574 -4087 5632 -4053
rect 5574 -4121 5586 -4087
rect 5620 -4121 5632 -4087
rect 5574 -4155 5632 -4121
rect 5574 -4189 5586 -4155
rect 5620 -4189 5632 -4155
rect 5574 -4204 5632 -4189
rect 5768 -4019 5826 -4004
rect 5768 -4053 5780 -4019
rect 5814 -4053 5826 -4019
rect 5768 -4087 5826 -4053
rect 5768 -4121 5780 -4087
rect 5814 -4121 5826 -4087
rect 5768 -4155 5826 -4121
rect 5768 -4189 5780 -4155
rect 5814 -4189 5826 -4155
rect 5768 -4204 5826 -4189
rect 6026 -4019 6084 -4004
rect 6026 -4053 6038 -4019
rect 6072 -4053 6084 -4019
rect 6026 -4087 6084 -4053
rect 6026 -4121 6038 -4087
rect 6072 -4121 6084 -4087
rect 6026 -4155 6084 -4121
rect 6026 -4189 6038 -4155
rect 6072 -4189 6084 -4155
rect 6026 -4204 6084 -4189
rect 6284 -4019 6342 -4004
rect 6284 -4053 6296 -4019
rect 6330 -4053 6342 -4019
rect 6284 -4087 6342 -4053
rect 6284 -4121 6296 -4087
rect 6330 -4121 6342 -4087
rect 6284 -4155 6342 -4121
rect 6284 -4189 6296 -4155
rect 6330 -4189 6342 -4155
rect 6284 -4204 6342 -4189
rect 6542 -4019 6600 -4004
rect 6542 -4053 6554 -4019
rect 6588 -4053 6600 -4019
rect 6542 -4087 6600 -4053
rect 6542 -4121 6554 -4087
rect 6588 -4121 6600 -4087
rect 6542 -4155 6600 -4121
rect 6542 -4189 6554 -4155
rect 6588 -4189 6600 -4155
rect 6542 -4204 6600 -4189
rect 6800 -4019 6858 -4004
rect 6800 -4053 6812 -4019
rect 6846 -4053 6858 -4019
rect 6800 -4087 6858 -4053
rect 6800 -4121 6812 -4087
rect 6846 -4121 6858 -4087
rect 6800 -4155 6858 -4121
rect 6800 -4189 6812 -4155
rect 6846 -4189 6858 -4155
rect 6800 -4204 6858 -4189
rect 6994 -4019 7052 -4004
rect 6994 -4053 7006 -4019
rect 7040 -4053 7052 -4019
rect 6994 -4087 7052 -4053
rect 6994 -4121 7006 -4087
rect 7040 -4121 7052 -4087
rect 6994 -4155 7052 -4121
rect 6994 -4189 7006 -4155
rect 7040 -4189 7052 -4155
rect 6994 -4204 7052 -4189
rect 7252 -4019 7310 -4004
rect 7252 -4053 7264 -4019
rect 7298 -4053 7310 -4019
rect 7252 -4087 7310 -4053
rect 7252 -4121 7264 -4087
rect 7298 -4121 7310 -4087
rect 7252 -4155 7310 -4121
rect 7252 -4189 7264 -4155
rect 7298 -4189 7310 -4155
rect 7252 -4204 7310 -4189
rect 7510 -4019 7568 -4004
rect 7510 -4053 7522 -4019
rect 7556 -4053 7568 -4019
rect 7510 -4087 7568 -4053
rect 7510 -4121 7522 -4087
rect 7556 -4121 7568 -4087
rect 7510 -4155 7568 -4121
rect 7510 -4189 7522 -4155
rect 7556 -4189 7568 -4155
rect 7510 -4204 7568 -4189
rect 7768 -4019 7826 -4004
rect 7768 -4053 7780 -4019
rect 7814 -4053 7826 -4019
rect 7768 -4087 7826 -4053
rect 7768 -4121 7780 -4087
rect 7814 -4121 7826 -4087
rect 7768 -4155 7826 -4121
rect 7768 -4189 7780 -4155
rect 7814 -4189 7826 -4155
rect 7768 -4204 7826 -4189
rect 7962 -4019 8020 -4004
rect 7962 -4053 7974 -4019
rect 8008 -4053 8020 -4019
rect 7962 -4087 8020 -4053
rect 7962 -4121 7974 -4087
rect 8008 -4121 8020 -4087
rect 7962 -4155 8020 -4121
rect 7962 -4189 7974 -4155
rect 8008 -4189 8020 -4155
rect 7962 -4204 8020 -4189
rect 8220 -4019 8278 -4004
rect 8220 -4053 8232 -4019
rect 8266 -4053 8278 -4019
rect 8220 -4087 8278 -4053
rect 8220 -4121 8232 -4087
rect 8266 -4121 8278 -4087
rect 8220 -4155 8278 -4121
rect 8220 -4189 8232 -4155
rect 8266 -4189 8278 -4155
rect 8220 -4204 8278 -4189
rect 8478 -4019 8536 -4004
rect 8478 -4053 8490 -4019
rect 8524 -4053 8536 -4019
rect 8478 -4087 8536 -4053
rect 8478 -4121 8490 -4087
rect 8524 -4121 8536 -4087
rect 8478 -4155 8536 -4121
rect 8478 -4189 8490 -4155
rect 8524 -4189 8536 -4155
rect 8478 -4204 8536 -4189
rect 8736 -4019 8794 -4004
rect 8736 -4053 8748 -4019
rect 8782 -4053 8794 -4019
rect 8736 -4087 8794 -4053
rect 8736 -4121 8748 -4087
rect 8782 -4121 8794 -4087
rect 8736 -4155 8794 -4121
rect 8736 -4189 8748 -4155
rect 8782 -4189 8794 -4155
rect 8736 -4204 8794 -4189
rect 8994 -4019 9052 -4004
rect 8994 -4053 9006 -4019
rect 9040 -4053 9052 -4019
rect 8994 -4087 9052 -4053
rect 8994 -4121 9006 -4087
rect 9040 -4121 9052 -4087
rect 8994 -4155 9052 -4121
rect 8994 -4189 9006 -4155
rect 9040 -4189 9052 -4155
rect 8994 -4204 9052 -4189
rect 9188 -4019 9246 -4004
rect 9188 -4053 9200 -4019
rect 9234 -4053 9246 -4019
rect 9188 -4087 9246 -4053
rect 9188 -4121 9200 -4087
rect 9234 -4121 9246 -4087
rect 9188 -4155 9246 -4121
rect 9188 -4189 9200 -4155
rect 9234 -4189 9246 -4155
rect 9188 -4204 9246 -4189
rect 9446 -4019 9504 -4004
rect 9446 -4053 9458 -4019
rect 9492 -4053 9504 -4019
rect 9446 -4087 9504 -4053
rect 9446 -4121 9458 -4087
rect 9492 -4121 9504 -4087
rect 9446 -4155 9504 -4121
rect 9446 -4189 9458 -4155
rect 9492 -4189 9504 -4155
rect 9446 -4204 9504 -4189
rect 9676 -4019 9734 -4004
rect 9676 -4053 9688 -4019
rect 9722 -4053 9734 -4019
rect 9676 -4087 9734 -4053
rect 9676 -4121 9688 -4087
rect 9722 -4121 9734 -4087
rect 9676 -4155 9734 -4121
rect 9676 -4189 9688 -4155
rect 9722 -4189 9734 -4155
rect 9676 -4204 9734 -4189
rect 9934 -4019 9992 -4004
rect 9934 -4053 9946 -4019
rect 9980 -4053 9992 -4019
rect 9934 -4087 9992 -4053
rect 9934 -4121 9946 -4087
rect 9980 -4121 9992 -4087
rect 9934 -4155 9992 -4121
rect 9934 -4189 9946 -4155
rect 9980 -4189 9992 -4155
rect 9934 -4204 9992 -4189
rect 10128 -4019 10186 -4004
rect 10128 -4053 10140 -4019
rect 10174 -4053 10186 -4019
rect 10128 -4087 10186 -4053
rect 10128 -4121 10140 -4087
rect 10174 -4121 10186 -4087
rect 10128 -4155 10186 -4121
rect 10128 -4189 10140 -4155
rect 10174 -4189 10186 -4155
rect 10128 -4204 10186 -4189
rect 10386 -4019 10444 -4004
rect 10386 -4053 10398 -4019
rect 10432 -4053 10444 -4019
rect 10386 -4087 10444 -4053
rect 10386 -4121 10398 -4087
rect 10432 -4121 10444 -4087
rect 10386 -4155 10444 -4121
rect 10386 -4189 10398 -4155
rect 10432 -4189 10444 -4155
rect 10386 -4204 10444 -4189
rect 10644 -4019 10702 -4004
rect 10644 -4053 10656 -4019
rect 10690 -4053 10702 -4019
rect 10644 -4087 10702 -4053
rect 10644 -4121 10656 -4087
rect 10690 -4121 10702 -4087
rect 10644 -4155 10702 -4121
rect 10644 -4189 10656 -4155
rect 10690 -4189 10702 -4155
rect 10644 -4204 10702 -4189
rect 10902 -4019 10960 -4004
rect 10902 -4053 10914 -4019
rect 10948 -4053 10960 -4019
rect 10902 -4087 10960 -4053
rect 10902 -4121 10914 -4087
rect 10948 -4121 10960 -4087
rect 10902 -4155 10960 -4121
rect 10902 -4189 10914 -4155
rect 10948 -4189 10960 -4155
rect 10902 -4204 10960 -4189
rect 11160 -4019 11218 -4004
rect 11160 -4053 11172 -4019
rect 11206 -4053 11218 -4019
rect 11160 -4087 11218 -4053
rect 11160 -4121 11172 -4087
rect 11206 -4121 11218 -4087
rect 11160 -4155 11218 -4121
rect 11160 -4189 11172 -4155
rect 11206 -4189 11218 -4155
rect 11160 -4204 11218 -4189
rect 11354 -4019 11412 -4004
rect 11354 -4053 11366 -4019
rect 11400 -4053 11412 -4019
rect 11354 -4087 11412 -4053
rect 11354 -4121 11366 -4087
rect 11400 -4121 11412 -4087
rect 11354 -4155 11412 -4121
rect 11354 -4189 11366 -4155
rect 11400 -4189 11412 -4155
rect 11354 -4204 11412 -4189
rect 11612 -4019 11670 -4004
rect 11612 -4053 11624 -4019
rect 11658 -4053 11670 -4019
rect 11612 -4087 11670 -4053
rect 11612 -4121 11624 -4087
rect 11658 -4121 11670 -4087
rect 11612 -4155 11670 -4121
rect 11612 -4189 11624 -4155
rect 11658 -4189 11670 -4155
rect 11612 -4204 11670 -4189
rect 11870 -4019 11928 -4004
rect 11870 -4053 11882 -4019
rect 11916 -4053 11928 -4019
rect 11870 -4087 11928 -4053
rect 11870 -4121 11882 -4087
rect 11916 -4121 11928 -4087
rect 11870 -4155 11928 -4121
rect 11870 -4189 11882 -4155
rect 11916 -4189 11928 -4155
rect 11870 -4204 11928 -4189
rect 12128 -4019 12186 -4004
rect 12128 -4053 12140 -4019
rect 12174 -4053 12186 -4019
rect 12128 -4087 12186 -4053
rect 12128 -4121 12140 -4087
rect 12174 -4121 12186 -4087
rect 12128 -4155 12186 -4121
rect 12128 -4189 12140 -4155
rect 12174 -4189 12186 -4155
rect 12128 -4204 12186 -4189
rect 12322 -4019 12380 -4004
rect 12322 -4053 12334 -4019
rect 12368 -4053 12380 -4019
rect 12322 -4087 12380 -4053
rect 12322 -4121 12334 -4087
rect 12368 -4121 12380 -4087
rect 12322 -4155 12380 -4121
rect 12322 -4189 12334 -4155
rect 12368 -4189 12380 -4155
rect 12322 -4204 12380 -4189
rect 12580 -4019 12638 -4004
rect 12580 -4053 12592 -4019
rect 12626 -4053 12638 -4019
rect 12580 -4087 12638 -4053
rect 12580 -4121 12592 -4087
rect 12626 -4121 12638 -4087
rect 12580 -4155 12638 -4121
rect 12580 -4189 12592 -4155
rect 12626 -4189 12638 -4155
rect 12580 -4204 12638 -4189
rect 12838 -4019 12896 -4004
rect 12838 -4053 12850 -4019
rect 12884 -4053 12896 -4019
rect 12838 -4087 12896 -4053
rect 12838 -4121 12850 -4087
rect 12884 -4121 12896 -4087
rect 12838 -4155 12896 -4121
rect 12838 -4189 12850 -4155
rect 12884 -4189 12896 -4155
rect 12838 -4204 12896 -4189
rect 13096 -4019 13154 -4004
rect 13096 -4053 13108 -4019
rect 13142 -4053 13154 -4019
rect 13096 -4087 13154 -4053
rect 13096 -4121 13108 -4087
rect 13142 -4121 13154 -4087
rect 13096 -4155 13154 -4121
rect 13096 -4189 13108 -4155
rect 13142 -4189 13154 -4155
rect 13096 -4204 13154 -4189
rect 13354 -4019 13412 -4004
rect 13354 -4053 13366 -4019
rect 13400 -4053 13412 -4019
rect 13354 -4087 13412 -4053
rect 13354 -4121 13366 -4087
rect 13400 -4121 13412 -4087
rect 13354 -4155 13412 -4121
rect 13354 -4189 13366 -4155
rect 13400 -4189 13412 -4155
rect 13354 -4204 13412 -4189
rect 13548 -4019 13606 -4004
rect 13548 -4053 13560 -4019
rect 13594 -4053 13606 -4019
rect 13548 -4087 13606 -4053
rect 13548 -4121 13560 -4087
rect 13594 -4121 13606 -4087
rect 13548 -4155 13606 -4121
rect 13548 -4189 13560 -4155
rect 13594 -4189 13606 -4155
rect 13548 -4204 13606 -4189
rect 13806 -4019 13864 -4004
rect 13806 -4053 13818 -4019
rect 13852 -4053 13864 -4019
rect 13806 -4087 13864 -4053
rect 13806 -4121 13818 -4087
rect 13852 -4121 13864 -4087
rect 13806 -4155 13864 -4121
rect 13806 -4189 13818 -4155
rect 13852 -4189 13864 -4155
rect 13806 -4204 13864 -4189
rect 14034 -4019 14092 -4004
rect 14034 -4053 14046 -4019
rect 14080 -4053 14092 -4019
rect 14034 -4087 14092 -4053
rect 14034 -4121 14046 -4087
rect 14080 -4121 14092 -4087
rect 14034 -4155 14092 -4121
rect 14034 -4189 14046 -4155
rect 14080 -4189 14092 -4155
rect 14034 -4204 14092 -4189
rect 14292 -4019 14350 -4004
rect 14292 -4053 14304 -4019
rect 14338 -4053 14350 -4019
rect 14292 -4087 14350 -4053
rect 14292 -4121 14304 -4087
rect 14338 -4121 14350 -4087
rect 14292 -4155 14350 -4121
rect 14292 -4189 14304 -4155
rect 14338 -4189 14350 -4155
rect 14292 -4204 14350 -4189
rect 14485 -4019 14543 -4004
rect 14485 -4053 14497 -4019
rect 14531 -4053 14543 -4019
rect 14485 -4087 14543 -4053
rect 14485 -4121 14497 -4087
rect 14531 -4121 14543 -4087
rect 14485 -4155 14543 -4121
rect 14485 -4189 14497 -4155
rect 14531 -4189 14543 -4155
rect 14485 -4204 14543 -4189
rect 14743 -4019 14801 -4004
rect 14743 -4053 14755 -4019
rect 14789 -4053 14801 -4019
rect 14743 -4087 14801 -4053
rect 14743 -4121 14755 -4087
rect 14789 -4121 14801 -4087
rect 14743 -4155 14801 -4121
rect 14743 -4189 14755 -4155
rect 14789 -4189 14801 -4155
rect 14743 -4204 14801 -4189
rect 15001 -4019 15059 -4004
rect 15001 -4053 15013 -4019
rect 15047 -4053 15059 -4019
rect 15001 -4087 15059 -4053
rect 15001 -4121 15013 -4087
rect 15047 -4121 15059 -4087
rect 15001 -4155 15059 -4121
rect 15001 -4189 15013 -4155
rect 15047 -4189 15059 -4155
rect 15001 -4204 15059 -4189
rect 15259 -4019 15317 -4004
rect 15259 -4053 15271 -4019
rect 15305 -4053 15317 -4019
rect 15259 -4087 15317 -4053
rect 15259 -4121 15271 -4087
rect 15305 -4121 15317 -4087
rect 15259 -4155 15317 -4121
rect 15259 -4189 15271 -4155
rect 15305 -4189 15317 -4155
rect 15259 -4204 15317 -4189
rect 15517 -4019 15575 -4004
rect 15517 -4053 15529 -4019
rect 15563 -4053 15575 -4019
rect 15517 -4087 15575 -4053
rect 15517 -4121 15529 -4087
rect 15563 -4121 15575 -4087
rect 15517 -4155 15575 -4121
rect 15517 -4189 15529 -4155
rect 15563 -4189 15575 -4155
rect 15517 -4204 15575 -4189
rect 15711 -4019 15769 -4004
rect 15711 -4053 15723 -4019
rect 15757 -4053 15769 -4019
rect 15711 -4087 15769 -4053
rect 15711 -4121 15723 -4087
rect 15757 -4121 15769 -4087
rect 15711 -4155 15769 -4121
rect 15711 -4189 15723 -4155
rect 15757 -4189 15769 -4155
rect 15711 -4204 15769 -4189
rect 15969 -4019 16027 -4004
rect 15969 -4053 15981 -4019
rect 16015 -4053 16027 -4019
rect 15969 -4087 16027 -4053
rect 15969 -4121 15981 -4087
rect 16015 -4121 16027 -4087
rect 15969 -4155 16027 -4121
rect 15969 -4189 15981 -4155
rect 16015 -4189 16027 -4155
rect 15969 -4204 16027 -4189
rect 16227 -4019 16285 -4004
rect 16227 -4053 16239 -4019
rect 16273 -4053 16285 -4019
rect 16227 -4087 16285 -4053
rect 16227 -4121 16239 -4087
rect 16273 -4121 16285 -4087
rect 16227 -4155 16285 -4121
rect 16227 -4189 16239 -4155
rect 16273 -4189 16285 -4155
rect 16227 -4204 16285 -4189
rect 16485 -4019 16543 -4004
rect 16485 -4053 16497 -4019
rect 16531 -4053 16543 -4019
rect 16485 -4087 16543 -4053
rect 16485 -4121 16497 -4087
rect 16531 -4121 16543 -4087
rect 16485 -4155 16543 -4121
rect 16485 -4189 16497 -4155
rect 16531 -4189 16543 -4155
rect 16485 -4204 16543 -4189
rect 16679 -4019 16737 -4004
rect 16679 -4053 16691 -4019
rect 16725 -4053 16737 -4019
rect 16679 -4087 16737 -4053
rect 16679 -4121 16691 -4087
rect 16725 -4121 16737 -4087
rect 16679 -4155 16737 -4121
rect 16679 -4189 16691 -4155
rect 16725 -4189 16737 -4155
rect 16679 -4204 16737 -4189
rect 16937 -4019 16995 -4004
rect 16937 -4053 16949 -4019
rect 16983 -4053 16995 -4019
rect 16937 -4087 16995 -4053
rect 16937 -4121 16949 -4087
rect 16983 -4121 16995 -4087
rect 16937 -4155 16995 -4121
rect 16937 -4189 16949 -4155
rect 16983 -4189 16995 -4155
rect 16937 -4204 16995 -4189
rect 17195 -4019 17253 -4004
rect 17195 -4053 17207 -4019
rect 17241 -4053 17253 -4019
rect 17195 -4087 17253 -4053
rect 17195 -4121 17207 -4087
rect 17241 -4121 17253 -4087
rect 17195 -4155 17253 -4121
rect 17195 -4189 17207 -4155
rect 17241 -4189 17253 -4155
rect 17195 -4204 17253 -4189
rect 17453 -4019 17511 -4004
rect 17453 -4053 17465 -4019
rect 17499 -4053 17511 -4019
rect 17453 -4087 17511 -4053
rect 17453 -4121 17465 -4087
rect 17499 -4121 17511 -4087
rect 17453 -4155 17511 -4121
rect 17453 -4189 17465 -4155
rect 17499 -4189 17511 -4155
rect 17453 -4204 17511 -4189
rect 17711 -4019 17769 -4004
rect 17711 -4053 17723 -4019
rect 17757 -4053 17769 -4019
rect 17711 -4087 17769 -4053
rect 17711 -4121 17723 -4087
rect 17757 -4121 17769 -4087
rect 17711 -4155 17769 -4121
rect 17711 -4189 17723 -4155
rect 17757 -4189 17769 -4155
rect 17711 -4204 17769 -4189
rect 17905 -4019 17963 -4004
rect 17905 -4053 17917 -4019
rect 17951 -4053 17963 -4019
rect 17905 -4087 17963 -4053
rect 17905 -4121 17917 -4087
rect 17951 -4121 17963 -4087
rect 17905 -4155 17963 -4121
rect 17905 -4189 17917 -4155
rect 17951 -4189 17963 -4155
rect 17905 -4204 17963 -4189
rect 18163 -4019 18221 -4004
rect 18163 -4053 18175 -4019
rect 18209 -4053 18221 -4019
rect 18163 -4087 18221 -4053
rect 18163 -4121 18175 -4087
rect 18209 -4121 18221 -4087
rect 18163 -4155 18221 -4121
rect 18163 -4189 18175 -4155
rect 18209 -4189 18221 -4155
rect 18163 -4204 18221 -4189
rect 959 -4575 1017 -4560
rect 959 -4609 971 -4575
rect 1005 -4609 1017 -4575
rect 959 -4643 1017 -4609
rect 959 -4677 971 -4643
rect 1005 -4677 1017 -4643
rect 959 -4711 1017 -4677
rect 959 -4745 971 -4711
rect 1005 -4745 1017 -4711
rect 959 -4760 1017 -4745
rect 1217 -4575 1275 -4560
rect 1217 -4609 1229 -4575
rect 1263 -4609 1275 -4575
rect 1217 -4643 1275 -4609
rect 1217 -4677 1229 -4643
rect 1263 -4677 1275 -4643
rect 1217 -4711 1275 -4677
rect 1217 -4745 1229 -4711
rect 1263 -4745 1275 -4711
rect 1217 -4760 1275 -4745
rect 1411 -4575 1469 -4560
rect 1411 -4609 1423 -4575
rect 1457 -4609 1469 -4575
rect 1411 -4643 1469 -4609
rect 1411 -4677 1423 -4643
rect 1457 -4677 1469 -4643
rect 1411 -4711 1469 -4677
rect 1411 -4745 1423 -4711
rect 1457 -4745 1469 -4711
rect 1411 -4760 1469 -4745
rect 1669 -4575 1727 -4560
rect 1669 -4609 1681 -4575
rect 1715 -4609 1727 -4575
rect 1669 -4643 1727 -4609
rect 1669 -4677 1681 -4643
rect 1715 -4677 1727 -4643
rect 1669 -4711 1727 -4677
rect 1669 -4745 1681 -4711
rect 1715 -4745 1727 -4711
rect 1669 -4760 1727 -4745
rect 1927 -4575 1985 -4560
rect 1927 -4609 1939 -4575
rect 1973 -4609 1985 -4575
rect 1927 -4643 1985 -4609
rect 1927 -4677 1939 -4643
rect 1973 -4677 1985 -4643
rect 1927 -4711 1985 -4677
rect 1927 -4745 1939 -4711
rect 1973 -4745 1985 -4711
rect 1927 -4760 1985 -4745
rect 2185 -4575 2243 -4560
rect 2185 -4609 2197 -4575
rect 2231 -4609 2243 -4575
rect 2185 -4643 2243 -4609
rect 2185 -4677 2197 -4643
rect 2231 -4677 2243 -4643
rect 2185 -4711 2243 -4677
rect 2185 -4745 2197 -4711
rect 2231 -4745 2243 -4711
rect 2185 -4760 2243 -4745
rect 2443 -4575 2501 -4560
rect 2443 -4609 2455 -4575
rect 2489 -4609 2501 -4575
rect 2443 -4643 2501 -4609
rect 2443 -4677 2455 -4643
rect 2489 -4677 2501 -4643
rect 2443 -4711 2501 -4677
rect 2443 -4745 2455 -4711
rect 2489 -4745 2501 -4711
rect 2443 -4760 2501 -4745
rect 2637 -4575 2695 -4560
rect 2637 -4609 2649 -4575
rect 2683 -4609 2695 -4575
rect 2637 -4643 2695 -4609
rect 2637 -4677 2649 -4643
rect 2683 -4677 2695 -4643
rect 2637 -4711 2695 -4677
rect 2637 -4745 2649 -4711
rect 2683 -4745 2695 -4711
rect 2637 -4760 2695 -4745
rect 2895 -4575 2953 -4560
rect 2895 -4609 2907 -4575
rect 2941 -4609 2953 -4575
rect 2895 -4643 2953 -4609
rect 2895 -4677 2907 -4643
rect 2941 -4677 2953 -4643
rect 2895 -4711 2953 -4677
rect 2895 -4745 2907 -4711
rect 2941 -4745 2953 -4711
rect 2895 -4760 2953 -4745
rect 3153 -4575 3211 -4560
rect 3153 -4609 3165 -4575
rect 3199 -4609 3211 -4575
rect 3153 -4643 3211 -4609
rect 3153 -4677 3165 -4643
rect 3199 -4677 3211 -4643
rect 3153 -4711 3211 -4677
rect 3153 -4745 3165 -4711
rect 3199 -4745 3211 -4711
rect 3153 -4760 3211 -4745
rect 3411 -4575 3469 -4560
rect 3411 -4609 3423 -4575
rect 3457 -4609 3469 -4575
rect 3411 -4643 3469 -4609
rect 3411 -4677 3423 -4643
rect 3457 -4677 3469 -4643
rect 3411 -4711 3469 -4677
rect 3411 -4745 3423 -4711
rect 3457 -4745 3469 -4711
rect 3411 -4760 3469 -4745
rect 3605 -4575 3663 -4560
rect 3605 -4609 3617 -4575
rect 3651 -4609 3663 -4575
rect 3605 -4643 3663 -4609
rect 3605 -4677 3617 -4643
rect 3651 -4677 3663 -4643
rect 3605 -4711 3663 -4677
rect 3605 -4745 3617 -4711
rect 3651 -4745 3663 -4711
rect 3605 -4760 3663 -4745
rect 3863 -4575 3921 -4560
rect 3863 -4609 3875 -4575
rect 3909 -4609 3921 -4575
rect 3863 -4643 3921 -4609
rect 3863 -4677 3875 -4643
rect 3909 -4677 3921 -4643
rect 3863 -4711 3921 -4677
rect 3863 -4745 3875 -4711
rect 3909 -4745 3921 -4711
rect 3863 -4760 3921 -4745
rect 4121 -4575 4179 -4560
rect 4121 -4609 4133 -4575
rect 4167 -4609 4179 -4575
rect 4121 -4643 4179 -4609
rect 4121 -4677 4133 -4643
rect 4167 -4677 4179 -4643
rect 4121 -4711 4179 -4677
rect 4121 -4745 4133 -4711
rect 4167 -4745 4179 -4711
rect 4121 -4760 4179 -4745
rect 4379 -4575 4437 -4560
rect 4379 -4609 4391 -4575
rect 4425 -4609 4437 -4575
rect 4379 -4643 4437 -4609
rect 4379 -4677 4391 -4643
rect 4425 -4677 4437 -4643
rect 4379 -4711 4437 -4677
rect 4379 -4745 4391 -4711
rect 4425 -4745 4437 -4711
rect 4379 -4760 4437 -4745
rect 4637 -4575 4695 -4560
rect 4637 -4609 4649 -4575
rect 4683 -4609 4695 -4575
rect 4637 -4643 4695 -4609
rect 4637 -4677 4649 -4643
rect 4683 -4677 4695 -4643
rect 4637 -4711 4695 -4677
rect 4637 -4745 4649 -4711
rect 4683 -4745 4695 -4711
rect 4637 -4760 4695 -4745
rect 4830 -4575 4888 -4560
rect 4830 -4609 4842 -4575
rect 4876 -4609 4888 -4575
rect 4830 -4643 4888 -4609
rect 4830 -4677 4842 -4643
rect 4876 -4677 4888 -4643
rect 4830 -4711 4888 -4677
rect 4830 -4745 4842 -4711
rect 4876 -4745 4888 -4711
rect 4830 -4760 4888 -4745
rect 5088 -4575 5146 -4560
rect 5088 -4609 5100 -4575
rect 5134 -4609 5146 -4575
rect 5088 -4643 5146 -4609
rect 5088 -4677 5100 -4643
rect 5134 -4677 5146 -4643
rect 5088 -4711 5146 -4677
rect 5088 -4745 5100 -4711
rect 5134 -4745 5146 -4711
rect 5088 -4760 5146 -4745
rect 5316 -4575 5374 -4560
rect 5316 -4609 5328 -4575
rect 5362 -4609 5374 -4575
rect 5316 -4643 5374 -4609
rect 5316 -4677 5328 -4643
rect 5362 -4677 5374 -4643
rect 5316 -4711 5374 -4677
rect 5316 -4745 5328 -4711
rect 5362 -4745 5374 -4711
rect 5316 -4760 5374 -4745
rect 5574 -4575 5632 -4560
rect 5574 -4609 5586 -4575
rect 5620 -4609 5632 -4575
rect 5574 -4643 5632 -4609
rect 5574 -4677 5586 -4643
rect 5620 -4677 5632 -4643
rect 5574 -4711 5632 -4677
rect 5574 -4745 5586 -4711
rect 5620 -4745 5632 -4711
rect 5574 -4760 5632 -4745
rect 5768 -4575 5826 -4560
rect 5768 -4609 5780 -4575
rect 5814 -4609 5826 -4575
rect 5768 -4643 5826 -4609
rect 5768 -4677 5780 -4643
rect 5814 -4677 5826 -4643
rect 5768 -4711 5826 -4677
rect 5768 -4745 5780 -4711
rect 5814 -4745 5826 -4711
rect 5768 -4760 5826 -4745
rect 6026 -4575 6084 -4560
rect 6026 -4609 6038 -4575
rect 6072 -4609 6084 -4575
rect 6026 -4643 6084 -4609
rect 6026 -4677 6038 -4643
rect 6072 -4677 6084 -4643
rect 6026 -4711 6084 -4677
rect 6026 -4745 6038 -4711
rect 6072 -4745 6084 -4711
rect 6026 -4760 6084 -4745
rect 6284 -4575 6342 -4560
rect 6284 -4609 6296 -4575
rect 6330 -4609 6342 -4575
rect 6284 -4643 6342 -4609
rect 6284 -4677 6296 -4643
rect 6330 -4677 6342 -4643
rect 6284 -4711 6342 -4677
rect 6284 -4745 6296 -4711
rect 6330 -4745 6342 -4711
rect 6284 -4760 6342 -4745
rect 6542 -4575 6600 -4560
rect 6542 -4609 6554 -4575
rect 6588 -4609 6600 -4575
rect 6542 -4643 6600 -4609
rect 6542 -4677 6554 -4643
rect 6588 -4677 6600 -4643
rect 6542 -4711 6600 -4677
rect 6542 -4745 6554 -4711
rect 6588 -4745 6600 -4711
rect 6542 -4760 6600 -4745
rect 6800 -4575 6858 -4560
rect 6800 -4609 6812 -4575
rect 6846 -4609 6858 -4575
rect 6800 -4643 6858 -4609
rect 6800 -4677 6812 -4643
rect 6846 -4677 6858 -4643
rect 6800 -4711 6858 -4677
rect 6800 -4745 6812 -4711
rect 6846 -4745 6858 -4711
rect 6800 -4760 6858 -4745
rect 6994 -4575 7052 -4560
rect 6994 -4609 7006 -4575
rect 7040 -4609 7052 -4575
rect 6994 -4643 7052 -4609
rect 6994 -4677 7006 -4643
rect 7040 -4677 7052 -4643
rect 6994 -4711 7052 -4677
rect 6994 -4745 7006 -4711
rect 7040 -4745 7052 -4711
rect 6994 -4760 7052 -4745
rect 7252 -4575 7310 -4560
rect 7252 -4609 7264 -4575
rect 7298 -4609 7310 -4575
rect 7252 -4643 7310 -4609
rect 7252 -4677 7264 -4643
rect 7298 -4677 7310 -4643
rect 7252 -4711 7310 -4677
rect 7252 -4745 7264 -4711
rect 7298 -4745 7310 -4711
rect 7252 -4760 7310 -4745
rect 7510 -4575 7568 -4560
rect 7510 -4609 7522 -4575
rect 7556 -4609 7568 -4575
rect 7510 -4643 7568 -4609
rect 7510 -4677 7522 -4643
rect 7556 -4677 7568 -4643
rect 7510 -4711 7568 -4677
rect 7510 -4745 7522 -4711
rect 7556 -4745 7568 -4711
rect 7510 -4760 7568 -4745
rect 7768 -4575 7826 -4560
rect 7768 -4609 7780 -4575
rect 7814 -4609 7826 -4575
rect 7768 -4643 7826 -4609
rect 7768 -4677 7780 -4643
rect 7814 -4677 7826 -4643
rect 7768 -4711 7826 -4677
rect 7768 -4745 7780 -4711
rect 7814 -4745 7826 -4711
rect 7768 -4760 7826 -4745
rect 7962 -4575 8020 -4560
rect 7962 -4609 7974 -4575
rect 8008 -4609 8020 -4575
rect 7962 -4643 8020 -4609
rect 7962 -4677 7974 -4643
rect 8008 -4677 8020 -4643
rect 7962 -4711 8020 -4677
rect 7962 -4745 7974 -4711
rect 8008 -4745 8020 -4711
rect 7962 -4760 8020 -4745
rect 8220 -4575 8278 -4560
rect 8220 -4609 8232 -4575
rect 8266 -4609 8278 -4575
rect 8220 -4643 8278 -4609
rect 8220 -4677 8232 -4643
rect 8266 -4677 8278 -4643
rect 8220 -4711 8278 -4677
rect 8220 -4745 8232 -4711
rect 8266 -4745 8278 -4711
rect 8220 -4760 8278 -4745
rect 8478 -4575 8536 -4560
rect 8478 -4609 8490 -4575
rect 8524 -4609 8536 -4575
rect 8478 -4643 8536 -4609
rect 8478 -4677 8490 -4643
rect 8524 -4677 8536 -4643
rect 8478 -4711 8536 -4677
rect 8478 -4745 8490 -4711
rect 8524 -4745 8536 -4711
rect 8478 -4760 8536 -4745
rect 8736 -4575 8794 -4560
rect 8736 -4609 8748 -4575
rect 8782 -4609 8794 -4575
rect 8736 -4643 8794 -4609
rect 8736 -4677 8748 -4643
rect 8782 -4677 8794 -4643
rect 8736 -4711 8794 -4677
rect 8736 -4745 8748 -4711
rect 8782 -4745 8794 -4711
rect 8736 -4760 8794 -4745
rect 8994 -4575 9052 -4560
rect 8994 -4609 9006 -4575
rect 9040 -4609 9052 -4575
rect 8994 -4643 9052 -4609
rect 8994 -4677 9006 -4643
rect 9040 -4677 9052 -4643
rect 8994 -4711 9052 -4677
rect 8994 -4745 9006 -4711
rect 9040 -4745 9052 -4711
rect 8994 -4760 9052 -4745
rect 9188 -4575 9246 -4560
rect 9188 -4609 9200 -4575
rect 9234 -4609 9246 -4575
rect 9188 -4643 9246 -4609
rect 9188 -4677 9200 -4643
rect 9234 -4677 9246 -4643
rect 9188 -4711 9246 -4677
rect 9188 -4745 9200 -4711
rect 9234 -4745 9246 -4711
rect 9188 -4760 9246 -4745
rect 9446 -4575 9504 -4560
rect 9446 -4609 9458 -4575
rect 9492 -4609 9504 -4575
rect 9446 -4643 9504 -4609
rect 9446 -4677 9458 -4643
rect 9492 -4677 9504 -4643
rect 9446 -4711 9504 -4677
rect 9446 -4745 9458 -4711
rect 9492 -4745 9504 -4711
rect 9446 -4760 9504 -4745
rect 9676 -4575 9734 -4560
rect 9676 -4609 9688 -4575
rect 9722 -4609 9734 -4575
rect 9676 -4643 9734 -4609
rect 9676 -4677 9688 -4643
rect 9722 -4677 9734 -4643
rect 9676 -4711 9734 -4677
rect 9676 -4745 9688 -4711
rect 9722 -4745 9734 -4711
rect 9676 -4760 9734 -4745
rect 9934 -4575 9992 -4560
rect 9934 -4609 9946 -4575
rect 9980 -4609 9992 -4575
rect 9934 -4643 9992 -4609
rect 9934 -4677 9946 -4643
rect 9980 -4677 9992 -4643
rect 9934 -4711 9992 -4677
rect 9934 -4745 9946 -4711
rect 9980 -4745 9992 -4711
rect 9934 -4760 9992 -4745
rect 10128 -4575 10186 -4560
rect 10128 -4609 10140 -4575
rect 10174 -4609 10186 -4575
rect 10128 -4643 10186 -4609
rect 10128 -4677 10140 -4643
rect 10174 -4677 10186 -4643
rect 10128 -4711 10186 -4677
rect 10128 -4745 10140 -4711
rect 10174 -4745 10186 -4711
rect 10128 -4760 10186 -4745
rect 10386 -4575 10444 -4560
rect 10386 -4609 10398 -4575
rect 10432 -4609 10444 -4575
rect 10386 -4643 10444 -4609
rect 10386 -4677 10398 -4643
rect 10432 -4677 10444 -4643
rect 10386 -4711 10444 -4677
rect 10386 -4745 10398 -4711
rect 10432 -4745 10444 -4711
rect 10386 -4760 10444 -4745
rect 10644 -4575 10702 -4560
rect 10644 -4609 10656 -4575
rect 10690 -4609 10702 -4575
rect 10644 -4643 10702 -4609
rect 10644 -4677 10656 -4643
rect 10690 -4677 10702 -4643
rect 10644 -4711 10702 -4677
rect 10644 -4745 10656 -4711
rect 10690 -4745 10702 -4711
rect 10644 -4760 10702 -4745
rect 10902 -4575 10960 -4560
rect 10902 -4609 10914 -4575
rect 10948 -4609 10960 -4575
rect 10902 -4643 10960 -4609
rect 10902 -4677 10914 -4643
rect 10948 -4677 10960 -4643
rect 10902 -4711 10960 -4677
rect 10902 -4745 10914 -4711
rect 10948 -4745 10960 -4711
rect 10902 -4760 10960 -4745
rect 11160 -4575 11218 -4560
rect 11160 -4609 11172 -4575
rect 11206 -4609 11218 -4575
rect 11160 -4643 11218 -4609
rect 11160 -4677 11172 -4643
rect 11206 -4677 11218 -4643
rect 11160 -4711 11218 -4677
rect 11160 -4745 11172 -4711
rect 11206 -4745 11218 -4711
rect 11160 -4760 11218 -4745
rect 11354 -4575 11412 -4560
rect 11354 -4609 11366 -4575
rect 11400 -4609 11412 -4575
rect 11354 -4643 11412 -4609
rect 11354 -4677 11366 -4643
rect 11400 -4677 11412 -4643
rect 11354 -4711 11412 -4677
rect 11354 -4745 11366 -4711
rect 11400 -4745 11412 -4711
rect 11354 -4760 11412 -4745
rect 11612 -4575 11670 -4560
rect 11612 -4609 11624 -4575
rect 11658 -4609 11670 -4575
rect 11612 -4643 11670 -4609
rect 11612 -4677 11624 -4643
rect 11658 -4677 11670 -4643
rect 11612 -4711 11670 -4677
rect 11612 -4745 11624 -4711
rect 11658 -4745 11670 -4711
rect 11612 -4760 11670 -4745
rect 11870 -4575 11928 -4560
rect 11870 -4609 11882 -4575
rect 11916 -4609 11928 -4575
rect 11870 -4643 11928 -4609
rect 11870 -4677 11882 -4643
rect 11916 -4677 11928 -4643
rect 11870 -4711 11928 -4677
rect 11870 -4745 11882 -4711
rect 11916 -4745 11928 -4711
rect 11870 -4760 11928 -4745
rect 12128 -4575 12186 -4560
rect 12128 -4609 12140 -4575
rect 12174 -4609 12186 -4575
rect 12128 -4643 12186 -4609
rect 12128 -4677 12140 -4643
rect 12174 -4677 12186 -4643
rect 12128 -4711 12186 -4677
rect 12128 -4745 12140 -4711
rect 12174 -4745 12186 -4711
rect 12128 -4760 12186 -4745
rect 12322 -4575 12380 -4560
rect 12322 -4609 12334 -4575
rect 12368 -4609 12380 -4575
rect 12322 -4643 12380 -4609
rect 12322 -4677 12334 -4643
rect 12368 -4677 12380 -4643
rect 12322 -4711 12380 -4677
rect 12322 -4745 12334 -4711
rect 12368 -4745 12380 -4711
rect 12322 -4760 12380 -4745
rect 12580 -4575 12638 -4560
rect 12580 -4609 12592 -4575
rect 12626 -4609 12638 -4575
rect 12580 -4643 12638 -4609
rect 12580 -4677 12592 -4643
rect 12626 -4677 12638 -4643
rect 12580 -4711 12638 -4677
rect 12580 -4745 12592 -4711
rect 12626 -4745 12638 -4711
rect 12580 -4760 12638 -4745
rect 12838 -4575 12896 -4560
rect 12838 -4609 12850 -4575
rect 12884 -4609 12896 -4575
rect 12838 -4643 12896 -4609
rect 12838 -4677 12850 -4643
rect 12884 -4677 12896 -4643
rect 12838 -4711 12896 -4677
rect 12838 -4745 12850 -4711
rect 12884 -4745 12896 -4711
rect 12838 -4760 12896 -4745
rect 13096 -4575 13154 -4560
rect 13096 -4609 13108 -4575
rect 13142 -4609 13154 -4575
rect 13096 -4643 13154 -4609
rect 13096 -4677 13108 -4643
rect 13142 -4677 13154 -4643
rect 13096 -4711 13154 -4677
rect 13096 -4745 13108 -4711
rect 13142 -4745 13154 -4711
rect 13096 -4760 13154 -4745
rect 13354 -4575 13412 -4560
rect 13354 -4609 13366 -4575
rect 13400 -4609 13412 -4575
rect 13354 -4643 13412 -4609
rect 13354 -4677 13366 -4643
rect 13400 -4677 13412 -4643
rect 13354 -4711 13412 -4677
rect 13354 -4745 13366 -4711
rect 13400 -4745 13412 -4711
rect 13354 -4760 13412 -4745
rect 13548 -4575 13606 -4560
rect 13548 -4609 13560 -4575
rect 13594 -4609 13606 -4575
rect 13548 -4643 13606 -4609
rect 13548 -4677 13560 -4643
rect 13594 -4677 13606 -4643
rect 13548 -4711 13606 -4677
rect 13548 -4745 13560 -4711
rect 13594 -4745 13606 -4711
rect 13548 -4760 13606 -4745
rect 13806 -4575 13864 -4560
rect 13806 -4609 13818 -4575
rect 13852 -4609 13864 -4575
rect 13806 -4643 13864 -4609
rect 13806 -4677 13818 -4643
rect 13852 -4677 13864 -4643
rect 13806 -4711 13864 -4677
rect 13806 -4745 13818 -4711
rect 13852 -4745 13864 -4711
rect 13806 -4760 13864 -4745
rect 14034 -4575 14092 -4560
rect 14034 -4609 14046 -4575
rect 14080 -4609 14092 -4575
rect 14034 -4643 14092 -4609
rect 14034 -4677 14046 -4643
rect 14080 -4677 14092 -4643
rect 14034 -4711 14092 -4677
rect 14034 -4745 14046 -4711
rect 14080 -4745 14092 -4711
rect 14034 -4760 14092 -4745
rect 14292 -4575 14350 -4560
rect 14292 -4609 14304 -4575
rect 14338 -4609 14350 -4575
rect 14292 -4643 14350 -4609
rect 14292 -4677 14304 -4643
rect 14338 -4677 14350 -4643
rect 14292 -4711 14350 -4677
rect 14292 -4745 14304 -4711
rect 14338 -4745 14350 -4711
rect 14292 -4760 14350 -4745
rect 14485 -4575 14543 -4560
rect 14485 -4609 14497 -4575
rect 14531 -4609 14543 -4575
rect 14485 -4643 14543 -4609
rect 14485 -4677 14497 -4643
rect 14531 -4677 14543 -4643
rect 14485 -4711 14543 -4677
rect 14485 -4745 14497 -4711
rect 14531 -4745 14543 -4711
rect 14485 -4760 14543 -4745
rect 14743 -4575 14801 -4560
rect 14743 -4609 14755 -4575
rect 14789 -4609 14801 -4575
rect 14743 -4643 14801 -4609
rect 14743 -4677 14755 -4643
rect 14789 -4677 14801 -4643
rect 14743 -4711 14801 -4677
rect 14743 -4745 14755 -4711
rect 14789 -4745 14801 -4711
rect 14743 -4760 14801 -4745
rect 15001 -4575 15059 -4560
rect 15001 -4609 15013 -4575
rect 15047 -4609 15059 -4575
rect 15001 -4643 15059 -4609
rect 15001 -4677 15013 -4643
rect 15047 -4677 15059 -4643
rect 15001 -4711 15059 -4677
rect 15001 -4745 15013 -4711
rect 15047 -4745 15059 -4711
rect 15001 -4760 15059 -4745
rect 15259 -4575 15317 -4560
rect 15259 -4609 15271 -4575
rect 15305 -4609 15317 -4575
rect 15259 -4643 15317 -4609
rect 15259 -4677 15271 -4643
rect 15305 -4677 15317 -4643
rect 15259 -4711 15317 -4677
rect 15259 -4745 15271 -4711
rect 15305 -4745 15317 -4711
rect 15259 -4760 15317 -4745
rect 15517 -4575 15575 -4560
rect 15517 -4609 15529 -4575
rect 15563 -4609 15575 -4575
rect 15517 -4643 15575 -4609
rect 15517 -4677 15529 -4643
rect 15563 -4677 15575 -4643
rect 15517 -4711 15575 -4677
rect 15517 -4745 15529 -4711
rect 15563 -4745 15575 -4711
rect 15517 -4760 15575 -4745
rect 15711 -4575 15769 -4560
rect 15711 -4609 15723 -4575
rect 15757 -4609 15769 -4575
rect 15711 -4643 15769 -4609
rect 15711 -4677 15723 -4643
rect 15757 -4677 15769 -4643
rect 15711 -4711 15769 -4677
rect 15711 -4745 15723 -4711
rect 15757 -4745 15769 -4711
rect 15711 -4760 15769 -4745
rect 15969 -4575 16027 -4560
rect 15969 -4609 15981 -4575
rect 16015 -4609 16027 -4575
rect 15969 -4643 16027 -4609
rect 15969 -4677 15981 -4643
rect 16015 -4677 16027 -4643
rect 15969 -4711 16027 -4677
rect 15969 -4745 15981 -4711
rect 16015 -4745 16027 -4711
rect 15969 -4760 16027 -4745
rect 16227 -4575 16285 -4560
rect 16227 -4609 16239 -4575
rect 16273 -4609 16285 -4575
rect 16227 -4643 16285 -4609
rect 16227 -4677 16239 -4643
rect 16273 -4677 16285 -4643
rect 16227 -4711 16285 -4677
rect 16227 -4745 16239 -4711
rect 16273 -4745 16285 -4711
rect 16227 -4760 16285 -4745
rect 16485 -4575 16543 -4560
rect 16485 -4609 16497 -4575
rect 16531 -4609 16543 -4575
rect 16485 -4643 16543 -4609
rect 16485 -4677 16497 -4643
rect 16531 -4677 16543 -4643
rect 16485 -4711 16543 -4677
rect 16485 -4745 16497 -4711
rect 16531 -4745 16543 -4711
rect 16485 -4760 16543 -4745
rect 16679 -4575 16737 -4560
rect 16679 -4609 16691 -4575
rect 16725 -4609 16737 -4575
rect 16679 -4643 16737 -4609
rect 16679 -4677 16691 -4643
rect 16725 -4677 16737 -4643
rect 16679 -4711 16737 -4677
rect 16679 -4745 16691 -4711
rect 16725 -4745 16737 -4711
rect 16679 -4760 16737 -4745
rect 16937 -4575 16995 -4560
rect 16937 -4609 16949 -4575
rect 16983 -4609 16995 -4575
rect 16937 -4643 16995 -4609
rect 16937 -4677 16949 -4643
rect 16983 -4677 16995 -4643
rect 16937 -4711 16995 -4677
rect 16937 -4745 16949 -4711
rect 16983 -4745 16995 -4711
rect 16937 -4760 16995 -4745
rect 17195 -4575 17253 -4560
rect 17195 -4609 17207 -4575
rect 17241 -4609 17253 -4575
rect 17195 -4643 17253 -4609
rect 17195 -4677 17207 -4643
rect 17241 -4677 17253 -4643
rect 17195 -4711 17253 -4677
rect 17195 -4745 17207 -4711
rect 17241 -4745 17253 -4711
rect 17195 -4760 17253 -4745
rect 17453 -4575 17511 -4560
rect 17453 -4609 17465 -4575
rect 17499 -4609 17511 -4575
rect 17453 -4643 17511 -4609
rect 17453 -4677 17465 -4643
rect 17499 -4677 17511 -4643
rect 17453 -4711 17511 -4677
rect 17453 -4745 17465 -4711
rect 17499 -4745 17511 -4711
rect 17453 -4760 17511 -4745
rect 17711 -4575 17769 -4560
rect 17711 -4609 17723 -4575
rect 17757 -4609 17769 -4575
rect 17711 -4643 17769 -4609
rect 17711 -4677 17723 -4643
rect 17757 -4677 17769 -4643
rect 17711 -4711 17769 -4677
rect 17711 -4745 17723 -4711
rect 17757 -4745 17769 -4711
rect 17711 -4760 17769 -4745
rect 17905 -4575 17963 -4560
rect 17905 -4609 17917 -4575
rect 17951 -4609 17963 -4575
rect 17905 -4643 17963 -4609
rect 17905 -4677 17917 -4643
rect 17951 -4677 17963 -4643
rect 17905 -4711 17963 -4677
rect 17905 -4745 17917 -4711
rect 17951 -4745 17963 -4711
rect 17905 -4760 17963 -4745
rect 18163 -4575 18221 -4560
rect 18163 -4609 18175 -4575
rect 18209 -4609 18221 -4575
rect 18163 -4643 18221 -4609
rect 18163 -4677 18175 -4643
rect 18209 -4677 18221 -4643
rect 18163 -4711 18221 -4677
rect 18163 -4745 18175 -4711
rect 18209 -4745 18221 -4711
rect 18163 -4760 18221 -4745
rect 959 -5565 1017 -5550
rect 959 -5599 971 -5565
rect 1005 -5599 1017 -5565
rect 959 -5633 1017 -5599
rect 959 -5667 971 -5633
rect 1005 -5667 1017 -5633
rect 959 -5701 1017 -5667
rect 959 -5735 971 -5701
rect 1005 -5735 1017 -5701
rect 959 -5750 1017 -5735
rect 1217 -5565 1275 -5550
rect 1217 -5599 1229 -5565
rect 1263 -5599 1275 -5565
rect 1217 -5633 1275 -5599
rect 1217 -5667 1229 -5633
rect 1263 -5667 1275 -5633
rect 1217 -5701 1275 -5667
rect 1217 -5735 1229 -5701
rect 1263 -5735 1275 -5701
rect 1217 -5750 1275 -5735
rect 1411 -5565 1469 -5550
rect 1411 -5599 1423 -5565
rect 1457 -5599 1469 -5565
rect 1411 -5633 1469 -5599
rect 1411 -5667 1423 -5633
rect 1457 -5667 1469 -5633
rect 1411 -5701 1469 -5667
rect 1411 -5735 1423 -5701
rect 1457 -5735 1469 -5701
rect 1411 -5750 1469 -5735
rect 1669 -5565 1727 -5550
rect 1669 -5599 1681 -5565
rect 1715 -5599 1727 -5565
rect 1669 -5633 1727 -5599
rect 1669 -5667 1681 -5633
rect 1715 -5667 1727 -5633
rect 1669 -5701 1727 -5667
rect 1669 -5735 1681 -5701
rect 1715 -5735 1727 -5701
rect 1669 -5750 1727 -5735
rect 1927 -5565 1985 -5550
rect 1927 -5599 1939 -5565
rect 1973 -5599 1985 -5565
rect 1927 -5633 1985 -5599
rect 1927 -5667 1939 -5633
rect 1973 -5667 1985 -5633
rect 1927 -5701 1985 -5667
rect 1927 -5735 1939 -5701
rect 1973 -5735 1985 -5701
rect 1927 -5750 1985 -5735
rect 2185 -5565 2243 -5550
rect 2185 -5599 2197 -5565
rect 2231 -5599 2243 -5565
rect 2185 -5633 2243 -5599
rect 2185 -5667 2197 -5633
rect 2231 -5667 2243 -5633
rect 2185 -5701 2243 -5667
rect 2185 -5735 2197 -5701
rect 2231 -5735 2243 -5701
rect 2185 -5750 2243 -5735
rect 2443 -5565 2501 -5550
rect 2443 -5599 2455 -5565
rect 2489 -5599 2501 -5565
rect 2443 -5633 2501 -5599
rect 2443 -5667 2455 -5633
rect 2489 -5667 2501 -5633
rect 2443 -5701 2501 -5667
rect 2443 -5735 2455 -5701
rect 2489 -5735 2501 -5701
rect 2443 -5750 2501 -5735
rect 2637 -5565 2695 -5550
rect 2637 -5599 2649 -5565
rect 2683 -5599 2695 -5565
rect 2637 -5633 2695 -5599
rect 2637 -5667 2649 -5633
rect 2683 -5667 2695 -5633
rect 2637 -5701 2695 -5667
rect 2637 -5735 2649 -5701
rect 2683 -5735 2695 -5701
rect 2637 -5750 2695 -5735
rect 2895 -5565 2953 -5550
rect 2895 -5599 2907 -5565
rect 2941 -5599 2953 -5565
rect 2895 -5633 2953 -5599
rect 2895 -5667 2907 -5633
rect 2941 -5667 2953 -5633
rect 2895 -5701 2953 -5667
rect 2895 -5735 2907 -5701
rect 2941 -5735 2953 -5701
rect 2895 -5750 2953 -5735
rect 3153 -5565 3211 -5550
rect 3153 -5599 3165 -5565
rect 3199 -5599 3211 -5565
rect 3153 -5633 3211 -5599
rect 3153 -5667 3165 -5633
rect 3199 -5667 3211 -5633
rect 3153 -5701 3211 -5667
rect 3153 -5735 3165 -5701
rect 3199 -5735 3211 -5701
rect 3153 -5750 3211 -5735
rect 3411 -5565 3469 -5550
rect 3411 -5599 3423 -5565
rect 3457 -5599 3469 -5565
rect 3411 -5633 3469 -5599
rect 3411 -5667 3423 -5633
rect 3457 -5667 3469 -5633
rect 3411 -5701 3469 -5667
rect 3411 -5735 3423 -5701
rect 3457 -5735 3469 -5701
rect 3411 -5750 3469 -5735
rect 3605 -5565 3663 -5550
rect 3605 -5599 3617 -5565
rect 3651 -5599 3663 -5565
rect 3605 -5633 3663 -5599
rect 3605 -5667 3617 -5633
rect 3651 -5667 3663 -5633
rect 3605 -5701 3663 -5667
rect 3605 -5735 3617 -5701
rect 3651 -5735 3663 -5701
rect 3605 -5750 3663 -5735
rect 3863 -5565 3921 -5550
rect 3863 -5599 3875 -5565
rect 3909 -5599 3921 -5565
rect 3863 -5633 3921 -5599
rect 3863 -5667 3875 -5633
rect 3909 -5667 3921 -5633
rect 3863 -5701 3921 -5667
rect 3863 -5735 3875 -5701
rect 3909 -5735 3921 -5701
rect 3863 -5750 3921 -5735
rect 4121 -5565 4179 -5550
rect 4121 -5599 4133 -5565
rect 4167 -5599 4179 -5565
rect 4121 -5633 4179 -5599
rect 4121 -5667 4133 -5633
rect 4167 -5667 4179 -5633
rect 4121 -5701 4179 -5667
rect 4121 -5735 4133 -5701
rect 4167 -5735 4179 -5701
rect 4121 -5750 4179 -5735
rect 4379 -5565 4437 -5550
rect 4379 -5599 4391 -5565
rect 4425 -5599 4437 -5565
rect 4379 -5633 4437 -5599
rect 4379 -5667 4391 -5633
rect 4425 -5667 4437 -5633
rect 4379 -5701 4437 -5667
rect 4379 -5735 4391 -5701
rect 4425 -5735 4437 -5701
rect 4379 -5750 4437 -5735
rect 4637 -5565 4695 -5550
rect 4637 -5599 4649 -5565
rect 4683 -5599 4695 -5565
rect 4637 -5633 4695 -5599
rect 4637 -5667 4649 -5633
rect 4683 -5667 4695 -5633
rect 4637 -5701 4695 -5667
rect 4637 -5735 4649 -5701
rect 4683 -5735 4695 -5701
rect 4637 -5750 4695 -5735
rect 4830 -5565 4888 -5550
rect 4830 -5599 4842 -5565
rect 4876 -5599 4888 -5565
rect 4830 -5633 4888 -5599
rect 4830 -5667 4842 -5633
rect 4876 -5667 4888 -5633
rect 4830 -5701 4888 -5667
rect 4830 -5735 4842 -5701
rect 4876 -5735 4888 -5701
rect 4830 -5750 4888 -5735
rect 5088 -5565 5146 -5550
rect 5088 -5599 5100 -5565
rect 5134 -5599 5146 -5565
rect 5088 -5633 5146 -5599
rect 5088 -5667 5100 -5633
rect 5134 -5667 5146 -5633
rect 5088 -5701 5146 -5667
rect 5088 -5735 5100 -5701
rect 5134 -5735 5146 -5701
rect 5088 -5750 5146 -5735
rect 5316 -5565 5374 -5550
rect 5316 -5599 5328 -5565
rect 5362 -5599 5374 -5565
rect 5316 -5633 5374 -5599
rect 5316 -5667 5328 -5633
rect 5362 -5667 5374 -5633
rect 5316 -5701 5374 -5667
rect 5316 -5735 5328 -5701
rect 5362 -5735 5374 -5701
rect 5316 -5750 5374 -5735
rect 5574 -5565 5632 -5550
rect 5574 -5599 5586 -5565
rect 5620 -5599 5632 -5565
rect 5574 -5633 5632 -5599
rect 5574 -5667 5586 -5633
rect 5620 -5667 5632 -5633
rect 5574 -5701 5632 -5667
rect 5574 -5735 5586 -5701
rect 5620 -5735 5632 -5701
rect 5574 -5750 5632 -5735
rect 5768 -5565 5826 -5550
rect 5768 -5599 5780 -5565
rect 5814 -5599 5826 -5565
rect 5768 -5633 5826 -5599
rect 5768 -5667 5780 -5633
rect 5814 -5667 5826 -5633
rect 5768 -5701 5826 -5667
rect 5768 -5735 5780 -5701
rect 5814 -5735 5826 -5701
rect 5768 -5750 5826 -5735
rect 6026 -5565 6084 -5550
rect 6026 -5599 6038 -5565
rect 6072 -5599 6084 -5565
rect 6026 -5633 6084 -5599
rect 6026 -5667 6038 -5633
rect 6072 -5667 6084 -5633
rect 6026 -5701 6084 -5667
rect 6026 -5735 6038 -5701
rect 6072 -5735 6084 -5701
rect 6026 -5750 6084 -5735
rect 6284 -5565 6342 -5550
rect 6284 -5599 6296 -5565
rect 6330 -5599 6342 -5565
rect 6284 -5633 6342 -5599
rect 6284 -5667 6296 -5633
rect 6330 -5667 6342 -5633
rect 6284 -5701 6342 -5667
rect 6284 -5735 6296 -5701
rect 6330 -5735 6342 -5701
rect 6284 -5750 6342 -5735
rect 6542 -5565 6600 -5550
rect 6542 -5599 6554 -5565
rect 6588 -5599 6600 -5565
rect 6542 -5633 6600 -5599
rect 6542 -5667 6554 -5633
rect 6588 -5667 6600 -5633
rect 6542 -5701 6600 -5667
rect 6542 -5735 6554 -5701
rect 6588 -5735 6600 -5701
rect 6542 -5750 6600 -5735
rect 6800 -5565 6858 -5550
rect 6800 -5599 6812 -5565
rect 6846 -5599 6858 -5565
rect 6800 -5633 6858 -5599
rect 6800 -5667 6812 -5633
rect 6846 -5667 6858 -5633
rect 6800 -5701 6858 -5667
rect 6800 -5735 6812 -5701
rect 6846 -5735 6858 -5701
rect 6800 -5750 6858 -5735
rect 6994 -5565 7052 -5550
rect 6994 -5599 7006 -5565
rect 7040 -5599 7052 -5565
rect 6994 -5633 7052 -5599
rect 6994 -5667 7006 -5633
rect 7040 -5667 7052 -5633
rect 6994 -5701 7052 -5667
rect 6994 -5735 7006 -5701
rect 7040 -5735 7052 -5701
rect 6994 -5750 7052 -5735
rect 7252 -5565 7310 -5550
rect 7252 -5599 7264 -5565
rect 7298 -5599 7310 -5565
rect 7252 -5633 7310 -5599
rect 7252 -5667 7264 -5633
rect 7298 -5667 7310 -5633
rect 7252 -5701 7310 -5667
rect 7252 -5735 7264 -5701
rect 7298 -5735 7310 -5701
rect 7252 -5750 7310 -5735
rect 7510 -5565 7568 -5550
rect 7510 -5599 7522 -5565
rect 7556 -5599 7568 -5565
rect 7510 -5633 7568 -5599
rect 7510 -5667 7522 -5633
rect 7556 -5667 7568 -5633
rect 7510 -5701 7568 -5667
rect 7510 -5735 7522 -5701
rect 7556 -5735 7568 -5701
rect 7510 -5750 7568 -5735
rect 7768 -5565 7826 -5550
rect 7768 -5599 7780 -5565
rect 7814 -5599 7826 -5565
rect 7768 -5633 7826 -5599
rect 7768 -5667 7780 -5633
rect 7814 -5667 7826 -5633
rect 7768 -5701 7826 -5667
rect 7768 -5735 7780 -5701
rect 7814 -5735 7826 -5701
rect 7768 -5750 7826 -5735
rect 7962 -5565 8020 -5550
rect 7962 -5599 7974 -5565
rect 8008 -5599 8020 -5565
rect 7962 -5633 8020 -5599
rect 7962 -5667 7974 -5633
rect 8008 -5667 8020 -5633
rect 7962 -5701 8020 -5667
rect 7962 -5735 7974 -5701
rect 8008 -5735 8020 -5701
rect 7962 -5750 8020 -5735
rect 8220 -5565 8278 -5550
rect 8220 -5599 8232 -5565
rect 8266 -5599 8278 -5565
rect 8220 -5633 8278 -5599
rect 8220 -5667 8232 -5633
rect 8266 -5667 8278 -5633
rect 8220 -5701 8278 -5667
rect 8220 -5735 8232 -5701
rect 8266 -5735 8278 -5701
rect 8220 -5750 8278 -5735
rect 8478 -5565 8536 -5550
rect 8478 -5599 8490 -5565
rect 8524 -5599 8536 -5565
rect 8478 -5633 8536 -5599
rect 8478 -5667 8490 -5633
rect 8524 -5667 8536 -5633
rect 8478 -5701 8536 -5667
rect 8478 -5735 8490 -5701
rect 8524 -5735 8536 -5701
rect 8478 -5750 8536 -5735
rect 8736 -5565 8794 -5550
rect 8736 -5599 8748 -5565
rect 8782 -5599 8794 -5565
rect 8736 -5633 8794 -5599
rect 8736 -5667 8748 -5633
rect 8782 -5667 8794 -5633
rect 8736 -5701 8794 -5667
rect 8736 -5735 8748 -5701
rect 8782 -5735 8794 -5701
rect 8736 -5750 8794 -5735
rect 8994 -5565 9052 -5550
rect 8994 -5599 9006 -5565
rect 9040 -5599 9052 -5565
rect 8994 -5633 9052 -5599
rect 8994 -5667 9006 -5633
rect 9040 -5667 9052 -5633
rect 8994 -5701 9052 -5667
rect 8994 -5735 9006 -5701
rect 9040 -5735 9052 -5701
rect 8994 -5750 9052 -5735
rect 9188 -5565 9246 -5550
rect 9188 -5599 9200 -5565
rect 9234 -5599 9246 -5565
rect 9188 -5633 9246 -5599
rect 9188 -5667 9200 -5633
rect 9234 -5667 9246 -5633
rect 9188 -5701 9246 -5667
rect 9188 -5735 9200 -5701
rect 9234 -5735 9246 -5701
rect 9188 -5750 9246 -5735
rect 9446 -5565 9504 -5550
rect 9446 -5599 9458 -5565
rect 9492 -5599 9504 -5565
rect 9446 -5633 9504 -5599
rect 9446 -5667 9458 -5633
rect 9492 -5667 9504 -5633
rect 9446 -5701 9504 -5667
rect 9446 -5735 9458 -5701
rect 9492 -5735 9504 -5701
rect 9446 -5750 9504 -5735
rect 9676 -5565 9734 -5550
rect 9676 -5599 9688 -5565
rect 9722 -5599 9734 -5565
rect 9676 -5633 9734 -5599
rect 9676 -5667 9688 -5633
rect 9722 -5667 9734 -5633
rect 9676 -5701 9734 -5667
rect 9676 -5735 9688 -5701
rect 9722 -5735 9734 -5701
rect 9676 -5750 9734 -5735
rect 9934 -5565 9992 -5550
rect 9934 -5599 9946 -5565
rect 9980 -5599 9992 -5565
rect 9934 -5633 9992 -5599
rect 9934 -5667 9946 -5633
rect 9980 -5667 9992 -5633
rect 9934 -5701 9992 -5667
rect 9934 -5735 9946 -5701
rect 9980 -5735 9992 -5701
rect 9934 -5750 9992 -5735
rect 10128 -5565 10186 -5550
rect 10128 -5599 10140 -5565
rect 10174 -5599 10186 -5565
rect 10128 -5633 10186 -5599
rect 10128 -5667 10140 -5633
rect 10174 -5667 10186 -5633
rect 10128 -5701 10186 -5667
rect 10128 -5735 10140 -5701
rect 10174 -5735 10186 -5701
rect 10128 -5750 10186 -5735
rect 10386 -5565 10444 -5550
rect 10386 -5599 10398 -5565
rect 10432 -5599 10444 -5565
rect 10386 -5633 10444 -5599
rect 10386 -5667 10398 -5633
rect 10432 -5667 10444 -5633
rect 10386 -5701 10444 -5667
rect 10386 -5735 10398 -5701
rect 10432 -5735 10444 -5701
rect 10386 -5750 10444 -5735
rect 10644 -5565 10702 -5550
rect 10644 -5599 10656 -5565
rect 10690 -5599 10702 -5565
rect 10644 -5633 10702 -5599
rect 10644 -5667 10656 -5633
rect 10690 -5667 10702 -5633
rect 10644 -5701 10702 -5667
rect 10644 -5735 10656 -5701
rect 10690 -5735 10702 -5701
rect 10644 -5750 10702 -5735
rect 10902 -5565 10960 -5550
rect 10902 -5599 10914 -5565
rect 10948 -5599 10960 -5565
rect 10902 -5633 10960 -5599
rect 10902 -5667 10914 -5633
rect 10948 -5667 10960 -5633
rect 10902 -5701 10960 -5667
rect 10902 -5735 10914 -5701
rect 10948 -5735 10960 -5701
rect 10902 -5750 10960 -5735
rect 11160 -5565 11218 -5550
rect 11160 -5599 11172 -5565
rect 11206 -5599 11218 -5565
rect 11160 -5633 11218 -5599
rect 11160 -5667 11172 -5633
rect 11206 -5667 11218 -5633
rect 11160 -5701 11218 -5667
rect 11160 -5735 11172 -5701
rect 11206 -5735 11218 -5701
rect 11160 -5750 11218 -5735
rect 11354 -5565 11412 -5550
rect 11354 -5599 11366 -5565
rect 11400 -5599 11412 -5565
rect 11354 -5633 11412 -5599
rect 11354 -5667 11366 -5633
rect 11400 -5667 11412 -5633
rect 11354 -5701 11412 -5667
rect 11354 -5735 11366 -5701
rect 11400 -5735 11412 -5701
rect 11354 -5750 11412 -5735
rect 11612 -5565 11670 -5550
rect 11612 -5599 11624 -5565
rect 11658 -5599 11670 -5565
rect 11612 -5633 11670 -5599
rect 11612 -5667 11624 -5633
rect 11658 -5667 11670 -5633
rect 11612 -5701 11670 -5667
rect 11612 -5735 11624 -5701
rect 11658 -5735 11670 -5701
rect 11612 -5750 11670 -5735
rect 11870 -5565 11928 -5550
rect 11870 -5599 11882 -5565
rect 11916 -5599 11928 -5565
rect 11870 -5633 11928 -5599
rect 11870 -5667 11882 -5633
rect 11916 -5667 11928 -5633
rect 11870 -5701 11928 -5667
rect 11870 -5735 11882 -5701
rect 11916 -5735 11928 -5701
rect 11870 -5750 11928 -5735
rect 12128 -5565 12186 -5550
rect 12128 -5599 12140 -5565
rect 12174 -5599 12186 -5565
rect 12128 -5633 12186 -5599
rect 12128 -5667 12140 -5633
rect 12174 -5667 12186 -5633
rect 12128 -5701 12186 -5667
rect 12128 -5735 12140 -5701
rect 12174 -5735 12186 -5701
rect 12128 -5750 12186 -5735
rect 12322 -5565 12380 -5550
rect 12322 -5599 12334 -5565
rect 12368 -5599 12380 -5565
rect 12322 -5633 12380 -5599
rect 12322 -5667 12334 -5633
rect 12368 -5667 12380 -5633
rect 12322 -5701 12380 -5667
rect 12322 -5735 12334 -5701
rect 12368 -5735 12380 -5701
rect 12322 -5750 12380 -5735
rect 12580 -5565 12638 -5550
rect 12580 -5599 12592 -5565
rect 12626 -5599 12638 -5565
rect 12580 -5633 12638 -5599
rect 12580 -5667 12592 -5633
rect 12626 -5667 12638 -5633
rect 12580 -5701 12638 -5667
rect 12580 -5735 12592 -5701
rect 12626 -5735 12638 -5701
rect 12580 -5750 12638 -5735
rect 12838 -5565 12896 -5550
rect 12838 -5599 12850 -5565
rect 12884 -5599 12896 -5565
rect 12838 -5633 12896 -5599
rect 12838 -5667 12850 -5633
rect 12884 -5667 12896 -5633
rect 12838 -5701 12896 -5667
rect 12838 -5735 12850 -5701
rect 12884 -5735 12896 -5701
rect 12838 -5750 12896 -5735
rect 13096 -5565 13154 -5550
rect 13096 -5599 13108 -5565
rect 13142 -5599 13154 -5565
rect 13096 -5633 13154 -5599
rect 13096 -5667 13108 -5633
rect 13142 -5667 13154 -5633
rect 13096 -5701 13154 -5667
rect 13096 -5735 13108 -5701
rect 13142 -5735 13154 -5701
rect 13096 -5750 13154 -5735
rect 13354 -5565 13412 -5550
rect 13354 -5599 13366 -5565
rect 13400 -5599 13412 -5565
rect 13354 -5633 13412 -5599
rect 13354 -5667 13366 -5633
rect 13400 -5667 13412 -5633
rect 13354 -5701 13412 -5667
rect 13354 -5735 13366 -5701
rect 13400 -5735 13412 -5701
rect 13354 -5750 13412 -5735
rect 13548 -5565 13606 -5550
rect 13548 -5599 13560 -5565
rect 13594 -5599 13606 -5565
rect 13548 -5633 13606 -5599
rect 13548 -5667 13560 -5633
rect 13594 -5667 13606 -5633
rect 13548 -5701 13606 -5667
rect 13548 -5735 13560 -5701
rect 13594 -5735 13606 -5701
rect 13548 -5750 13606 -5735
rect 13806 -5565 13864 -5550
rect 13806 -5599 13818 -5565
rect 13852 -5599 13864 -5565
rect 13806 -5633 13864 -5599
rect 13806 -5667 13818 -5633
rect 13852 -5667 13864 -5633
rect 13806 -5701 13864 -5667
rect 13806 -5735 13818 -5701
rect 13852 -5735 13864 -5701
rect 13806 -5750 13864 -5735
rect 14034 -5565 14092 -5550
rect 14034 -5599 14046 -5565
rect 14080 -5599 14092 -5565
rect 14034 -5633 14092 -5599
rect 14034 -5667 14046 -5633
rect 14080 -5667 14092 -5633
rect 14034 -5701 14092 -5667
rect 14034 -5735 14046 -5701
rect 14080 -5735 14092 -5701
rect 14034 -5750 14092 -5735
rect 14292 -5565 14350 -5550
rect 14292 -5599 14304 -5565
rect 14338 -5599 14350 -5565
rect 14292 -5633 14350 -5599
rect 14292 -5667 14304 -5633
rect 14338 -5667 14350 -5633
rect 14292 -5701 14350 -5667
rect 14292 -5735 14304 -5701
rect 14338 -5735 14350 -5701
rect 14292 -5750 14350 -5735
rect 14485 -5565 14543 -5550
rect 14485 -5599 14497 -5565
rect 14531 -5599 14543 -5565
rect 14485 -5633 14543 -5599
rect 14485 -5667 14497 -5633
rect 14531 -5667 14543 -5633
rect 14485 -5701 14543 -5667
rect 14485 -5735 14497 -5701
rect 14531 -5735 14543 -5701
rect 14485 -5750 14543 -5735
rect 14743 -5565 14801 -5550
rect 14743 -5599 14755 -5565
rect 14789 -5599 14801 -5565
rect 14743 -5633 14801 -5599
rect 14743 -5667 14755 -5633
rect 14789 -5667 14801 -5633
rect 14743 -5701 14801 -5667
rect 14743 -5735 14755 -5701
rect 14789 -5735 14801 -5701
rect 14743 -5750 14801 -5735
rect 15001 -5565 15059 -5550
rect 15001 -5599 15013 -5565
rect 15047 -5599 15059 -5565
rect 15001 -5633 15059 -5599
rect 15001 -5667 15013 -5633
rect 15047 -5667 15059 -5633
rect 15001 -5701 15059 -5667
rect 15001 -5735 15013 -5701
rect 15047 -5735 15059 -5701
rect 15001 -5750 15059 -5735
rect 15259 -5565 15317 -5550
rect 15259 -5599 15271 -5565
rect 15305 -5599 15317 -5565
rect 15259 -5633 15317 -5599
rect 15259 -5667 15271 -5633
rect 15305 -5667 15317 -5633
rect 15259 -5701 15317 -5667
rect 15259 -5735 15271 -5701
rect 15305 -5735 15317 -5701
rect 15259 -5750 15317 -5735
rect 15517 -5565 15575 -5550
rect 15517 -5599 15529 -5565
rect 15563 -5599 15575 -5565
rect 15517 -5633 15575 -5599
rect 15517 -5667 15529 -5633
rect 15563 -5667 15575 -5633
rect 15517 -5701 15575 -5667
rect 15517 -5735 15529 -5701
rect 15563 -5735 15575 -5701
rect 15517 -5750 15575 -5735
rect 15711 -5565 15769 -5550
rect 15711 -5599 15723 -5565
rect 15757 -5599 15769 -5565
rect 15711 -5633 15769 -5599
rect 15711 -5667 15723 -5633
rect 15757 -5667 15769 -5633
rect 15711 -5701 15769 -5667
rect 15711 -5735 15723 -5701
rect 15757 -5735 15769 -5701
rect 15711 -5750 15769 -5735
rect 15969 -5565 16027 -5550
rect 15969 -5599 15981 -5565
rect 16015 -5599 16027 -5565
rect 15969 -5633 16027 -5599
rect 15969 -5667 15981 -5633
rect 16015 -5667 16027 -5633
rect 15969 -5701 16027 -5667
rect 15969 -5735 15981 -5701
rect 16015 -5735 16027 -5701
rect 15969 -5750 16027 -5735
rect 16227 -5565 16285 -5550
rect 16227 -5599 16239 -5565
rect 16273 -5599 16285 -5565
rect 16227 -5633 16285 -5599
rect 16227 -5667 16239 -5633
rect 16273 -5667 16285 -5633
rect 16227 -5701 16285 -5667
rect 16227 -5735 16239 -5701
rect 16273 -5735 16285 -5701
rect 16227 -5750 16285 -5735
rect 16485 -5565 16543 -5550
rect 16485 -5599 16497 -5565
rect 16531 -5599 16543 -5565
rect 16485 -5633 16543 -5599
rect 16485 -5667 16497 -5633
rect 16531 -5667 16543 -5633
rect 16485 -5701 16543 -5667
rect 16485 -5735 16497 -5701
rect 16531 -5735 16543 -5701
rect 16485 -5750 16543 -5735
rect 16679 -5565 16737 -5550
rect 16679 -5599 16691 -5565
rect 16725 -5599 16737 -5565
rect 16679 -5633 16737 -5599
rect 16679 -5667 16691 -5633
rect 16725 -5667 16737 -5633
rect 16679 -5701 16737 -5667
rect 16679 -5735 16691 -5701
rect 16725 -5735 16737 -5701
rect 16679 -5750 16737 -5735
rect 16937 -5565 16995 -5550
rect 16937 -5599 16949 -5565
rect 16983 -5599 16995 -5565
rect 16937 -5633 16995 -5599
rect 16937 -5667 16949 -5633
rect 16983 -5667 16995 -5633
rect 16937 -5701 16995 -5667
rect 16937 -5735 16949 -5701
rect 16983 -5735 16995 -5701
rect 16937 -5750 16995 -5735
rect 17195 -5565 17253 -5550
rect 17195 -5599 17207 -5565
rect 17241 -5599 17253 -5565
rect 17195 -5633 17253 -5599
rect 17195 -5667 17207 -5633
rect 17241 -5667 17253 -5633
rect 17195 -5701 17253 -5667
rect 17195 -5735 17207 -5701
rect 17241 -5735 17253 -5701
rect 17195 -5750 17253 -5735
rect 17453 -5565 17511 -5550
rect 17453 -5599 17465 -5565
rect 17499 -5599 17511 -5565
rect 17453 -5633 17511 -5599
rect 17453 -5667 17465 -5633
rect 17499 -5667 17511 -5633
rect 17453 -5701 17511 -5667
rect 17453 -5735 17465 -5701
rect 17499 -5735 17511 -5701
rect 17453 -5750 17511 -5735
rect 17711 -5565 17769 -5550
rect 17711 -5599 17723 -5565
rect 17757 -5599 17769 -5565
rect 17711 -5633 17769 -5599
rect 17711 -5667 17723 -5633
rect 17757 -5667 17769 -5633
rect 17711 -5701 17769 -5667
rect 17711 -5735 17723 -5701
rect 17757 -5735 17769 -5701
rect 17711 -5750 17769 -5735
rect 17905 -5565 17963 -5550
rect 17905 -5599 17917 -5565
rect 17951 -5599 17963 -5565
rect 17905 -5633 17963 -5599
rect 17905 -5667 17917 -5633
rect 17951 -5667 17963 -5633
rect 17905 -5701 17963 -5667
rect 17905 -5735 17917 -5701
rect 17951 -5735 17963 -5701
rect 17905 -5750 17963 -5735
rect 18163 -5565 18221 -5550
rect 18163 -5599 18175 -5565
rect 18209 -5599 18221 -5565
rect 18163 -5633 18221 -5599
rect 18163 -5667 18175 -5633
rect 18209 -5667 18221 -5633
rect 18163 -5701 18221 -5667
rect 18163 -5735 18175 -5701
rect 18209 -5735 18221 -5701
rect 18163 -5750 18221 -5735
rect 959 -6255 1017 -6240
rect 959 -6289 971 -6255
rect 1005 -6289 1017 -6255
rect 959 -6323 1017 -6289
rect 959 -6357 971 -6323
rect 1005 -6357 1017 -6323
rect 959 -6391 1017 -6357
rect 959 -6425 971 -6391
rect 1005 -6425 1017 -6391
rect 959 -6440 1017 -6425
rect 1217 -6255 1275 -6240
rect 1217 -6289 1229 -6255
rect 1263 -6289 1275 -6255
rect 1217 -6323 1275 -6289
rect 1217 -6357 1229 -6323
rect 1263 -6357 1275 -6323
rect 1217 -6391 1275 -6357
rect 1217 -6425 1229 -6391
rect 1263 -6425 1275 -6391
rect 1217 -6440 1275 -6425
rect 1411 -6255 1469 -6240
rect 1411 -6289 1423 -6255
rect 1457 -6289 1469 -6255
rect 1411 -6323 1469 -6289
rect 1411 -6357 1423 -6323
rect 1457 -6357 1469 -6323
rect 1411 -6391 1469 -6357
rect 1411 -6425 1423 -6391
rect 1457 -6425 1469 -6391
rect 1411 -6440 1469 -6425
rect 1669 -6255 1727 -6240
rect 1669 -6289 1681 -6255
rect 1715 -6289 1727 -6255
rect 1669 -6323 1727 -6289
rect 1669 -6357 1681 -6323
rect 1715 -6357 1727 -6323
rect 1669 -6391 1727 -6357
rect 1669 -6425 1681 -6391
rect 1715 -6425 1727 -6391
rect 1669 -6440 1727 -6425
rect 1927 -6255 1985 -6240
rect 1927 -6289 1939 -6255
rect 1973 -6289 1985 -6255
rect 1927 -6323 1985 -6289
rect 1927 -6357 1939 -6323
rect 1973 -6357 1985 -6323
rect 1927 -6391 1985 -6357
rect 1927 -6425 1939 -6391
rect 1973 -6425 1985 -6391
rect 1927 -6440 1985 -6425
rect 2185 -6255 2243 -6240
rect 2185 -6289 2197 -6255
rect 2231 -6289 2243 -6255
rect 2185 -6323 2243 -6289
rect 2185 -6357 2197 -6323
rect 2231 -6357 2243 -6323
rect 2185 -6391 2243 -6357
rect 2185 -6425 2197 -6391
rect 2231 -6425 2243 -6391
rect 2185 -6440 2243 -6425
rect 2443 -6255 2501 -6240
rect 2443 -6289 2455 -6255
rect 2489 -6289 2501 -6255
rect 2443 -6323 2501 -6289
rect 2443 -6357 2455 -6323
rect 2489 -6357 2501 -6323
rect 2443 -6391 2501 -6357
rect 2443 -6425 2455 -6391
rect 2489 -6425 2501 -6391
rect 2443 -6440 2501 -6425
rect 2637 -6255 2695 -6240
rect 2637 -6289 2649 -6255
rect 2683 -6289 2695 -6255
rect 2637 -6323 2695 -6289
rect 2637 -6357 2649 -6323
rect 2683 -6357 2695 -6323
rect 2637 -6391 2695 -6357
rect 2637 -6425 2649 -6391
rect 2683 -6425 2695 -6391
rect 2637 -6440 2695 -6425
rect 2895 -6255 2953 -6240
rect 2895 -6289 2907 -6255
rect 2941 -6289 2953 -6255
rect 2895 -6323 2953 -6289
rect 2895 -6357 2907 -6323
rect 2941 -6357 2953 -6323
rect 2895 -6391 2953 -6357
rect 2895 -6425 2907 -6391
rect 2941 -6425 2953 -6391
rect 2895 -6440 2953 -6425
rect 3153 -6255 3211 -6240
rect 3153 -6289 3165 -6255
rect 3199 -6289 3211 -6255
rect 3153 -6323 3211 -6289
rect 3153 -6357 3165 -6323
rect 3199 -6357 3211 -6323
rect 3153 -6391 3211 -6357
rect 3153 -6425 3165 -6391
rect 3199 -6425 3211 -6391
rect 3153 -6440 3211 -6425
rect 3411 -6255 3469 -6240
rect 3411 -6289 3423 -6255
rect 3457 -6289 3469 -6255
rect 3411 -6323 3469 -6289
rect 3411 -6357 3423 -6323
rect 3457 -6357 3469 -6323
rect 3411 -6391 3469 -6357
rect 3411 -6425 3423 -6391
rect 3457 -6425 3469 -6391
rect 3411 -6440 3469 -6425
rect 3605 -6255 3663 -6240
rect 3605 -6289 3617 -6255
rect 3651 -6289 3663 -6255
rect 3605 -6323 3663 -6289
rect 3605 -6357 3617 -6323
rect 3651 -6357 3663 -6323
rect 3605 -6391 3663 -6357
rect 3605 -6425 3617 -6391
rect 3651 -6425 3663 -6391
rect 3605 -6440 3663 -6425
rect 3863 -6255 3921 -6240
rect 3863 -6289 3875 -6255
rect 3909 -6289 3921 -6255
rect 3863 -6323 3921 -6289
rect 3863 -6357 3875 -6323
rect 3909 -6357 3921 -6323
rect 3863 -6391 3921 -6357
rect 3863 -6425 3875 -6391
rect 3909 -6425 3921 -6391
rect 3863 -6440 3921 -6425
rect 4121 -6255 4179 -6240
rect 4121 -6289 4133 -6255
rect 4167 -6289 4179 -6255
rect 4121 -6323 4179 -6289
rect 4121 -6357 4133 -6323
rect 4167 -6357 4179 -6323
rect 4121 -6391 4179 -6357
rect 4121 -6425 4133 -6391
rect 4167 -6425 4179 -6391
rect 4121 -6440 4179 -6425
rect 4379 -6255 4437 -6240
rect 4379 -6289 4391 -6255
rect 4425 -6289 4437 -6255
rect 4379 -6323 4437 -6289
rect 4379 -6357 4391 -6323
rect 4425 -6357 4437 -6323
rect 4379 -6391 4437 -6357
rect 4379 -6425 4391 -6391
rect 4425 -6425 4437 -6391
rect 4379 -6440 4437 -6425
rect 4637 -6255 4695 -6240
rect 4637 -6289 4649 -6255
rect 4683 -6289 4695 -6255
rect 4637 -6323 4695 -6289
rect 4637 -6357 4649 -6323
rect 4683 -6357 4695 -6323
rect 4637 -6391 4695 -6357
rect 4637 -6425 4649 -6391
rect 4683 -6425 4695 -6391
rect 4637 -6440 4695 -6425
rect 4830 -6255 4888 -6240
rect 4830 -6289 4842 -6255
rect 4876 -6289 4888 -6255
rect 4830 -6323 4888 -6289
rect 4830 -6357 4842 -6323
rect 4876 -6357 4888 -6323
rect 4830 -6391 4888 -6357
rect 4830 -6425 4842 -6391
rect 4876 -6425 4888 -6391
rect 4830 -6440 4888 -6425
rect 5088 -6255 5146 -6240
rect 5088 -6289 5100 -6255
rect 5134 -6289 5146 -6255
rect 5088 -6323 5146 -6289
rect 5088 -6357 5100 -6323
rect 5134 -6357 5146 -6323
rect 5088 -6391 5146 -6357
rect 5088 -6425 5100 -6391
rect 5134 -6425 5146 -6391
rect 5088 -6440 5146 -6425
rect 5316 -6255 5374 -6240
rect 5316 -6289 5328 -6255
rect 5362 -6289 5374 -6255
rect 5316 -6323 5374 -6289
rect 5316 -6357 5328 -6323
rect 5362 -6357 5374 -6323
rect 5316 -6391 5374 -6357
rect 5316 -6425 5328 -6391
rect 5362 -6425 5374 -6391
rect 5316 -6440 5374 -6425
rect 5574 -6255 5632 -6240
rect 5574 -6289 5586 -6255
rect 5620 -6289 5632 -6255
rect 5574 -6323 5632 -6289
rect 5574 -6357 5586 -6323
rect 5620 -6357 5632 -6323
rect 5574 -6391 5632 -6357
rect 5574 -6425 5586 -6391
rect 5620 -6425 5632 -6391
rect 5574 -6440 5632 -6425
rect 5768 -6255 5826 -6240
rect 5768 -6289 5780 -6255
rect 5814 -6289 5826 -6255
rect 5768 -6323 5826 -6289
rect 5768 -6357 5780 -6323
rect 5814 -6357 5826 -6323
rect 5768 -6391 5826 -6357
rect 5768 -6425 5780 -6391
rect 5814 -6425 5826 -6391
rect 5768 -6440 5826 -6425
rect 6026 -6255 6084 -6240
rect 6026 -6289 6038 -6255
rect 6072 -6289 6084 -6255
rect 6026 -6323 6084 -6289
rect 6026 -6357 6038 -6323
rect 6072 -6357 6084 -6323
rect 6026 -6391 6084 -6357
rect 6026 -6425 6038 -6391
rect 6072 -6425 6084 -6391
rect 6026 -6440 6084 -6425
rect 6284 -6255 6342 -6240
rect 6284 -6289 6296 -6255
rect 6330 -6289 6342 -6255
rect 6284 -6323 6342 -6289
rect 6284 -6357 6296 -6323
rect 6330 -6357 6342 -6323
rect 6284 -6391 6342 -6357
rect 6284 -6425 6296 -6391
rect 6330 -6425 6342 -6391
rect 6284 -6440 6342 -6425
rect 6542 -6255 6600 -6240
rect 6542 -6289 6554 -6255
rect 6588 -6289 6600 -6255
rect 6542 -6323 6600 -6289
rect 6542 -6357 6554 -6323
rect 6588 -6357 6600 -6323
rect 6542 -6391 6600 -6357
rect 6542 -6425 6554 -6391
rect 6588 -6425 6600 -6391
rect 6542 -6440 6600 -6425
rect 6800 -6255 6858 -6240
rect 6800 -6289 6812 -6255
rect 6846 -6289 6858 -6255
rect 6800 -6323 6858 -6289
rect 6800 -6357 6812 -6323
rect 6846 -6357 6858 -6323
rect 6800 -6391 6858 -6357
rect 6800 -6425 6812 -6391
rect 6846 -6425 6858 -6391
rect 6800 -6440 6858 -6425
rect 6994 -6255 7052 -6240
rect 6994 -6289 7006 -6255
rect 7040 -6289 7052 -6255
rect 6994 -6323 7052 -6289
rect 6994 -6357 7006 -6323
rect 7040 -6357 7052 -6323
rect 6994 -6391 7052 -6357
rect 6994 -6425 7006 -6391
rect 7040 -6425 7052 -6391
rect 6994 -6440 7052 -6425
rect 7252 -6255 7310 -6240
rect 7252 -6289 7264 -6255
rect 7298 -6289 7310 -6255
rect 7252 -6323 7310 -6289
rect 7252 -6357 7264 -6323
rect 7298 -6357 7310 -6323
rect 7252 -6391 7310 -6357
rect 7252 -6425 7264 -6391
rect 7298 -6425 7310 -6391
rect 7252 -6440 7310 -6425
rect 7510 -6255 7568 -6240
rect 7510 -6289 7522 -6255
rect 7556 -6289 7568 -6255
rect 7510 -6323 7568 -6289
rect 7510 -6357 7522 -6323
rect 7556 -6357 7568 -6323
rect 7510 -6391 7568 -6357
rect 7510 -6425 7522 -6391
rect 7556 -6425 7568 -6391
rect 7510 -6440 7568 -6425
rect 7768 -6255 7826 -6240
rect 7768 -6289 7780 -6255
rect 7814 -6289 7826 -6255
rect 7768 -6323 7826 -6289
rect 7768 -6357 7780 -6323
rect 7814 -6357 7826 -6323
rect 7768 -6391 7826 -6357
rect 7768 -6425 7780 -6391
rect 7814 -6425 7826 -6391
rect 7768 -6440 7826 -6425
rect 7962 -6255 8020 -6240
rect 7962 -6289 7974 -6255
rect 8008 -6289 8020 -6255
rect 7962 -6323 8020 -6289
rect 7962 -6357 7974 -6323
rect 8008 -6357 8020 -6323
rect 7962 -6391 8020 -6357
rect 7962 -6425 7974 -6391
rect 8008 -6425 8020 -6391
rect 7962 -6440 8020 -6425
rect 8220 -6255 8278 -6240
rect 8220 -6289 8232 -6255
rect 8266 -6289 8278 -6255
rect 8220 -6323 8278 -6289
rect 8220 -6357 8232 -6323
rect 8266 -6357 8278 -6323
rect 8220 -6391 8278 -6357
rect 8220 -6425 8232 -6391
rect 8266 -6425 8278 -6391
rect 8220 -6440 8278 -6425
rect 8478 -6255 8536 -6240
rect 8478 -6289 8490 -6255
rect 8524 -6289 8536 -6255
rect 8478 -6323 8536 -6289
rect 8478 -6357 8490 -6323
rect 8524 -6357 8536 -6323
rect 8478 -6391 8536 -6357
rect 8478 -6425 8490 -6391
rect 8524 -6425 8536 -6391
rect 8478 -6440 8536 -6425
rect 8736 -6255 8794 -6240
rect 8736 -6289 8748 -6255
rect 8782 -6289 8794 -6255
rect 8736 -6323 8794 -6289
rect 8736 -6357 8748 -6323
rect 8782 -6357 8794 -6323
rect 8736 -6391 8794 -6357
rect 8736 -6425 8748 -6391
rect 8782 -6425 8794 -6391
rect 8736 -6440 8794 -6425
rect 8994 -6255 9052 -6240
rect 8994 -6289 9006 -6255
rect 9040 -6289 9052 -6255
rect 8994 -6323 9052 -6289
rect 8994 -6357 9006 -6323
rect 9040 -6357 9052 -6323
rect 8994 -6391 9052 -6357
rect 8994 -6425 9006 -6391
rect 9040 -6425 9052 -6391
rect 8994 -6440 9052 -6425
rect 9188 -6255 9246 -6240
rect 9188 -6289 9200 -6255
rect 9234 -6289 9246 -6255
rect 9188 -6323 9246 -6289
rect 9188 -6357 9200 -6323
rect 9234 -6357 9246 -6323
rect 9188 -6391 9246 -6357
rect 9188 -6425 9200 -6391
rect 9234 -6425 9246 -6391
rect 9188 -6440 9246 -6425
rect 9446 -6255 9504 -6240
rect 9446 -6289 9458 -6255
rect 9492 -6289 9504 -6255
rect 9446 -6323 9504 -6289
rect 9446 -6357 9458 -6323
rect 9492 -6357 9504 -6323
rect 9446 -6391 9504 -6357
rect 9446 -6425 9458 -6391
rect 9492 -6425 9504 -6391
rect 9446 -6440 9504 -6425
rect 9676 -6255 9734 -6240
rect 9676 -6289 9688 -6255
rect 9722 -6289 9734 -6255
rect 9676 -6323 9734 -6289
rect 9676 -6357 9688 -6323
rect 9722 -6357 9734 -6323
rect 9676 -6391 9734 -6357
rect 9676 -6425 9688 -6391
rect 9722 -6425 9734 -6391
rect 9676 -6440 9734 -6425
rect 9934 -6255 9992 -6240
rect 9934 -6289 9946 -6255
rect 9980 -6289 9992 -6255
rect 9934 -6323 9992 -6289
rect 9934 -6357 9946 -6323
rect 9980 -6357 9992 -6323
rect 9934 -6391 9992 -6357
rect 9934 -6425 9946 -6391
rect 9980 -6425 9992 -6391
rect 9934 -6440 9992 -6425
rect 10128 -6255 10186 -6240
rect 10128 -6289 10140 -6255
rect 10174 -6289 10186 -6255
rect 10128 -6323 10186 -6289
rect 10128 -6357 10140 -6323
rect 10174 -6357 10186 -6323
rect 10128 -6391 10186 -6357
rect 10128 -6425 10140 -6391
rect 10174 -6425 10186 -6391
rect 10128 -6440 10186 -6425
rect 10386 -6255 10444 -6240
rect 10386 -6289 10398 -6255
rect 10432 -6289 10444 -6255
rect 10386 -6323 10444 -6289
rect 10386 -6357 10398 -6323
rect 10432 -6357 10444 -6323
rect 10386 -6391 10444 -6357
rect 10386 -6425 10398 -6391
rect 10432 -6425 10444 -6391
rect 10386 -6440 10444 -6425
rect 10644 -6255 10702 -6240
rect 10644 -6289 10656 -6255
rect 10690 -6289 10702 -6255
rect 10644 -6323 10702 -6289
rect 10644 -6357 10656 -6323
rect 10690 -6357 10702 -6323
rect 10644 -6391 10702 -6357
rect 10644 -6425 10656 -6391
rect 10690 -6425 10702 -6391
rect 10644 -6440 10702 -6425
rect 10902 -6255 10960 -6240
rect 10902 -6289 10914 -6255
rect 10948 -6289 10960 -6255
rect 10902 -6323 10960 -6289
rect 10902 -6357 10914 -6323
rect 10948 -6357 10960 -6323
rect 10902 -6391 10960 -6357
rect 10902 -6425 10914 -6391
rect 10948 -6425 10960 -6391
rect 10902 -6440 10960 -6425
rect 11160 -6255 11218 -6240
rect 11160 -6289 11172 -6255
rect 11206 -6289 11218 -6255
rect 11160 -6323 11218 -6289
rect 11160 -6357 11172 -6323
rect 11206 -6357 11218 -6323
rect 11160 -6391 11218 -6357
rect 11160 -6425 11172 -6391
rect 11206 -6425 11218 -6391
rect 11160 -6440 11218 -6425
rect 11354 -6255 11412 -6240
rect 11354 -6289 11366 -6255
rect 11400 -6289 11412 -6255
rect 11354 -6323 11412 -6289
rect 11354 -6357 11366 -6323
rect 11400 -6357 11412 -6323
rect 11354 -6391 11412 -6357
rect 11354 -6425 11366 -6391
rect 11400 -6425 11412 -6391
rect 11354 -6440 11412 -6425
rect 11612 -6255 11670 -6240
rect 11612 -6289 11624 -6255
rect 11658 -6289 11670 -6255
rect 11612 -6323 11670 -6289
rect 11612 -6357 11624 -6323
rect 11658 -6357 11670 -6323
rect 11612 -6391 11670 -6357
rect 11612 -6425 11624 -6391
rect 11658 -6425 11670 -6391
rect 11612 -6440 11670 -6425
rect 11870 -6255 11928 -6240
rect 11870 -6289 11882 -6255
rect 11916 -6289 11928 -6255
rect 11870 -6323 11928 -6289
rect 11870 -6357 11882 -6323
rect 11916 -6357 11928 -6323
rect 11870 -6391 11928 -6357
rect 11870 -6425 11882 -6391
rect 11916 -6425 11928 -6391
rect 11870 -6440 11928 -6425
rect 12128 -6255 12186 -6240
rect 12128 -6289 12140 -6255
rect 12174 -6289 12186 -6255
rect 12128 -6323 12186 -6289
rect 12128 -6357 12140 -6323
rect 12174 -6357 12186 -6323
rect 12128 -6391 12186 -6357
rect 12128 -6425 12140 -6391
rect 12174 -6425 12186 -6391
rect 12128 -6440 12186 -6425
rect 12322 -6255 12380 -6240
rect 12322 -6289 12334 -6255
rect 12368 -6289 12380 -6255
rect 12322 -6323 12380 -6289
rect 12322 -6357 12334 -6323
rect 12368 -6357 12380 -6323
rect 12322 -6391 12380 -6357
rect 12322 -6425 12334 -6391
rect 12368 -6425 12380 -6391
rect 12322 -6440 12380 -6425
rect 12580 -6255 12638 -6240
rect 12580 -6289 12592 -6255
rect 12626 -6289 12638 -6255
rect 12580 -6323 12638 -6289
rect 12580 -6357 12592 -6323
rect 12626 -6357 12638 -6323
rect 12580 -6391 12638 -6357
rect 12580 -6425 12592 -6391
rect 12626 -6425 12638 -6391
rect 12580 -6440 12638 -6425
rect 12838 -6255 12896 -6240
rect 12838 -6289 12850 -6255
rect 12884 -6289 12896 -6255
rect 12838 -6323 12896 -6289
rect 12838 -6357 12850 -6323
rect 12884 -6357 12896 -6323
rect 12838 -6391 12896 -6357
rect 12838 -6425 12850 -6391
rect 12884 -6425 12896 -6391
rect 12838 -6440 12896 -6425
rect 13096 -6255 13154 -6240
rect 13096 -6289 13108 -6255
rect 13142 -6289 13154 -6255
rect 13096 -6323 13154 -6289
rect 13096 -6357 13108 -6323
rect 13142 -6357 13154 -6323
rect 13096 -6391 13154 -6357
rect 13096 -6425 13108 -6391
rect 13142 -6425 13154 -6391
rect 13096 -6440 13154 -6425
rect 13354 -6255 13412 -6240
rect 13354 -6289 13366 -6255
rect 13400 -6289 13412 -6255
rect 13354 -6323 13412 -6289
rect 13354 -6357 13366 -6323
rect 13400 -6357 13412 -6323
rect 13354 -6391 13412 -6357
rect 13354 -6425 13366 -6391
rect 13400 -6425 13412 -6391
rect 13354 -6440 13412 -6425
rect 13548 -6255 13606 -6240
rect 13548 -6289 13560 -6255
rect 13594 -6289 13606 -6255
rect 13548 -6323 13606 -6289
rect 13548 -6357 13560 -6323
rect 13594 -6357 13606 -6323
rect 13548 -6391 13606 -6357
rect 13548 -6425 13560 -6391
rect 13594 -6425 13606 -6391
rect 13548 -6440 13606 -6425
rect 13806 -6255 13864 -6240
rect 13806 -6289 13818 -6255
rect 13852 -6289 13864 -6255
rect 13806 -6323 13864 -6289
rect 13806 -6357 13818 -6323
rect 13852 -6357 13864 -6323
rect 13806 -6391 13864 -6357
rect 13806 -6425 13818 -6391
rect 13852 -6425 13864 -6391
rect 13806 -6440 13864 -6425
rect 14034 -6255 14092 -6240
rect 14034 -6289 14046 -6255
rect 14080 -6289 14092 -6255
rect 14034 -6323 14092 -6289
rect 14034 -6357 14046 -6323
rect 14080 -6357 14092 -6323
rect 14034 -6391 14092 -6357
rect 14034 -6425 14046 -6391
rect 14080 -6425 14092 -6391
rect 14034 -6440 14092 -6425
rect 14292 -6255 14350 -6240
rect 14292 -6289 14304 -6255
rect 14338 -6289 14350 -6255
rect 14292 -6323 14350 -6289
rect 14292 -6357 14304 -6323
rect 14338 -6357 14350 -6323
rect 14292 -6391 14350 -6357
rect 14292 -6425 14304 -6391
rect 14338 -6425 14350 -6391
rect 14292 -6440 14350 -6425
rect 14485 -6255 14543 -6240
rect 14485 -6289 14497 -6255
rect 14531 -6289 14543 -6255
rect 14485 -6323 14543 -6289
rect 14485 -6357 14497 -6323
rect 14531 -6357 14543 -6323
rect 14485 -6391 14543 -6357
rect 14485 -6425 14497 -6391
rect 14531 -6425 14543 -6391
rect 14485 -6440 14543 -6425
rect 14743 -6255 14801 -6240
rect 14743 -6289 14755 -6255
rect 14789 -6289 14801 -6255
rect 14743 -6323 14801 -6289
rect 14743 -6357 14755 -6323
rect 14789 -6357 14801 -6323
rect 14743 -6391 14801 -6357
rect 14743 -6425 14755 -6391
rect 14789 -6425 14801 -6391
rect 14743 -6440 14801 -6425
rect 15001 -6255 15059 -6240
rect 15001 -6289 15013 -6255
rect 15047 -6289 15059 -6255
rect 15001 -6323 15059 -6289
rect 15001 -6357 15013 -6323
rect 15047 -6357 15059 -6323
rect 15001 -6391 15059 -6357
rect 15001 -6425 15013 -6391
rect 15047 -6425 15059 -6391
rect 15001 -6440 15059 -6425
rect 15259 -6255 15317 -6240
rect 15259 -6289 15271 -6255
rect 15305 -6289 15317 -6255
rect 15259 -6323 15317 -6289
rect 15259 -6357 15271 -6323
rect 15305 -6357 15317 -6323
rect 15259 -6391 15317 -6357
rect 15259 -6425 15271 -6391
rect 15305 -6425 15317 -6391
rect 15259 -6440 15317 -6425
rect 15517 -6255 15575 -6240
rect 15517 -6289 15529 -6255
rect 15563 -6289 15575 -6255
rect 15517 -6323 15575 -6289
rect 15517 -6357 15529 -6323
rect 15563 -6357 15575 -6323
rect 15517 -6391 15575 -6357
rect 15517 -6425 15529 -6391
rect 15563 -6425 15575 -6391
rect 15517 -6440 15575 -6425
rect 15711 -6255 15769 -6240
rect 15711 -6289 15723 -6255
rect 15757 -6289 15769 -6255
rect 15711 -6323 15769 -6289
rect 15711 -6357 15723 -6323
rect 15757 -6357 15769 -6323
rect 15711 -6391 15769 -6357
rect 15711 -6425 15723 -6391
rect 15757 -6425 15769 -6391
rect 15711 -6440 15769 -6425
rect 15969 -6255 16027 -6240
rect 15969 -6289 15981 -6255
rect 16015 -6289 16027 -6255
rect 15969 -6323 16027 -6289
rect 15969 -6357 15981 -6323
rect 16015 -6357 16027 -6323
rect 15969 -6391 16027 -6357
rect 15969 -6425 15981 -6391
rect 16015 -6425 16027 -6391
rect 15969 -6440 16027 -6425
rect 16227 -6255 16285 -6240
rect 16227 -6289 16239 -6255
rect 16273 -6289 16285 -6255
rect 16227 -6323 16285 -6289
rect 16227 -6357 16239 -6323
rect 16273 -6357 16285 -6323
rect 16227 -6391 16285 -6357
rect 16227 -6425 16239 -6391
rect 16273 -6425 16285 -6391
rect 16227 -6440 16285 -6425
rect 16485 -6255 16543 -6240
rect 16485 -6289 16497 -6255
rect 16531 -6289 16543 -6255
rect 16485 -6323 16543 -6289
rect 16485 -6357 16497 -6323
rect 16531 -6357 16543 -6323
rect 16485 -6391 16543 -6357
rect 16485 -6425 16497 -6391
rect 16531 -6425 16543 -6391
rect 16485 -6440 16543 -6425
rect 16679 -6255 16737 -6240
rect 16679 -6289 16691 -6255
rect 16725 -6289 16737 -6255
rect 16679 -6323 16737 -6289
rect 16679 -6357 16691 -6323
rect 16725 -6357 16737 -6323
rect 16679 -6391 16737 -6357
rect 16679 -6425 16691 -6391
rect 16725 -6425 16737 -6391
rect 16679 -6440 16737 -6425
rect 16937 -6255 16995 -6240
rect 16937 -6289 16949 -6255
rect 16983 -6289 16995 -6255
rect 16937 -6323 16995 -6289
rect 16937 -6357 16949 -6323
rect 16983 -6357 16995 -6323
rect 16937 -6391 16995 -6357
rect 16937 -6425 16949 -6391
rect 16983 -6425 16995 -6391
rect 16937 -6440 16995 -6425
rect 17195 -6255 17253 -6240
rect 17195 -6289 17207 -6255
rect 17241 -6289 17253 -6255
rect 17195 -6323 17253 -6289
rect 17195 -6357 17207 -6323
rect 17241 -6357 17253 -6323
rect 17195 -6391 17253 -6357
rect 17195 -6425 17207 -6391
rect 17241 -6425 17253 -6391
rect 17195 -6440 17253 -6425
rect 17453 -6255 17511 -6240
rect 17453 -6289 17465 -6255
rect 17499 -6289 17511 -6255
rect 17453 -6323 17511 -6289
rect 17453 -6357 17465 -6323
rect 17499 -6357 17511 -6323
rect 17453 -6391 17511 -6357
rect 17453 -6425 17465 -6391
rect 17499 -6425 17511 -6391
rect 17453 -6440 17511 -6425
rect 17711 -6255 17769 -6240
rect 17711 -6289 17723 -6255
rect 17757 -6289 17769 -6255
rect 17711 -6323 17769 -6289
rect 17711 -6357 17723 -6323
rect 17757 -6357 17769 -6323
rect 17711 -6391 17769 -6357
rect 17711 -6425 17723 -6391
rect 17757 -6425 17769 -6391
rect 17711 -6440 17769 -6425
rect 17905 -6255 17963 -6240
rect 17905 -6289 17917 -6255
rect 17951 -6289 17963 -6255
rect 17905 -6323 17963 -6289
rect 17905 -6357 17917 -6323
rect 17951 -6357 17963 -6323
rect 17905 -6391 17963 -6357
rect 17905 -6425 17917 -6391
rect 17951 -6425 17963 -6391
rect 17905 -6440 17963 -6425
rect 18163 -6255 18221 -6240
rect 18163 -6289 18175 -6255
rect 18209 -6289 18221 -6255
rect 18163 -6323 18221 -6289
rect 18163 -6357 18175 -6323
rect 18209 -6357 18221 -6323
rect 18163 -6391 18221 -6357
rect 18163 -6425 18175 -6391
rect 18209 -6425 18221 -6391
rect 18163 -6440 18221 -6425
rect 959 -7212 1017 -7197
rect 959 -7246 971 -7212
rect 1005 -7246 1017 -7212
rect 959 -7280 1017 -7246
rect 959 -7314 971 -7280
rect 1005 -7314 1017 -7280
rect 959 -7348 1017 -7314
rect 959 -7382 971 -7348
rect 1005 -7382 1017 -7348
rect 959 -7397 1017 -7382
rect 1217 -7212 1275 -7197
rect 1217 -7246 1229 -7212
rect 1263 -7246 1275 -7212
rect 1217 -7280 1275 -7246
rect 1217 -7314 1229 -7280
rect 1263 -7314 1275 -7280
rect 1217 -7348 1275 -7314
rect 1217 -7382 1229 -7348
rect 1263 -7382 1275 -7348
rect 1217 -7397 1275 -7382
rect 1411 -7212 1469 -7197
rect 1411 -7246 1423 -7212
rect 1457 -7246 1469 -7212
rect 1411 -7280 1469 -7246
rect 1411 -7314 1423 -7280
rect 1457 -7314 1469 -7280
rect 1411 -7348 1469 -7314
rect 1411 -7382 1423 -7348
rect 1457 -7382 1469 -7348
rect 1411 -7397 1469 -7382
rect 1669 -7212 1727 -7197
rect 1669 -7246 1681 -7212
rect 1715 -7246 1727 -7212
rect 1669 -7280 1727 -7246
rect 1669 -7314 1681 -7280
rect 1715 -7314 1727 -7280
rect 1669 -7348 1727 -7314
rect 1669 -7382 1681 -7348
rect 1715 -7382 1727 -7348
rect 1669 -7397 1727 -7382
rect 1927 -7212 1985 -7197
rect 1927 -7246 1939 -7212
rect 1973 -7246 1985 -7212
rect 1927 -7280 1985 -7246
rect 1927 -7314 1939 -7280
rect 1973 -7314 1985 -7280
rect 1927 -7348 1985 -7314
rect 1927 -7382 1939 -7348
rect 1973 -7382 1985 -7348
rect 1927 -7397 1985 -7382
rect 2185 -7212 2243 -7197
rect 2185 -7246 2197 -7212
rect 2231 -7246 2243 -7212
rect 2185 -7280 2243 -7246
rect 2185 -7314 2197 -7280
rect 2231 -7314 2243 -7280
rect 2185 -7348 2243 -7314
rect 2185 -7382 2197 -7348
rect 2231 -7382 2243 -7348
rect 2185 -7397 2243 -7382
rect 2443 -7212 2501 -7197
rect 2443 -7246 2455 -7212
rect 2489 -7246 2501 -7212
rect 2443 -7280 2501 -7246
rect 2443 -7314 2455 -7280
rect 2489 -7314 2501 -7280
rect 2443 -7348 2501 -7314
rect 2443 -7382 2455 -7348
rect 2489 -7382 2501 -7348
rect 2443 -7397 2501 -7382
rect 2637 -7212 2695 -7197
rect 2637 -7246 2649 -7212
rect 2683 -7246 2695 -7212
rect 2637 -7280 2695 -7246
rect 2637 -7314 2649 -7280
rect 2683 -7314 2695 -7280
rect 2637 -7348 2695 -7314
rect 2637 -7382 2649 -7348
rect 2683 -7382 2695 -7348
rect 2637 -7397 2695 -7382
rect 2895 -7212 2953 -7197
rect 2895 -7246 2907 -7212
rect 2941 -7246 2953 -7212
rect 2895 -7280 2953 -7246
rect 2895 -7314 2907 -7280
rect 2941 -7314 2953 -7280
rect 2895 -7348 2953 -7314
rect 2895 -7382 2907 -7348
rect 2941 -7382 2953 -7348
rect 2895 -7397 2953 -7382
rect 3153 -7212 3211 -7197
rect 3153 -7246 3165 -7212
rect 3199 -7246 3211 -7212
rect 3153 -7280 3211 -7246
rect 3153 -7314 3165 -7280
rect 3199 -7314 3211 -7280
rect 3153 -7348 3211 -7314
rect 3153 -7382 3165 -7348
rect 3199 -7382 3211 -7348
rect 3153 -7397 3211 -7382
rect 3411 -7212 3469 -7197
rect 3411 -7246 3423 -7212
rect 3457 -7246 3469 -7212
rect 3411 -7280 3469 -7246
rect 3411 -7314 3423 -7280
rect 3457 -7314 3469 -7280
rect 3411 -7348 3469 -7314
rect 3411 -7382 3423 -7348
rect 3457 -7382 3469 -7348
rect 3411 -7397 3469 -7382
rect 3605 -7212 3663 -7197
rect 3605 -7246 3617 -7212
rect 3651 -7246 3663 -7212
rect 3605 -7280 3663 -7246
rect 3605 -7314 3617 -7280
rect 3651 -7314 3663 -7280
rect 3605 -7348 3663 -7314
rect 3605 -7382 3617 -7348
rect 3651 -7382 3663 -7348
rect 3605 -7397 3663 -7382
rect 3863 -7212 3921 -7197
rect 3863 -7246 3875 -7212
rect 3909 -7246 3921 -7212
rect 3863 -7280 3921 -7246
rect 3863 -7314 3875 -7280
rect 3909 -7314 3921 -7280
rect 3863 -7348 3921 -7314
rect 3863 -7382 3875 -7348
rect 3909 -7382 3921 -7348
rect 3863 -7397 3921 -7382
rect 4121 -7212 4179 -7197
rect 4121 -7246 4133 -7212
rect 4167 -7246 4179 -7212
rect 4121 -7280 4179 -7246
rect 4121 -7314 4133 -7280
rect 4167 -7314 4179 -7280
rect 4121 -7348 4179 -7314
rect 4121 -7382 4133 -7348
rect 4167 -7382 4179 -7348
rect 4121 -7397 4179 -7382
rect 4379 -7212 4437 -7197
rect 4379 -7246 4391 -7212
rect 4425 -7246 4437 -7212
rect 4379 -7280 4437 -7246
rect 4379 -7314 4391 -7280
rect 4425 -7314 4437 -7280
rect 4379 -7348 4437 -7314
rect 4379 -7382 4391 -7348
rect 4425 -7382 4437 -7348
rect 4379 -7397 4437 -7382
rect 4637 -7212 4695 -7197
rect 4637 -7246 4649 -7212
rect 4683 -7246 4695 -7212
rect 4637 -7280 4695 -7246
rect 4637 -7314 4649 -7280
rect 4683 -7314 4695 -7280
rect 4637 -7348 4695 -7314
rect 4637 -7382 4649 -7348
rect 4683 -7382 4695 -7348
rect 4637 -7397 4695 -7382
rect 4830 -7212 4888 -7197
rect 4830 -7246 4842 -7212
rect 4876 -7246 4888 -7212
rect 4830 -7280 4888 -7246
rect 4830 -7314 4842 -7280
rect 4876 -7314 4888 -7280
rect 4830 -7348 4888 -7314
rect 4830 -7382 4842 -7348
rect 4876 -7382 4888 -7348
rect 4830 -7397 4888 -7382
rect 5088 -7212 5146 -7197
rect 5088 -7246 5100 -7212
rect 5134 -7246 5146 -7212
rect 5088 -7280 5146 -7246
rect 5088 -7314 5100 -7280
rect 5134 -7314 5146 -7280
rect 5088 -7348 5146 -7314
rect 5088 -7382 5100 -7348
rect 5134 -7382 5146 -7348
rect 5088 -7397 5146 -7382
rect 5316 -7212 5374 -7197
rect 5316 -7246 5328 -7212
rect 5362 -7246 5374 -7212
rect 5316 -7280 5374 -7246
rect 5316 -7314 5328 -7280
rect 5362 -7314 5374 -7280
rect 5316 -7348 5374 -7314
rect 5316 -7382 5328 -7348
rect 5362 -7382 5374 -7348
rect 5316 -7397 5374 -7382
rect 5574 -7212 5632 -7197
rect 5574 -7246 5586 -7212
rect 5620 -7246 5632 -7212
rect 5574 -7280 5632 -7246
rect 5574 -7314 5586 -7280
rect 5620 -7314 5632 -7280
rect 5574 -7348 5632 -7314
rect 5574 -7382 5586 -7348
rect 5620 -7382 5632 -7348
rect 5574 -7397 5632 -7382
rect 5768 -7212 5826 -7197
rect 5768 -7246 5780 -7212
rect 5814 -7246 5826 -7212
rect 5768 -7280 5826 -7246
rect 5768 -7314 5780 -7280
rect 5814 -7314 5826 -7280
rect 5768 -7348 5826 -7314
rect 5768 -7382 5780 -7348
rect 5814 -7382 5826 -7348
rect 5768 -7397 5826 -7382
rect 6026 -7212 6084 -7197
rect 6026 -7246 6038 -7212
rect 6072 -7246 6084 -7212
rect 6026 -7280 6084 -7246
rect 6026 -7314 6038 -7280
rect 6072 -7314 6084 -7280
rect 6026 -7348 6084 -7314
rect 6026 -7382 6038 -7348
rect 6072 -7382 6084 -7348
rect 6026 -7397 6084 -7382
rect 6284 -7212 6342 -7197
rect 6284 -7246 6296 -7212
rect 6330 -7246 6342 -7212
rect 6284 -7280 6342 -7246
rect 6284 -7314 6296 -7280
rect 6330 -7314 6342 -7280
rect 6284 -7348 6342 -7314
rect 6284 -7382 6296 -7348
rect 6330 -7382 6342 -7348
rect 6284 -7397 6342 -7382
rect 6542 -7212 6600 -7197
rect 6542 -7246 6554 -7212
rect 6588 -7246 6600 -7212
rect 6542 -7280 6600 -7246
rect 6542 -7314 6554 -7280
rect 6588 -7314 6600 -7280
rect 6542 -7348 6600 -7314
rect 6542 -7382 6554 -7348
rect 6588 -7382 6600 -7348
rect 6542 -7397 6600 -7382
rect 6800 -7212 6858 -7197
rect 6800 -7246 6812 -7212
rect 6846 -7246 6858 -7212
rect 6800 -7280 6858 -7246
rect 6800 -7314 6812 -7280
rect 6846 -7314 6858 -7280
rect 6800 -7348 6858 -7314
rect 6800 -7382 6812 -7348
rect 6846 -7382 6858 -7348
rect 6800 -7397 6858 -7382
rect 6994 -7212 7052 -7197
rect 6994 -7246 7006 -7212
rect 7040 -7246 7052 -7212
rect 6994 -7280 7052 -7246
rect 6994 -7314 7006 -7280
rect 7040 -7314 7052 -7280
rect 6994 -7348 7052 -7314
rect 6994 -7382 7006 -7348
rect 7040 -7382 7052 -7348
rect 6994 -7397 7052 -7382
rect 7252 -7212 7310 -7197
rect 7252 -7246 7264 -7212
rect 7298 -7246 7310 -7212
rect 7252 -7280 7310 -7246
rect 7252 -7314 7264 -7280
rect 7298 -7314 7310 -7280
rect 7252 -7348 7310 -7314
rect 7252 -7382 7264 -7348
rect 7298 -7382 7310 -7348
rect 7252 -7397 7310 -7382
rect 7510 -7212 7568 -7197
rect 7510 -7246 7522 -7212
rect 7556 -7246 7568 -7212
rect 7510 -7280 7568 -7246
rect 7510 -7314 7522 -7280
rect 7556 -7314 7568 -7280
rect 7510 -7348 7568 -7314
rect 7510 -7382 7522 -7348
rect 7556 -7382 7568 -7348
rect 7510 -7397 7568 -7382
rect 7768 -7212 7826 -7197
rect 7768 -7246 7780 -7212
rect 7814 -7246 7826 -7212
rect 7768 -7280 7826 -7246
rect 7768 -7314 7780 -7280
rect 7814 -7314 7826 -7280
rect 7768 -7348 7826 -7314
rect 7768 -7382 7780 -7348
rect 7814 -7382 7826 -7348
rect 7768 -7397 7826 -7382
rect 7962 -7212 8020 -7197
rect 7962 -7246 7974 -7212
rect 8008 -7246 8020 -7212
rect 7962 -7280 8020 -7246
rect 7962 -7314 7974 -7280
rect 8008 -7314 8020 -7280
rect 7962 -7348 8020 -7314
rect 7962 -7382 7974 -7348
rect 8008 -7382 8020 -7348
rect 7962 -7397 8020 -7382
rect 8220 -7212 8278 -7197
rect 8220 -7246 8232 -7212
rect 8266 -7246 8278 -7212
rect 8220 -7280 8278 -7246
rect 8220 -7314 8232 -7280
rect 8266 -7314 8278 -7280
rect 8220 -7348 8278 -7314
rect 8220 -7382 8232 -7348
rect 8266 -7382 8278 -7348
rect 8220 -7397 8278 -7382
rect 8478 -7212 8536 -7197
rect 8478 -7246 8490 -7212
rect 8524 -7246 8536 -7212
rect 8478 -7280 8536 -7246
rect 8478 -7314 8490 -7280
rect 8524 -7314 8536 -7280
rect 8478 -7348 8536 -7314
rect 8478 -7382 8490 -7348
rect 8524 -7382 8536 -7348
rect 8478 -7397 8536 -7382
rect 8736 -7212 8794 -7197
rect 8736 -7246 8748 -7212
rect 8782 -7246 8794 -7212
rect 8736 -7280 8794 -7246
rect 8736 -7314 8748 -7280
rect 8782 -7314 8794 -7280
rect 8736 -7348 8794 -7314
rect 8736 -7382 8748 -7348
rect 8782 -7382 8794 -7348
rect 8736 -7397 8794 -7382
rect 8994 -7212 9052 -7197
rect 8994 -7246 9006 -7212
rect 9040 -7246 9052 -7212
rect 8994 -7280 9052 -7246
rect 8994 -7314 9006 -7280
rect 9040 -7314 9052 -7280
rect 8994 -7348 9052 -7314
rect 8994 -7382 9006 -7348
rect 9040 -7382 9052 -7348
rect 8994 -7397 9052 -7382
rect 9188 -7212 9246 -7197
rect 9188 -7246 9200 -7212
rect 9234 -7246 9246 -7212
rect 9188 -7280 9246 -7246
rect 9188 -7314 9200 -7280
rect 9234 -7314 9246 -7280
rect 9188 -7348 9246 -7314
rect 9188 -7382 9200 -7348
rect 9234 -7382 9246 -7348
rect 9188 -7397 9246 -7382
rect 9446 -7212 9504 -7197
rect 9446 -7246 9458 -7212
rect 9492 -7246 9504 -7212
rect 9446 -7280 9504 -7246
rect 9446 -7314 9458 -7280
rect 9492 -7314 9504 -7280
rect 9446 -7348 9504 -7314
rect 9446 -7382 9458 -7348
rect 9492 -7382 9504 -7348
rect 9446 -7397 9504 -7382
rect 9676 -7212 9734 -7197
rect 9676 -7246 9688 -7212
rect 9722 -7246 9734 -7212
rect 9676 -7280 9734 -7246
rect 9676 -7314 9688 -7280
rect 9722 -7314 9734 -7280
rect 9676 -7348 9734 -7314
rect 9676 -7382 9688 -7348
rect 9722 -7382 9734 -7348
rect 9676 -7397 9734 -7382
rect 9934 -7212 9992 -7197
rect 9934 -7246 9946 -7212
rect 9980 -7246 9992 -7212
rect 9934 -7280 9992 -7246
rect 9934 -7314 9946 -7280
rect 9980 -7314 9992 -7280
rect 9934 -7348 9992 -7314
rect 9934 -7382 9946 -7348
rect 9980 -7382 9992 -7348
rect 9934 -7397 9992 -7382
rect 10128 -7212 10186 -7197
rect 10128 -7246 10140 -7212
rect 10174 -7246 10186 -7212
rect 10128 -7280 10186 -7246
rect 10128 -7314 10140 -7280
rect 10174 -7314 10186 -7280
rect 10128 -7348 10186 -7314
rect 10128 -7382 10140 -7348
rect 10174 -7382 10186 -7348
rect 10128 -7397 10186 -7382
rect 10386 -7212 10444 -7197
rect 10386 -7246 10398 -7212
rect 10432 -7246 10444 -7212
rect 10386 -7280 10444 -7246
rect 10386 -7314 10398 -7280
rect 10432 -7314 10444 -7280
rect 10386 -7348 10444 -7314
rect 10386 -7382 10398 -7348
rect 10432 -7382 10444 -7348
rect 10386 -7397 10444 -7382
rect 10644 -7212 10702 -7197
rect 10644 -7246 10656 -7212
rect 10690 -7246 10702 -7212
rect 10644 -7280 10702 -7246
rect 10644 -7314 10656 -7280
rect 10690 -7314 10702 -7280
rect 10644 -7348 10702 -7314
rect 10644 -7382 10656 -7348
rect 10690 -7382 10702 -7348
rect 10644 -7397 10702 -7382
rect 10902 -7212 10960 -7197
rect 10902 -7246 10914 -7212
rect 10948 -7246 10960 -7212
rect 10902 -7280 10960 -7246
rect 10902 -7314 10914 -7280
rect 10948 -7314 10960 -7280
rect 10902 -7348 10960 -7314
rect 10902 -7382 10914 -7348
rect 10948 -7382 10960 -7348
rect 10902 -7397 10960 -7382
rect 11160 -7212 11218 -7197
rect 11160 -7246 11172 -7212
rect 11206 -7246 11218 -7212
rect 11160 -7280 11218 -7246
rect 11160 -7314 11172 -7280
rect 11206 -7314 11218 -7280
rect 11160 -7348 11218 -7314
rect 11160 -7382 11172 -7348
rect 11206 -7382 11218 -7348
rect 11160 -7397 11218 -7382
rect 11354 -7212 11412 -7197
rect 11354 -7246 11366 -7212
rect 11400 -7246 11412 -7212
rect 11354 -7280 11412 -7246
rect 11354 -7314 11366 -7280
rect 11400 -7314 11412 -7280
rect 11354 -7348 11412 -7314
rect 11354 -7382 11366 -7348
rect 11400 -7382 11412 -7348
rect 11354 -7397 11412 -7382
rect 11612 -7212 11670 -7197
rect 11612 -7246 11624 -7212
rect 11658 -7246 11670 -7212
rect 11612 -7280 11670 -7246
rect 11612 -7314 11624 -7280
rect 11658 -7314 11670 -7280
rect 11612 -7348 11670 -7314
rect 11612 -7382 11624 -7348
rect 11658 -7382 11670 -7348
rect 11612 -7397 11670 -7382
rect 11870 -7212 11928 -7197
rect 11870 -7246 11882 -7212
rect 11916 -7246 11928 -7212
rect 11870 -7280 11928 -7246
rect 11870 -7314 11882 -7280
rect 11916 -7314 11928 -7280
rect 11870 -7348 11928 -7314
rect 11870 -7382 11882 -7348
rect 11916 -7382 11928 -7348
rect 11870 -7397 11928 -7382
rect 12128 -7212 12186 -7197
rect 12128 -7246 12140 -7212
rect 12174 -7246 12186 -7212
rect 12128 -7280 12186 -7246
rect 12128 -7314 12140 -7280
rect 12174 -7314 12186 -7280
rect 12128 -7348 12186 -7314
rect 12128 -7382 12140 -7348
rect 12174 -7382 12186 -7348
rect 12128 -7397 12186 -7382
rect 12322 -7212 12380 -7197
rect 12322 -7246 12334 -7212
rect 12368 -7246 12380 -7212
rect 12322 -7280 12380 -7246
rect 12322 -7314 12334 -7280
rect 12368 -7314 12380 -7280
rect 12322 -7348 12380 -7314
rect 12322 -7382 12334 -7348
rect 12368 -7382 12380 -7348
rect 12322 -7397 12380 -7382
rect 12580 -7212 12638 -7197
rect 12580 -7246 12592 -7212
rect 12626 -7246 12638 -7212
rect 12580 -7280 12638 -7246
rect 12580 -7314 12592 -7280
rect 12626 -7314 12638 -7280
rect 12580 -7348 12638 -7314
rect 12580 -7382 12592 -7348
rect 12626 -7382 12638 -7348
rect 12580 -7397 12638 -7382
rect 12838 -7212 12896 -7197
rect 12838 -7246 12850 -7212
rect 12884 -7246 12896 -7212
rect 12838 -7280 12896 -7246
rect 12838 -7314 12850 -7280
rect 12884 -7314 12896 -7280
rect 12838 -7348 12896 -7314
rect 12838 -7382 12850 -7348
rect 12884 -7382 12896 -7348
rect 12838 -7397 12896 -7382
rect 13096 -7212 13154 -7197
rect 13096 -7246 13108 -7212
rect 13142 -7246 13154 -7212
rect 13096 -7280 13154 -7246
rect 13096 -7314 13108 -7280
rect 13142 -7314 13154 -7280
rect 13096 -7348 13154 -7314
rect 13096 -7382 13108 -7348
rect 13142 -7382 13154 -7348
rect 13096 -7397 13154 -7382
rect 13354 -7212 13412 -7197
rect 13354 -7246 13366 -7212
rect 13400 -7246 13412 -7212
rect 13354 -7280 13412 -7246
rect 13354 -7314 13366 -7280
rect 13400 -7314 13412 -7280
rect 13354 -7348 13412 -7314
rect 13354 -7382 13366 -7348
rect 13400 -7382 13412 -7348
rect 13354 -7397 13412 -7382
rect 13548 -7212 13606 -7197
rect 13548 -7246 13560 -7212
rect 13594 -7246 13606 -7212
rect 13548 -7280 13606 -7246
rect 13548 -7314 13560 -7280
rect 13594 -7314 13606 -7280
rect 13548 -7348 13606 -7314
rect 13548 -7382 13560 -7348
rect 13594 -7382 13606 -7348
rect 13548 -7397 13606 -7382
rect 13806 -7212 13864 -7197
rect 13806 -7246 13818 -7212
rect 13852 -7246 13864 -7212
rect 13806 -7280 13864 -7246
rect 13806 -7314 13818 -7280
rect 13852 -7314 13864 -7280
rect 13806 -7348 13864 -7314
rect 13806 -7382 13818 -7348
rect 13852 -7382 13864 -7348
rect 13806 -7397 13864 -7382
rect 14034 -7212 14092 -7197
rect 14034 -7246 14046 -7212
rect 14080 -7246 14092 -7212
rect 14034 -7280 14092 -7246
rect 14034 -7314 14046 -7280
rect 14080 -7314 14092 -7280
rect 14034 -7348 14092 -7314
rect 14034 -7382 14046 -7348
rect 14080 -7382 14092 -7348
rect 14034 -7397 14092 -7382
rect 14292 -7212 14350 -7197
rect 14292 -7246 14304 -7212
rect 14338 -7246 14350 -7212
rect 14292 -7280 14350 -7246
rect 14292 -7314 14304 -7280
rect 14338 -7314 14350 -7280
rect 14292 -7348 14350 -7314
rect 14292 -7382 14304 -7348
rect 14338 -7382 14350 -7348
rect 14292 -7397 14350 -7382
rect 14485 -7212 14543 -7197
rect 14485 -7246 14497 -7212
rect 14531 -7246 14543 -7212
rect 14485 -7280 14543 -7246
rect 14485 -7314 14497 -7280
rect 14531 -7314 14543 -7280
rect 14485 -7348 14543 -7314
rect 14485 -7382 14497 -7348
rect 14531 -7382 14543 -7348
rect 14485 -7397 14543 -7382
rect 14743 -7212 14801 -7197
rect 14743 -7246 14755 -7212
rect 14789 -7246 14801 -7212
rect 14743 -7280 14801 -7246
rect 14743 -7314 14755 -7280
rect 14789 -7314 14801 -7280
rect 14743 -7348 14801 -7314
rect 14743 -7382 14755 -7348
rect 14789 -7382 14801 -7348
rect 14743 -7397 14801 -7382
rect 15001 -7212 15059 -7197
rect 15001 -7246 15013 -7212
rect 15047 -7246 15059 -7212
rect 15001 -7280 15059 -7246
rect 15001 -7314 15013 -7280
rect 15047 -7314 15059 -7280
rect 15001 -7348 15059 -7314
rect 15001 -7382 15013 -7348
rect 15047 -7382 15059 -7348
rect 15001 -7397 15059 -7382
rect 15259 -7212 15317 -7197
rect 15259 -7246 15271 -7212
rect 15305 -7246 15317 -7212
rect 15259 -7280 15317 -7246
rect 15259 -7314 15271 -7280
rect 15305 -7314 15317 -7280
rect 15259 -7348 15317 -7314
rect 15259 -7382 15271 -7348
rect 15305 -7382 15317 -7348
rect 15259 -7397 15317 -7382
rect 15517 -7212 15575 -7197
rect 15517 -7246 15529 -7212
rect 15563 -7246 15575 -7212
rect 15517 -7280 15575 -7246
rect 15517 -7314 15529 -7280
rect 15563 -7314 15575 -7280
rect 15517 -7348 15575 -7314
rect 15517 -7382 15529 -7348
rect 15563 -7382 15575 -7348
rect 15517 -7397 15575 -7382
rect 15711 -7212 15769 -7197
rect 15711 -7246 15723 -7212
rect 15757 -7246 15769 -7212
rect 15711 -7280 15769 -7246
rect 15711 -7314 15723 -7280
rect 15757 -7314 15769 -7280
rect 15711 -7348 15769 -7314
rect 15711 -7382 15723 -7348
rect 15757 -7382 15769 -7348
rect 15711 -7397 15769 -7382
rect 15969 -7212 16027 -7197
rect 15969 -7246 15981 -7212
rect 16015 -7246 16027 -7212
rect 15969 -7280 16027 -7246
rect 15969 -7314 15981 -7280
rect 16015 -7314 16027 -7280
rect 15969 -7348 16027 -7314
rect 15969 -7382 15981 -7348
rect 16015 -7382 16027 -7348
rect 15969 -7397 16027 -7382
rect 16227 -7212 16285 -7197
rect 16227 -7246 16239 -7212
rect 16273 -7246 16285 -7212
rect 16227 -7280 16285 -7246
rect 16227 -7314 16239 -7280
rect 16273 -7314 16285 -7280
rect 16227 -7348 16285 -7314
rect 16227 -7382 16239 -7348
rect 16273 -7382 16285 -7348
rect 16227 -7397 16285 -7382
rect 16485 -7212 16543 -7197
rect 16485 -7246 16497 -7212
rect 16531 -7246 16543 -7212
rect 16485 -7280 16543 -7246
rect 16485 -7314 16497 -7280
rect 16531 -7314 16543 -7280
rect 16485 -7348 16543 -7314
rect 16485 -7382 16497 -7348
rect 16531 -7382 16543 -7348
rect 16485 -7397 16543 -7382
rect 16679 -7212 16737 -7197
rect 16679 -7246 16691 -7212
rect 16725 -7246 16737 -7212
rect 16679 -7280 16737 -7246
rect 16679 -7314 16691 -7280
rect 16725 -7314 16737 -7280
rect 16679 -7348 16737 -7314
rect 16679 -7382 16691 -7348
rect 16725 -7382 16737 -7348
rect 16679 -7397 16737 -7382
rect 16937 -7212 16995 -7197
rect 16937 -7246 16949 -7212
rect 16983 -7246 16995 -7212
rect 16937 -7280 16995 -7246
rect 16937 -7314 16949 -7280
rect 16983 -7314 16995 -7280
rect 16937 -7348 16995 -7314
rect 16937 -7382 16949 -7348
rect 16983 -7382 16995 -7348
rect 16937 -7397 16995 -7382
rect 17195 -7212 17253 -7197
rect 17195 -7246 17207 -7212
rect 17241 -7246 17253 -7212
rect 17195 -7280 17253 -7246
rect 17195 -7314 17207 -7280
rect 17241 -7314 17253 -7280
rect 17195 -7348 17253 -7314
rect 17195 -7382 17207 -7348
rect 17241 -7382 17253 -7348
rect 17195 -7397 17253 -7382
rect 17453 -7212 17511 -7197
rect 17453 -7246 17465 -7212
rect 17499 -7246 17511 -7212
rect 17453 -7280 17511 -7246
rect 17453 -7314 17465 -7280
rect 17499 -7314 17511 -7280
rect 17453 -7348 17511 -7314
rect 17453 -7382 17465 -7348
rect 17499 -7382 17511 -7348
rect 17453 -7397 17511 -7382
rect 17711 -7212 17769 -7197
rect 17711 -7246 17723 -7212
rect 17757 -7246 17769 -7212
rect 17711 -7280 17769 -7246
rect 17711 -7314 17723 -7280
rect 17757 -7314 17769 -7280
rect 17711 -7348 17769 -7314
rect 17711 -7382 17723 -7348
rect 17757 -7382 17769 -7348
rect 17711 -7397 17769 -7382
rect 17905 -7212 17963 -7197
rect 17905 -7246 17917 -7212
rect 17951 -7246 17963 -7212
rect 17905 -7280 17963 -7246
rect 17905 -7314 17917 -7280
rect 17951 -7314 17963 -7280
rect 17905 -7348 17963 -7314
rect 17905 -7382 17917 -7348
rect 17951 -7382 17963 -7348
rect 17905 -7397 17963 -7382
rect 18163 -7212 18221 -7197
rect 18163 -7246 18175 -7212
rect 18209 -7246 18221 -7212
rect 18163 -7280 18221 -7246
rect 18163 -7314 18175 -7280
rect 18209 -7314 18221 -7280
rect 18163 -7348 18221 -7314
rect 18163 -7382 18175 -7348
rect 18209 -7382 18221 -7348
rect 18163 -7397 18221 -7382
rect 959 -7902 1017 -7887
rect 959 -7936 971 -7902
rect 1005 -7936 1017 -7902
rect 959 -7970 1017 -7936
rect 959 -8004 971 -7970
rect 1005 -8004 1017 -7970
rect 959 -8038 1017 -8004
rect 959 -8072 971 -8038
rect 1005 -8072 1017 -8038
rect 959 -8087 1017 -8072
rect 1217 -7902 1275 -7887
rect 1217 -7936 1229 -7902
rect 1263 -7936 1275 -7902
rect 1217 -7970 1275 -7936
rect 1217 -8004 1229 -7970
rect 1263 -8004 1275 -7970
rect 1217 -8038 1275 -8004
rect 1217 -8072 1229 -8038
rect 1263 -8072 1275 -8038
rect 1217 -8087 1275 -8072
rect 1411 -7902 1469 -7887
rect 1411 -7936 1423 -7902
rect 1457 -7936 1469 -7902
rect 1411 -7970 1469 -7936
rect 1411 -8004 1423 -7970
rect 1457 -8004 1469 -7970
rect 1411 -8038 1469 -8004
rect 1411 -8072 1423 -8038
rect 1457 -8072 1469 -8038
rect 1411 -8087 1469 -8072
rect 1669 -7902 1727 -7887
rect 1669 -7936 1681 -7902
rect 1715 -7936 1727 -7902
rect 1669 -7970 1727 -7936
rect 1669 -8004 1681 -7970
rect 1715 -8004 1727 -7970
rect 1669 -8038 1727 -8004
rect 1669 -8072 1681 -8038
rect 1715 -8072 1727 -8038
rect 1669 -8087 1727 -8072
rect 1927 -7902 1985 -7887
rect 1927 -7936 1939 -7902
rect 1973 -7936 1985 -7902
rect 1927 -7970 1985 -7936
rect 1927 -8004 1939 -7970
rect 1973 -8004 1985 -7970
rect 1927 -8038 1985 -8004
rect 1927 -8072 1939 -8038
rect 1973 -8072 1985 -8038
rect 1927 -8087 1985 -8072
rect 2185 -7902 2243 -7887
rect 2185 -7936 2197 -7902
rect 2231 -7936 2243 -7902
rect 2185 -7970 2243 -7936
rect 2185 -8004 2197 -7970
rect 2231 -8004 2243 -7970
rect 2185 -8038 2243 -8004
rect 2185 -8072 2197 -8038
rect 2231 -8072 2243 -8038
rect 2185 -8087 2243 -8072
rect 2443 -7902 2501 -7887
rect 2443 -7936 2455 -7902
rect 2489 -7936 2501 -7902
rect 2443 -7970 2501 -7936
rect 2443 -8004 2455 -7970
rect 2489 -8004 2501 -7970
rect 2443 -8038 2501 -8004
rect 2443 -8072 2455 -8038
rect 2489 -8072 2501 -8038
rect 2443 -8087 2501 -8072
rect 2637 -7902 2695 -7887
rect 2637 -7936 2649 -7902
rect 2683 -7936 2695 -7902
rect 2637 -7970 2695 -7936
rect 2637 -8004 2649 -7970
rect 2683 -8004 2695 -7970
rect 2637 -8038 2695 -8004
rect 2637 -8072 2649 -8038
rect 2683 -8072 2695 -8038
rect 2637 -8087 2695 -8072
rect 2895 -7902 2953 -7887
rect 2895 -7936 2907 -7902
rect 2941 -7936 2953 -7902
rect 2895 -7970 2953 -7936
rect 2895 -8004 2907 -7970
rect 2941 -8004 2953 -7970
rect 2895 -8038 2953 -8004
rect 2895 -8072 2907 -8038
rect 2941 -8072 2953 -8038
rect 2895 -8087 2953 -8072
rect 3153 -7902 3211 -7887
rect 3153 -7936 3165 -7902
rect 3199 -7936 3211 -7902
rect 3153 -7970 3211 -7936
rect 3153 -8004 3165 -7970
rect 3199 -8004 3211 -7970
rect 3153 -8038 3211 -8004
rect 3153 -8072 3165 -8038
rect 3199 -8072 3211 -8038
rect 3153 -8087 3211 -8072
rect 3411 -7902 3469 -7887
rect 3411 -7936 3423 -7902
rect 3457 -7936 3469 -7902
rect 3411 -7970 3469 -7936
rect 3411 -8004 3423 -7970
rect 3457 -8004 3469 -7970
rect 3411 -8038 3469 -8004
rect 3411 -8072 3423 -8038
rect 3457 -8072 3469 -8038
rect 3411 -8087 3469 -8072
rect 3605 -7902 3663 -7887
rect 3605 -7936 3617 -7902
rect 3651 -7936 3663 -7902
rect 3605 -7970 3663 -7936
rect 3605 -8004 3617 -7970
rect 3651 -8004 3663 -7970
rect 3605 -8038 3663 -8004
rect 3605 -8072 3617 -8038
rect 3651 -8072 3663 -8038
rect 3605 -8087 3663 -8072
rect 3863 -7902 3921 -7887
rect 3863 -7936 3875 -7902
rect 3909 -7936 3921 -7902
rect 3863 -7970 3921 -7936
rect 3863 -8004 3875 -7970
rect 3909 -8004 3921 -7970
rect 3863 -8038 3921 -8004
rect 3863 -8072 3875 -8038
rect 3909 -8072 3921 -8038
rect 3863 -8087 3921 -8072
rect 4121 -7902 4179 -7887
rect 4121 -7936 4133 -7902
rect 4167 -7936 4179 -7902
rect 4121 -7970 4179 -7936
rect 4121 -8004 4133 -7970
rect 4167 -8004 4179 -7970
rect 4121 -8038 4179 -8004
rect 4121 -8072 4133 -8038
rect 4167 -8072 4179 -8038
rect 4121 -8087 4179 -8072
rect 4379 -7902 4437 -7887
rect 4379 -7936 4391 -7902
rect 4425 -7936 4437 -7902
rect 4379 -7970 4437 -7936
rect 4379 -8004 4391 -7970
rect 4425 -8004 4437 -7970
rect 4379 -8038 4437 -8004
rect 4379 -8072 4391 -8038
rect 4425 -8072 4437 -8038
rect 4379 -8087 4437 -8072
rect 4637 -7902 4695 -7887
rect 4637 -7936 4649 -7902
rect 4683 -7936 4695 -7902
rect 4637 -7970 4695 -7936
rect 4637 -8004 4649 -7970
rect 4683 -8004 4695 -7970
rect 4637 -8038 4695 -8004
rect 4637 -8072 4649 -8038
rect 4683 -8072 4695 -8038
rect 4637 -8087 4695 -8072
rect 4830 -7902 4888 -7887
rect 4830 -7936 4842 -7902
rect 4876 -7936 4888 -7902
rect 4830 -7970 4888 -7936
rect 4830 -8004 4842 -7970
rect 4876 -8004 4888 -7970
rect 4830 -8038 4888 -8004
rect 4830 -8072 4842 -8038
rect 4876 -8072 4888 -8038
rect 4830 -8087 4888 -8072
rect 5088 -7902 5146 -7887
rect 5088 -7936 5100 -7902
rect 5134 -7936 5146 -7902
rect 5088 -7970 5146 -7936
rect 5088 -8004 5100 -7970
rect 5134 -8004 5146 -7970
rect 5088 -8038 5146 -8004
rect 5088 -8072 5100 -8038
rect 5134 -8072 5146 -8038
rect 5088 -8087 5146 -8072
rect 5316 -7902 5374 -7887
rect 5316 -7936 5328 -7902
rect 5362 -7936 5374 -7902
rect 5316 -7970 5374 -7936
rect 5316 -8004 5328 -7970
rect 5362 -8004 5374 -7970
rect 5316 -8038 5374 -8004
rect 5316 -8072 5328 -8038
rect 5362 -8072 5374 -8038
rect 5316 -8087 5374 -8072
rect 5574 -7902 5632 -7887
rect 5574 -7936 5586 -7902
rect 5620 -7936 5632 -7902
rect 5574 -7970 5632 -7936
rect 5574 -8004 5586 -7970
rect 5620 -8004 5632 -7970
rect 5574 -8038 5632 -8004
rect 5574 -8072 5586 -8038
rect 5620 -8072 5632 -8038
rect 5574 -8087 5632 -8072
rect 5768 -7902 5826 -7887
rect 5768 -7936 5780 -7902
rect 5814 -7936 5826 -7902
rect 5768 -7970 5826 -7936
rect 5768 -8004 5780 -7970
rect 5814 -8004 5826 -7970
rect 5768 -8038 5826 -8004
rect 5768 -8072 5780 -8038
rect 5814 -8072 5826 -8038
rect 5768 -8087 5826 -8072
rect 6026 -7902 6084 -7887
rect 6026 -7936 6038 -7902
rect 6072 -7936 6084 -7902
rect 6026 -7970 6084 -7936
rect 6026 -8004 6038 -7970
rect 6072 -8004 6084 -7970
rect 6026 -8038 6084 -8004
rect 6026 -8072 6038 -8038
rect 6072 -8072 6084 -8038
rect 6026 -8087 6084 -8072
rect 6284 -7902 6342 -7887
rect 6284 -7936 6296 -7902
rect 6330 -7936 6342 -7902
rect 6284 -7970 6342 -7936
rect 6284 -8004 6296 -7970
rect 6330 -8004 6342 -7970
rect 6284 -8038 6342 -8004
rect 6284 -8072 6296 -8038
rect 6330 -8072 6342 -8038
rect 6284 -8087 6342 -8072
rect 6542 -7902 6600 -7887
rect 6542 -7936 6554 -7902
rect 6588 -7936 6600 -7902
rect 6542 -7970 6600 -7936
rect 6542 -8004 6554 -7970
rect 6588 -8004 6600 -7970
rect 6542 -8038 6600 -8004
rect 6542 -8072 6554 -8038
rect 6588 -8072 6600 -8038
rect 6542 -8087 6600 -8072
rect 6800 -7902 6858 -7887
rect 6800 -7936 6812 -7902
rect 6846 -7936 6858 -7902
rect 6800 -7970 6858 -7936
rect 6800 -8004 6812 -7970
rect 6846 -8004 6858 -7970
rect 6800 -8038 6858 -8004
rect 6800 -8072 6812 -8038
rect 6846 -8072 6858 -8038
rect 6800 -8087 6858 -8072
rect 6994 -7902 7052 -7887
rect 6994 -7936 7006 -7902
rect 7040 -7936 7052 -7902
rect 6994 -7970 7052 -7936
rect 6994 -8004 7006 -7970
rect 7040 -8004 7052 -7970
rect 6994 -8038 7052 -8004
rect 6994 -8072 7006 -8038
rect 7040 -8072 7052 -8038
rect 6994 -8087 7052 -8072
rect 7252 -7902 7310 -7887
rect 7252 -7936 7264 -7902
rect 7298 -7936 7310 -7902
rect 7252 -7970 7310 -7936
rect 7252 -8004 7264 -7970
rect 7298 -8004 7310 -7970
rect 7252 -8038 7310 -8004
rect 7252 -8072 7264 -8038
rect 7298 -8072 7310 -8038
rect 7252 -8087 7310 -8072
rect 7510 -7902 7568 -7887
rect 7510 -7936 7522 -7902
rect 7556 -7936 7568 -7902
rect 7510 -7970 7568 -7936
rect 7510 -8004 7522 -7970
rect 7556 -8004 7568 -7970
rect 7510 -8038 7568 -8004
rect 7510 -8072 7522 -8038
rect 7556 -8072 7568 -8038
rect 7510 -8087 7568 -8072
rect 7768 -7902 7826 -7887
rect 7768 -7936 7780 -7902
rect 7814 -7936 7826 -7902
rect 7768 -7970 7826 -7936
rect 7768 -8004 7780 -7970
rect 7814 -8004 7826 -7970
rect 7768 -8038 7826 -8004
rect 7768 -8072 7780 -8038
rect 7814 -8072 7826 -8038
rect 7768 -8087 7826 -8072
rect 7962 -7902 8020 -7887
rect 7962 -7936 7974 -7902
rect 8008 -7936 8020 -7902
rect 7962 -7970 8020 -7936
rect 7962 -8004 7974 -7970
rect 8008 -8004 8020 -7970
rect 7962 -8038 8020 -8004
rect 7962 -8072 7974 -8038
rect 8008 -8072 8020 -8038
rect 7962 -8087 8020 -8072
rect 8220 -7902 8278 -7887
rect 8220 -7936 8232 -7902
rect 8266 -7936 8278 -7902
rect 8220 -7970 8278 -7936
rect 8220 -8004 8232 -7970
rect 8266 -8004 8278 -7970
rect 8220 -8038 8278 -8004
rect 8220 -8072 8232 -8038
rect 8266 -8072 8278 -8038
rect 8220 -8087 8278 -8072
rect 8478 -7902 8536 -7887
rect 8478 -7936 8490 -7902
rect 8524 -7936 8536 -7902
rect 8478 -7970 8536 -7936
rect 8478 -8004 8490 -7970
rect 8524 -8004 8536 -7970
rect 8478 -8038 8536 -8004
rect 8478 -8072 8490 -8038
rect 8524 -8072 8536 -8038
rect 8478 -8087 8536 -8072
rect 8736 -7902 8794 -7887
rect 8736 -7936 8748 -7902
rect 8782 -7936 8794 -7902
rect 8736 -7970 8794 -7936
rect 8736 -8004 8748 -7970
rect 8782 -8004 8794 -7970
rect 8736 -8038 8794 -8004
rect 8736 -8072 8748 -8038
rect 8782 -8072 8794 -8038
rect 8736 -8087 8794 -8072
rect 8994 -7902 9052 -7887
rect 8994 -7936 9006 -7902
rect 9040 -7936 9052 -7902
rect 8994 -7970 9052 -7936
rect 8994 -8004 9006 -7970
rect 9040 -8004 9052 -7970
rect 8994 -8038 9052 -8004
rect 8994 -8072 9006 -8038
rect 9040 -8072 9052 -8038
rect 8994 -8087 9052 -8072
rect 9188 -7902 9246 -7887
rect 9188 -7936 9200 -7902
rect 9234 -7936 9246 -7902
rect 9188 -7970 9246 -7936
rect 9188 -8004 9200 -7970
rect 9234 -8004 9246 -7970
rect 9188 -8038 9246 -8004
rect 9188 -8072 9200 -8038
rect 9234 -8072 9246 -8038
rect 9188 -8087 9246 -8072
rect 9446 -7902 9504 -7887
rect 9446 -7936 9458 -7902
rect 9492 -7936 9504 -7902
rect 9446 -7970 9504 -7936
rect 9446 -8004 9458 -7970
rect 9492 -8004 9504 -7970
rect 9446 -8038 9504 -8004
rect 9446 -8072 9458 -8038
rect 9492 -8072 9504 -8038
rect 9446 -8087 9504 -8072
rect 9676 -7902 9734 -7887
rect 9676 -7936 9688 -7902
rect 9722 -7936 9734 -7902
rect 9676 -7970 9734 -7936
rect 9676 -8004 9688 -7970
rect 9722 -8004 9734 -7970
rect 9676 -8038 9734 -8004
rect 9676 -8072 9688 -8038
rect 9722 -8072 9734 -8038
rect 9676 -8087 9734 -8072
rect 9934 -7902 9992 -7887
rect 9934 -7936 9946 -7902
rect 9980 -7936 9992 -7902
rect 9934 -7970 9992 -7936
rect 9934 -8004 9946 -7970
rect 9980 -8004 9992 -7970
rect 9934 -8038 9992 -8004
rect 9934 -8072 9946 -8038
rect 9980 -8072 9992 -8038
rect 9934 -8087 9992 -8072
rect 10128 -7902 10186 -7887
rect 10128 -7936 10140 -7902
rect 10174 -7936 10186 -7902
rect 10128 -7970 10186 -7936
rect 10128 -8004 10140 -7970
rect 10174 -8004 10186 -7970
rect 10128 -8038 10186 -8004
rect 10128 -8072 10140 -8038
rect 10174 -8072 10186 -8038
rect 10128 -8087 10186 -8072
rect 10386 -7902 10444 -7887
rect 10386 -7936 10398 -7902
rect 10432 -7936 10444 -7902
rect 10386 -7970 10444 -7936
rect 10386 -8004 10398 -7970
rect 10432 -8004 10444 -7970
rect 10386 -8038 10444 -8004
rect 10386 -8072 10398 -8038
rect 10432 -8072 10444 -8038
rect 10386 -8087 10444 -8072
rect 10644 -7902 10702 -7887
rect 10644 -7936 10656 -7902
rect 10690 -7936 10702 -7902
rect 10644 -7970 10702 -7936
rect 10644 -8004 10656 -7970
rect 10690 -8004 10702 -7970
rect 10644 -8038 10702 -8004
rect 10644 -8072 10656 -8038
rect 10690 -8072 10702 -8038
rect 10644 -8087 10702 -8072
rect 10902 -7902 10960 -7887
rect 10902 -7936 10914 -7902
rect 10948 -7936 10960 -7902
rect 10902 -7970 10960 -7936
rect 10902 -8004 10914 -7970
rect 10948 -8004 10960 -7970
rect 10902 -8038 10960 -8004
rect 10902 -8072 10914 -8038
rect 10948 -8072 10960 -8038
rect 10902 -8087 10960 -8072
rect 11160 -7902 11218 -7887
rect 11160 -7936 11172 -7902
rect 11206 -7936 11218 -7902
rect 11160 -7970 11218 -7936
rect 11160 -8004 11172 -7970
rect 11206 -8004 11218 -7970
rect 11160 -8038 11218 -8004
rect 11160 -8072 11172 -8038
rect 11206 -8072 11218 -8038
rect 11160 -8087 11218 -8072
rect 11354 -7902 11412 -7887
rect 11354 -7936 11366 -7902
rect 11400 -7936 11412 -7902
rect 11354 -7970 11412 -7936
rect 11354 -8004 11366 -7970
rect 11400 -8004 11412 -7970
rect 11354 -8038 11412 -8004
rect 11354 -8072 11366 -8038
rect 11400 -8072 11412 -8038
rect 11354 -8087 11412 -8072
rect 11612 -7902 11670 -7887
rect 11612 -7936 11624 -7902
rect 11658 -7936 11670 -7902
rect 11612 -7970 11670 -7936
rect 11612 -8004 11624 -7970
rect 11658 -8004 11670 -7970
rect 11612 -8038 11670 -8004
rect 11612 -8072 11624 -8038
rect 11658 -8072 11670 -8038
rect 11612 -8087 11670 -8072
rect 11870 -7902 11928 -7887
rect 11870 -7936 11882 -7902
rect 11916 -7936 11928 -7902
rect 11870 -7970 11928 -7936
rect 11870 -8004 11882 -7970
rect 11916 -8004 11928 -7970
rect 11870 -8038 11928 -8004
rect 11870 -8072 11882 -8038
rect 11916 -8072 11928 -8038
rect 11870 -8087 11928 -8072
rect 12128 -7902 12186 -7887
rect 12128 -7936 12140 -7902
rect 12174 -7936 12186 -7902
rect 12128 -7970 12186 -7936
rect 12128 -8004 12140 -7970
rect 12174 -8004 12186 -7970
rect 12128 -8038 12186 -8004
rect 12128 -8072 12140 -8038
rect 12174 -8072 12186 -8038
rect 12128 -8087 12186 -8072
rect 12322 -7902 12380 -7887
rect 12322 -7936 12334 -7902
rect 12368 -7936 12380 -7902
rect 12322 -7970 12380 -7936
rect 12322 -8004 12334 -7970
rect 12368 -8004 12380 -7970
rect 12322 -8038 12380 -8004
rect 12322 -8072 12334 -8038
rect 12368 -8072 12380 -8038
rect 12322 -8087 12380 -8072
rect 12580 -7902 12638 -7887
rect 12580 -7936 12592 -7902
rect 12626 -7936 12638 -7902
rect 12580 -7970 12638 -7936
rect 12580 -8004 12592 -7970
rect 12626 -8004 12638 -7970
rect 12580 -8038 12638 -8004
rect 12580 -8072 12592 -8038
rect 12626 -8072 12638 -8038
rect 12580 -8087 12638 -8072
rect 12838 -7902 12896 -7887
rect 12838 -7936 12850 -7902
rect 12884 -7936 12896 -7902
rect 12838 -7970 12896 -7936
rect 12838 -8004 12850 -7970
rect 12884 -8004 12896 -7970
rect 12838 -8038 12896 -8004
rect 12838 -8072 12850 -8038
rect 12884 -8072 12896 -8038
rect 12838 -8087 12896 -8072
rect 13096 -7902 13154 -7887
rect 13096 -7936 13108 -7902
rect 13142 -7936 13154 -7902
rect 13096 -7970 13154 -7936
rect 13096 -8004 13108 -7970
rect 13142 -8004 13154 -7970
rect 13096 -8038 13154 -8004
rect 13096 -8072 13108 -8038
rect 13142 -8072 13154 -8038
rect 13096 -8087 13154 -8072
rect 13354 -7902 13412 -7887
rect 13354 -7936 13366 -7902
rect 13400 -7936 13412 -7902
rect 13354 -7970 13412 -7936
rect 13354 -8004 13366 -7970
rect 13400 -8004 13412 -7970
rect 13354 -8038 13412 -8004
rect 13354 -8072 13366 -8038
rect 13400 -8072 13412 -8038
rect 13354 -8087 13412 -8072
rect 13548 -7902 13606 -7887
rect 13548 -7936 13560 -7902
rect 13594 -7936 13606 -7902
rect 13548 -7970 13606 -7936
rect 13548 -8004 13560 -7970
rect 13594 -8004 13606 -7970
rect 13548 -8038 13606 -8004
rect 13548 -8072 13560 -8038
rect 13594 -8072 13606 -8038
rect 13548 -8087 13606 -8072
rect 13806 -7902 13864 -7887
rect 13806 -7936 13818 -7902
rect 13852 -7936 13864 -7902
rect 13806 -7970 13864 -7936
rect 13806 -8004 13818 -7970
rect 13852 -8004 13864 -7970
rect 13806 -8038 13864 -8004
rect 13806 -8072 13818 -8038
rect 13852 -8072 13864 -8038
rect 13806 -8087 13864 -8072
rect 14034 -7902 14092 -7887
rect 14034 -7936 14046 -7902
rect 14080 -7936 14092 -7902
rect 14034 -7970 14092 -7936
rect 14034 -8004 14046 -7970
rect 14080 -8004 14092 -7970
rect 14034 -8038 14092 -8004
rect 14034 -8072 14046 -8038
rect 14080 -8072 14092 -8038
rect 14034 -8087 14092 -8072
rect 14292 -7902 14350 -7887
rect 14292 -7936 14304 -7902
rect 14338 -7936 14350 -7902
rect 14292 -7970 14350 -7936
rect 14292 -8004 14304 -7970
rect 14338 -8004 14350 -7970
rect 14292 -8038 14350 -8004
rect 14292 -8072 14304 -8038
rect 14338 -8072 14350 -8038
rect 14292 -8087 14350 -8072
rect 14485 -7902 14543 -7887
rect 14485 -7936 14497 -7902
rect 14531 -7936 14543 -7902
rect 14485 -7970 14543 -7936
rect 14485 -8004 14497 -7970
rect 14531 -8004 14543 -7970
rect 14485 -8038 14543 -8004
rect 14485 -8072 14497 -8038
rect 14531 -8072 14543 -8038
rect 14485 -8087 14543 -8072
rect 14743 -7902 14801 -7887
rect 14743 -7936 14755 -7902
rect 14789 -7936 14801 -7902
rect 14743 -7970 14801 -7936
rect 14743 -8004 14755 -7970
rect 14789 -8004 14801 -7970
rect 14743 -8038 14801 -8004
rect 14743 -8072 14755 -8038
rect 14789 -8072 14801 -8038
rect 14743 -8087 14801 -8072
rect 15001 -7902 15059 -7887
rect 15001 -7936 15013 -7902
rect 15047 -7936 15059 -7902
rect 15001 -7970 15059 -7936
rect 15001 -8004 15013 -7970
rect 15047 -8004 15059 -7970
rect 15001 -8038 15059 -8004
rect 15001 -8072 15013 -8038
rect 15047 -8072 15059 -8038
rect 15001 -8087 15059 -8072
rect 15259 -7902 15317 -7887
rect 15259 -7936 15271 -7902
rect 15305 -7936 15317 -7902
rect 15259 -7970 15317 -7936
rect 15259 -8004 15271 -7970
rect 15305 -8004 15317 -7970
rect 15259 -8038 15317 -8004
rect 15259 -8072 15271 -8038
rect 15305 -8072 15317 -8038
rect 15259 -8087 15317 -8072
rect 15517 -7902 15575 -7887
rect 15517 -7936 15529 -7902
rect 15563 -7936 15575 -7902
rect 15517 -7970 15575 -7936
rect 15517 -8004 15529 -7970
rect 15563 -8004 15575 -7970
rect 15517 -8038 15575 -8004
rect 15517 -8072 15529 -8038
rect 15563 -8072 15575 -8038
rect 15517 -8087 15575 -8072
rect 15711 -7902 15769 -7887
rect 15711 -7936 15723 -7902
rect 15757 -7936 15769 -7902
rect 15711 -7970 15769 -7936
rect 15711 -8004 15723 -7970
rect 15757 -8004 15769 -7970
rect 15711 -8038 15769 -8004
rect 15711 -8072 15723 -8038
rect 15757 -8072 15769 -8038
rect 15711 -8087 15769 -8072
rect 15969 -7902 16027 -7887
rect 15969 -7936 15981 -7902
rect 16015 -7936 16027 -7902
rect 15969 -7970 16027 -7936
rect 15969 -8004 15981 -7970
rect 16015 -8004 16027 -7970
rect 15969 -8038 16027 -8004
rect 15969 -8072 15981 -8038
rect 16015 -8072 16027 -8038
rect 15969 -8087 16027 -8072
rect 16227 -7902 16285 -7887
rect 16227 -7936 16239 -7902
rect 16273 -7936 16285 -7902
rect 16227 -7970 16285 -7936
rect 16227 -8004 16239 -7970
rect 16273 -8004 16285 -7970
rect 16227 -8038 16285 -8004
rect 16227 -8072 16239 -8038
rect 16273 -8072 16285 -8038
rect 16227 -8087 16285 -8072
rect 16485 -7902 16543 -7887
rect 16485 -7936 16497 -7902
rect 16531 -7936 16543 -7902
rect 16485 -7970 16543 -7936
rect 16485 -8004 16497 -7970
rect 16531 -8004 16543 -7970
rect 16485 -8038 16543 -8004
rect 16485 -8072 16497 -8038
rect 16531 -8072 16543 -8038
rect 16485 -8087 16543 -8072
rect 16679 -7902 16737 -7887
rect 16679 -7936 16691 -7902
rect 16725 -7936 16737 -7902
rect 16679 -7970 16737 -7936
rect 16679 -8004 16691 -7970
rect 16725 -8004 16737 -7970
rect 16679 -8038 16737 -8004
rect 16679 -8072 16691 -8038
rect 16725 -8072 16737 -8038
rect 16679 -8087 16737 -8072
rect 16937 -7902 16995 -7887
rect 16937 -7936 16949 -7902
rect 16983 -7936 16995 -7902
rect 16937 -7970 16995 -7936
rect 16937 -8004 16949 -7970
rect 16983 -8004 16995 -7970
rect 16937 -8038 16995 -8004
rect 16937 -8072 16949 -8038
rect 16983 -8072 16995 -8038
rect 16937 -8087 16995 -8072
rect 17195 -7902 17253 -7887
rect 17195 -7936 17207 -7902
rect 17241 -7936 17253 -7902
rect 17195 -7970 17253 -7936
rect 17195 -8004 17207 -7970
rect 17241 -8004 17253 -7970
rect 17195 -8038 17253 -8004
rect 17195 -8072 17207 -8038
rect 17241 -8072 17253 -8038
rect 17195 -8087 17253 -8072
rect 17453 -7902 17511 -7887
rect 17453 -7936 17465 -7902
rect 17499 -7936 17511 -7902
rect 17453 -7970 17511 -7936
rect 17453 -8004 17465 -7970
rect 17499 -8004 17511 -7970
rect 17453 -8038 17511 -8004
rect 17453 -8072 17465 -8038
rect 17499 -8072 17511 -8038
rect 17453 -8087 17511 -8072
rect 17711 -7902 17769 -7887
rect 17711 -7936 17723 -7902
rect 17757 -7936 17769 -7902
rect 17711 -7970 17769 -7936
rect 17711 -8004 17723 -7970
rect 17757 -8004 17769 -7970
rect 17711 -8038 17769 -8004
rect 17711 -8072 17723 -8038
rect 17757 -8072 17769 -8038
rect 17711 -8087 17769 -8072
rect 17905 -7902 17963 -7887
rect 17905 -7936 17917 -7902
rect 17951 -7936 17963 -7902
rect 17905 -7970 17963 -7936
rect 17905 -8004 17917 -7970
rect 17951 -8004 17963 -7970
rect 17905 -8038 17963 -8004
rect 17905 -8072 17917 -8038
rect 17951 -8072 17963 -8038
rect 17905 -8087 17963 -8072
rect 18163 -7902 18221 -7887
rect 18163 -7936 18175 -7902
rect 18209 -7936 18221 -7902
rect 18163 -7970 18221 -7936
rect 18163 -8004 18175 -7970
rect 18209 -8004 18221 -7970
rect 18163 -8038 18221 -8004
rect 18163 -8072 18175 -8038
rect 18209 -8072 18221 -8038
rect 18163 -8087 18221 -8072
rect 959 -8846 1017 -8831
rect 959 -8880 971 -8846
rect 1005 -8880 1017 -8846
rect 959 -8914 1017 -8880
rect 959 -8948 971 -8914
rect 1005 -8948 1017 -8914
rect 959 -8982 1017 -8948
rect 959 -9016 971 -8982
rect 1005 -9016 1017 -8982
rect 959 -9031 1017 -9016
rect 1217 -8846 1275 -8831
rect 1217 -8880 1229 -8846
rect 1263 -8880 1275 -8846
rect 1217 -8914 1275 -8880
rect 1217 -8948 1229 -8914
rect 1263 -8948 1275 -8914
rect 1217 -8982 1275 -8948
rect 1217 -9016 1229 -8982
rect 1263 -9016 1275 -8982
rect 1217 -9031 1275 -9016
rect 1411 -8846 1469 -8831
rect 1411 -8880 1423 -8846
rect 1457 -8880 1469 -8846
rect 1411 -8914 1469 -8880
rect 1411 -8948 1423 -8914
rect 1457 -8948 1469 -8914
rect 1411 -8982 1469 -8948
rect 1411 -9016 1423 -8982
rect 1457 -9016 1469 -8982
rect 1411 -9031 1469 -9016
rect 1669 -8846 1727 -8831
rect 1669 -8880 1681 -8846
rect 1715 -8880 1727 -8846
rect 1669 -8914 1727 -8880
rect 1669 -8948 1681 -8914
rect 1715 -8948 1727 -8914
rect 1669 -8982 1727 -8948
rect 1669 -9016 1681 -8982
rect 1715 -9016 1727 -8982
rect 1669 -9031 1727 -9016
rect 1927 -8846 1985 -8831
rect 1927 -8880 1939 -8846
rect 1973 -8880 1985 -8846
rect 1927 -8914 1985 -8880
rect 1927 -8948 1939 -8914
rect 1973 -8948 1985 -8914
rect 1927 -8982 1985 -8948
rect 1927 -9016 1939 -8982
rect 1973 -9016 1985 -8982
rect 1927 -9031 1985 -9016
rect 2185 -8846 2243 -8831
rect 2185 -8880 2197 -8846
rect 2231 -8880 2243 -8846
rect 2185 -8914 2243 -8880
rect 2185 -8948 2197 -8914
rect 2231 -8948 2243 -8914
rect 2185 -8982 2243 -8948
rect 2185 -9016 2197 -8982
rect 2231 -9016 2243 -8982
rect 2185 -9031 2243 -9016
rect 2443 -8846 2501 -8831
rect 2443 -8880 2455 -8846
rect 2489 -8880 2501 -8846
rect 2443 -8914 2501 -8880
rect 2443 -8948 2455 -8914
rect 2489 -8948 2501 -8914
rect 2443 -8982 2501 -8948
rect 2443 -9016 2455 -8982
rect 2489 -9016 2501 -8982
rect 2443 -9031 2501 -9016
rect 2637 -8846 2695 -8831
rect 2637 -8880 2649 -8846
rect 2683 -8880 2695 -8846
rect 2637 -8914 2695 -8880
rect 2637 -8948 2649 -8914
rect 2683 -8948 2695 -8914
rect 2637 -8982 2695 -8948
rect 2637 -9016 2649 -8982
rect 2683 -9016 2695 -8982
rect 2637 -9031 2695 -9016
rect 2895 -8846 2953 -8831
rect 2895 -8880 2907 -8846
rect 2941 -8880 2953 -8846
rect 2895 -8914 2953 -8880
rect 2895 -8948 2907 -8914
rect 2941 -8948 2953 -8914
rect 2895 -8982 2953 -8948
rect 2895 -9016 2907 -8982
rect 2941 -9016 2953 -8982
rect 2895 -9031 2953 -9016
rect 3153 -8846 3211 -8831
rect 3153 -8880 3165 -8846
rect 3199 -8880 3211 -8846
rect 3153 -8914 3211 -8880
rect 3153 -8948 3165 -8914
rect 3199 -8948 3211 -8914
rect 3153 -8982 3211 -8948
rect 3153 -9016 3165 -8982
rect 3199 -9016 3211 -8982
rect 3153 -9031 3211 -9016
rect 3411 -8846 3469 -8831
rect 3411 -8880 3423 -8846
rect 3457 -8880 3469 -8846
rect 3411 -8914 3469 -8880
rect 3411 -8948 3423 -8914
rect 3457 -8948 3469 -8914
rect 3411 -8982 3469 -8948
rect 3411 -9016 3423 -8982
rect 3457 -9016 3469 -8982
rect 3411 -9031 3469 -9016
rect 3605 -8846 3663 -8831
rect 3605 -8880 3617 -8846
rect 3651 -8880 3663 -8846
rect 3605 -8914 3663 -8880
rect 3605 -8948 3617 -8914
rect 3651 -8948 3663 -8914
rect 3605 -8982 3663 -8948
rect 3605 -9016 3617 -8982
rect 3651 -9016 3663 -8982
rect 3605 -9031 3663 -9016
rect 3863 -8846 3921 -8831
rect 3863 -8880 3875 -8846
rect 3909 -8880 3921 -8846
rect 3863 -8914 3921 -8880
rect 3863 -8948 3875 -8914
rect 3909 -8948 3921 -8914
rect 3863 -8982 3921 -8948
rect 3863 -9016 3875 -8982
rect 3909 -9016 3921 -8982
rect 3863 -9031 3921 -9016
rect 4121 -8846 4179 -8831
rect 4121 -8880 4133 -8846
rect 4167 -8880 4179 -8846
rect 4121 -8914 4179 -8880
rect 4121 -8948 4133 -8914
rect 4167 -8948 4179 -8914
rect 4121 -8982 4179 -8948
rect 4121 -9016 4133 -8982
rect 4167 -9016 4179 -8982
rect 4121 -9031 4179 -9016
rect 4379 -8846 4437 -8831
rect 4379 -8880 4391 -8846
rect 4425 -8880 4437 -8846
rect 4379 -8914 4437 -8880
rect 4379 -8948 4391 -8914
rect 4425 -8948 4437 -8914
rect 4379 -8982 4437 -8948
rect 4379 -9016 4391 -8982
rect 4425 -9016 4437 -8982
rect 4379 -9031 4437 -9016
rect 4637 -8846 4695 -8831
rect 4637 -8880 4649 -8846
rect 4683 -8880 4695 -8846
rect 4637 -8914 4695 -8880
rect 4637 -8948 4649 -8914
rect 4683 -8948 4695 -8914
rect 4637 -8982 4695 -8948
rect 4637 -9016 4649 -8982
rect 4683 -9016 4695 -8982
rect 4637 -9031 4695 -9016
rect 4830 -8846 4888 -8831
rect 4830 -8880 4842 -8846
rect 4876 -8880 4888 -8846
rect 4830 -8914 4888 -8880
rect 4830 -8948 4842 -8914
rect 4876 -8948 4888 -8914
rect 4830 -8982 4888 -8948
rect 4830 -9016 4842 -8982
rect 4876 -9016 4888 -8982
rect 4830 -9031 4888 -9016
rect 5088 -8846 5146 -8831
rect 5088 -8880 5100 -8846
rect 5134 -8880 5146 -8846
rect 5088 -8914 5146 -8880
rect 5088 -8948 5100 -8914
rect 5134 -8948 5146 -8914
rect 5088 -8982 5146 -8948
rect 5088 -9016 5100 -8982
rect 5134 -9016 5146 -8982
rect 5088 -9031 5146 -9016
rect 5316 -8846 5374 -8831
rect 5316 -8880 5328 -8846
rect 5362 -8880 5374 -8846
rect 5316 -8914 5374 -8880
rect 5316 -8948 5328 -8914
rect 5362 -8948 5374 -8914
rect 5316 -8982 5374 -8948
rect 5316 -9016 5328 -8982
rect 5362 -9016 5374 -8982
rect 5316 -9031 5374 -9016
rect 5574 -8846 5632 -8831
rect 5574 -8880 5586 -8846
rect 5620 -8880 5632 -8846
rect 5574 -8914 5632 -8880
rect 5574 -8948 5586 -8914
rect 5620 -8948 5632 -8914
rect 5574 -8982 5632 -8948
rect 5574 -9016 5586 -8982
rect 5620 -9016 5632 -8982
rect 5574 -9031 5632 -9016
rect 5768 -8846 5826 -8831
rect 5768 -8880 5780 -8846
rect 5814 -8880 5826 -8846
rect 5768 -8914 5826 -8880
rect 5768 -8948 5780 -8914
rect 5814 -8948 5826 -8914
rect 5768 -8982 5826 -8948
rect 5768 -9016 5780 -8982
rect 5814 -9016 5826 -8982
rect 5768 -9031 5826 -9016
rect 6026 -8846 6084 -8831
rect 6026 -8880 6038 -8846
rect 6072 -8880 6084 -8846
rect 6026 -8914 6084 -8880
rect 6026 -8948 6038 -8914
rect 6072 -8948 6084 -8914
rect 6026 -8982 6084 -8948
rect 6026 -9016 6038 -8982
rect 6072 -9016 6084 -8982
rect 6026 -9031 6084 -9016
rect 6284 -8846 6342 -8831
rect 6284 -8880 6296 -8846
rect 6330 -8880 6342 -8846
rect 6284 -8914 6342 -8880
rect 6284 -8948 6296 -8914
rect 6330 -8948 6342 -8914
rect 6284 -8982 6342 -8948
rect 6284 -9016 6296 -8982
rect 6330 -9016 6342 -8982
rect 6284 -9031 6342 -9016
rect 6542 -8846 6600 -8831
rect 6542 -8880 6554 -8846
rect 6588 -8880 6600 -8846
rect 6542 -8914 6600 -8880
rect 6542 -8948 6554 -8914
rect 6588 -8948 6600 -8914
rect 6542 -8982 6600 -8948
rect 6542 -9016 6554 -8982
rect 6588 -9016 6600 -8982
rect 6542 -9031 6600 -9016
rect 6800 -8846 6858 -8831
rect 6800 -8880 6812 -8846
rect 6846 -8880 6858 -8846
rect 6800 -8914 6858 -8880
rect 6800 -8948 6812 -8914
rect 6846 -8948 6858 -8914
rect 6800 -8982 6858 -8948
rect 6800 -9016 6812 -8982
rect 6846 -9016 6858 -8982
rect 6800 -9031 6858 -9016
rect 6994 -8846 7052 -8831
rect 6994 -8880 7006 -8846
rect 7040 -8880 7052 -8846
rect 6994 -8914 7052 -8880
rect 6994 -8948 7006 -8914
rect 7040 -8948 7052 -8914
rect 6994 -8982 7052 -8948
rect 6994 -9016 7006 -8982
rect 7040 -9016 7052 -8982
rect 6994 -9031 7052 -9016
rect 7252 -8846 7310 -8831
rect 7252 -8880 7264 -8846
rect 7298 -8880 7310 -8846
rect 7252 -8914 7310 -8880
rect 7252 -8948 7264 -8914
rect 7298 -8948 7310 -8914
rect 7252 -8982 7310 -8948
rect 7252 -9016 7264 -8982
rect 7298 -9016 7310 -8982
rect 7252 -9031 7310 -9016
rect 7510 -8846 7568 -8831
rect 7510 -8880 7522 -8846
rect 7556 -8880 7568 -8846
rect 7510 -8914 7568 -8880
rect 7510 -8948 7522 -8914
rect 7556 -8948 7568 -8914
rect 7510 -8982 7568 -8948
rect 7510 -9016 7522 -8982
rect 7556 -9016 7568 -8982
rect 7510 -9031 7568 -9016
rect 7768 -8846 7826 -8831
rect 7768 -8880 7780 -8846
rect 7814 -8880 7826 -8846
rect 7768 -8914 7826 -8880
rect 7768 -8948 7780 -8914
rect 7814 -8948 7826 -8914
rect 7768 -8982 7826 -8948
rect 7768 -9016 7780 -8982
rect 7814 -9016 7826 -8982
rect 7768 -9031 7826 -9016
rect 7962 -8846 8020 -8831
rect 7962 -8880 7974 -8846
rect 8008 -8880 8020 -8846
rect 7962 -8914 8020 -8880
rect 7962 -8948 7974 -8914
rect 8008 -8948 8020 -8914
rect 7962 -8982 8020 -8948
rect 7962 -9016 7974 -8982
rect 8008 -9016 8020 -8982
rect 7962 -9031 8020 -9016
rect 8220 -8846 8278 -8831
rect 8220 -8880 8232 -8846
rect 8266 -8880 8278 -8846
rect 8220 -8914 8278 -8880
rect 8220 -8948 8232 -8914
rect 8266 -8948 8278 -8914
rect 8220 -8982 8278 -8948
rect 8220 -9016 8232 -8982
rect 8266 -9016 8278 -8982
rect 8220 -9031 8278 -9016
rect 8478 -8846 8536 -8831
rect 8478 -8880 8490 -8846
rect 8524 -8880 8536 -8846
rect 8478 -8914 8536 -8880
rect 8478 -8948 8490 -8914
rect 8524 -8948 8536 -8914
rect 8478 -8982 8536 -8948
rect 8478 -9016 8490 -8982
rect 8524 -9016 8536 -8982
rect 8478 -9031 8536 -9016
rect 8736 -8846 8794 -8831
rect 8736 -8880 8748 -8846
rect 8782 -8880 8794 -8846
rect 8736 -8914 8794 -8880
rect 8736 -8948 8748 -8914
rect 8782 -8948 8794 -8914
rect 8736 -8982 8794 -8948
rect 8736 -9016 8748 -8982
rect 8782 -9016 8794 -8982
rect 8736 -9031 8794 -9016
rect 8994 -8846 9052 -8831
rect 8994 -8880 9006 -8846
rect 9040 -8880 9052 -8846
rect 8994 -8914 9052 -8880
rect 8994 -8948 9006 -8914
rect 9040 -8948 9052 -8914
rect 8994 -8982 9052 -8948
rect 8994 -9016 9006 -8982
rect 9040 -9016 9052 -8982
rect 8994 -9031 9052 -9016
rect 9188 -8846 9246 -8831
rect 9188 -8880 9200 -8846
rect 9234 -8880 9246 -8846
rect 9188 -8914 9246 -8880
rect 9188 -8948 9200 -8914
rect 9234 -8948 9246 -8914
rect 9188 -8982 9246 -8948
rect 9188 -9016 9200 -8982
rect 9234 -9016 9246 -8982
rect 9188 -9031 9246 -9016
rect 9446 -8846 9504 -8831
rect 9446 -8880 9458 -8846
rect 9492 -8880 9504 -8846
rect 9446 -8914 9504 -8880
rect 9446 -8948 9458 -8914
rect 9492 -8948 9504 -8914
rect 9446 -8982 9504 -8948
rect 9446 -9016 9458 -8982
rect 9492 -9016 9504 -8982
rect 9446 -9031 9504 -9016
rect 9676 -8846 9734 -8831
rect 9676 -8880 9688 -8846
rect 9722 -8880 9734 -8846
rect 9676 -8914 9734 -8880
rect 9676 -8948 9688 -8914
rect 9722 -8948 9734 -8914
rect 9676 -8982 9734 -8948
rect 9676 -9016 9688 -8982
rect 9722 -9016 9734 -8982
rect 9676 -9031 9734 -9016
rect 9934 -8846 9992 -8831
rect 9934 -8880 9946 -8846
rect 9980 -8880 9992 -8846
rect 9934 -8914 9992 -8880
rect 9934 -8948 9946 -8914
rect 9980 -8948 9992 -8914
rect 9934 -8982 9992 -8948
rect 9934 -9016 9946 -8982
rect 9980 -9016 9992 -8982
rect 9934 -9031 9992 -9016
rect 10128 -8846 10186 -8831
rect 10128 -8880 10140 -8846
rect 10174 -8880 10186 -8846
rect 10128 -8914 10186 -8880
rect 10128 -8948 10140 -8914
rect 10174 -8948 10186 -8914
rect 10128 -8982 10186 -8948
rect 10128 -9016 10140 -8982
rect 10174 -9016 10186 -8982
rect 10128 -9031 10186 -9016
rect 10386 -8846 10444 -8831
rect 10386 -8880 10398 -8846
rect 10432 -8880 10444 -8846
rect 10386 -8914 10444 -8880
rect 10386 -8948 10398 -8914
rect 10432 -8948 10444 -8914
rect 10386 -8982 10444 -8948
rect 10386 -9016 10398 -8982
rect 10432 -9016 10444 -8982
rect 10386 -9031 10444 -9016
rect 10644 -8846 10702 -8831
rect 10644 -8880 10656 -8846
rect 10690 -8880 10702 -8846
rect 10644 -8914 10702 -8880
rect 10644 -8948 10656 -8914
rect 10690 -8948 10702 -8914
rect 10644 -8982 10702 -8948
rect 10644 -9016 10656 -8982
rect 10690 -9016 10702 -8982
rect 10644 -9031 10702 -9016
rect 10902 -8846 10960 -8831
rect 10902 -8880 10914 -8846
rect 10948 -8880 10960 -8846
rect 10902 -8914 10960 -8880
rect 10902 -8948 10914 -8914
rect 10948 -8948 10960 -8914
rect 10902 -8982 10960 -8948
rect 10902 -9016 10914 -8982
rect 10948 -9016 10960 -8982
rect 10902 -9031 10960 -9016
rect 11160 -8846 11218 -8831
rect 11160 -8880 11172 -8846
rect 11206 -8880 11218 -8846
rect 11160 -8914 11218 -8880
rect 11160 -8948 11172 -8914
rect 11206 -8948 11218 -8914
rect 11160 -8982 11218 -8948
rect 11160 -9016 11172 -8982
rect 11206 -9016 11218 -8982
rect 11160 -9031 11218 -9016
rect 11354 -8846 11412 -8831
rect 11354 -8880 11366 -8846
rect 11400 -8880 11412 -8846
rect 11354 -8914 11412 -8880
rect 11354 -8948 11366 -8914
rect 11400 -8948 11412 -8914
rect 11354 -8982 11412 -8948
rect 11354 -9016 11366 -8982
rect 11400 -9016 11412 -8982
rect 11354 -9031 11412 -9016
rect 11612 -8846 11670 -8831
rect 11612 -8880 11624 -8846
rect 11658 -8880 11670 -8846
rect 11612 -8914 11670 -8880
rect 11612 -8948 11624 -8914
rect 11658 -8948 11670 -8914
rect 11612 -8982 11670 -8948
rect 11612 -9016 11624 -8982
rect 11658 -9016 11670 -8982
rect 11612 -9031 11670 -9016
rect 11870 -8846 11928 -8831
rect 11870 -8880 11882 -8846
rect 11916 -8880 11928 -8846
rect 11870 -8914 11928 -8880
rect 11870 -8948 11882 -8914
rect 11916 -8948 11928 -8914
rect 11870 -8982 11928 -8948
rect 11870 -9016 11882 -8982
rect 11916 -9016 11928 -8982
rect 11870 -9031 11928 -9016
rect 12128 -8846 12186 -8831
rect 12128 -8880 12140 -8846
rect 12174 -8880 12186 -8846
rect 12128 -8914 12186 -8880
rect 12128 -8948 12140 -8914
rect 12174 -8948 12186 -8914
rect 12128 -8982 12186 -8948
rect 12128 -9016 12140 -8982
rect 12174 -9016 12186 -8982
rect 12128 -9031 12186 -9016
rect 12322 -8846 12380 -8831
rect 12322 -8880 12334 -8846
rect 12368 -8880 12380 -8846
rect 12322 -8914 12380 -8880
rect 12322 -8948 12334 -8914
rect 12368 -8948 12380 -8914
rect 12322 -8982 12380 -8948
rect 12322 -9016 12334 -8982
rect 12368 -9016 12380 -8982
rect 12322 -9031 12380 -9016
rect 12580 -8846 12638 -8831
rect 12580 -8880 12592 -8846
rect 12626 -8880 12638 -8846
rect 12580 -8914 12638 -8880
rect 12580 -8948 12592 -8914
rect 12626 -8948 12638 -8914
rect 12580 -8982 12638 -8948
rect 12580 -9016 12592 -8982
rect 12626 -9016 12638 -8982
rect 12580 -9031 12638 -9016
rect 12838 -8846 12896 -8831
rect 12838 -8880 12850 -8846
rect 12884 -8880 12896 -8846
rect 12838 -8914 12896 -8880
rect 12838 -8948 12850 -8914
rect 12884 -8948 12896 -8914
rect 12838 -8982 12896 -8948
rect 12838 -9016 12850 -8982
rect 12884 -9016 12896 -8982
rect 12838 -9031 12896 -9016
rect 13096 -8846 13154 -8831
rect 13096 -8880 13108 -8846
rect 13142 -8880 13154 -8846
rect 13096 -8914 13154 -8880
rect 13096 -8948 13108 -8914
rect 13142 -8948 13154 -8914
rect 13096 -8982 13154 -8948
rect 13096 -9016 13108 -8982
rect 13142 -9016 13154 -8982
rect 13096 -9031 13154 -9016
rect 13354 -8846 13412 -8831
rect 13354 -8880 13366 -8846
rect 13400 -8880 13412 -8846
rect 13354 -8914 13412 -8880
rect 13354 -8948 13366 -8914
rect 13400 -8948 13412 -8914
rect 13354 -8982 13412 -8948
rect 13354 -9016 13366 -8982
rect 13400 -9016 13412 -8982
rect 13354 -9031 13412 -9016
rect 13548 -8846 13606 -8831
rect 13548 -8880 13560 -8846
rect 13594 -8880 13606 -8846
rect 13548 -8914 13606 -8880
rect 13548 -8948 13560 -8914
rect 13594 -8948 13606 -8914
rect 13548 -8982 13606 -8948
rect 13548 -9016 13560 -8982
rect 13594 -9016 13606 -8982
rect 13548 -9031 13606 -9016
rect 13806 -8846 13864 -8831
rect 13806 -8880 13818 -8846
rect 13852 -8880 13864 -8846
rect 13806 -8914 13864 -8880
rect 13806 -8948 13818 -8914
rect 13852 -8948 13864 -8914
rect 13806 -8982 13864 -8948
rect 13806 -9016 13818 -8982
rect 13852 -9016 13864 -8982
rect 13806 -9031 13864 -9016
rect 14034 -8846 14092 -8831
rect 14034 -8880 14046 -8846
rect 14080 -8880 14092 -8846
rect 14034 -8914 14092 -8880
rect 14034 -8948 14046 -8914
rect 14080 -8948 14092 -8914
rect 14034 -8982 14092 -8948
rect 14034 -9016 14046 -8982
rect 14080 -9016 14092 -8982
rect 14034 -9031 14092 -9016
rect 14292 -8846 14350 -8831
rect 14292 -8880 14304 -8846
rect 14338 -8880 14350 -8846
rect 14292 -8914 14350 -8880
rect 14292 -8948 14304 -8914
rect 14338 -8948 14350 -8914
rect 14292 -8982 14350 -8948
rect 14292 -9016 14304 -8982
rect 14338 -9016 14350 -8982
rect 14292 -9031 14350 -9016
rect 14485 -8846 14543 -8831
rect 14485 -8880 14497 -8846
rect 14531 -8880 14543 -8846
rect 14485 -8914 14543 -8880
rect 14485 -8948 14497 -8914
rect 14531 -8948 14543 -8914
rect 14485 -8982 14543 -8948
rect 14485 -9016 14497 -8982
rect 14531 -9016 14543 -8982
rect 14485 -9031 14543 -9016
rect 14743 -8846 14801 -8831
rect 14743 -8880 14755 -8846
rect 14789 -8880 14801 -8846
rect 14743 -8914 14801 -8880
rect 14743 -8948 14755 -8914
rect 14789 -8948 14801 -8914
rect 14743 -8982 14801 -8948
rect 14743 -9016 14755 -8982
rect 14789 -9016 14801 -8982
rect 14743 -9031 14801 -9016
rect 15001 -8846 15059 -8831
rect 15001 -8880 15013 -8846
rect 15047 -8880 15059 -8846
rect 15001 -8914 15059 -8880
rect 15001 -8948 15013 -8914
rect 15047 -8948 15059 -8914
rect 15001 -8982 15059 -8948
rect 15001 -9016 15013 -8982
rect 15047 -9016 15059 -8982
rect 15001 -9031 15059 -9016
rect 15259 -8846 15317 -8831
rect 15259 -8880 15271 -8846
rect 15305 -8880 15317 -8846
rect 15259 -8914 15317 -8880
rect 15259 -8948 15271 -8914
rect 15305 -8948 15317 -8914
rect 15259 -8982 15317 -8948
rect 15259 -9016 15271 -8982
rect 15305 -9016 15317 -8982
rect 15259 -9031 15317 -9016
rect 15517 -8846 15575 -8831
rect 15517 -8880 15529 -8846
rect 15563 -8880 15575 -8846
rect 15517 -8914 15575 -8880
rect 15517 -8948 15529 -8914
rect 15563 -8948 15575 -8914
rect 15517 -8982 15575 -8948
rect 15517 -9016 15529 -8982
rect 15563 -9016 15575 -8982
rect 15517 -9031 15575 -9016
rect 15711 -8846 15769 -8831
rect 15711 -8880 15723 -8846
rect 15757 -8880 15769 -8846
rect 15711 -8914 15769 -8880
rect 15711 -8948 15723 -8914
rect 15757 -8948 15769 -8914
rect 15711 -8982 15769 -8948
rect 15711 -9016 15723 -8982
rect 15757 -9016 15769 -8982
rect 15711 -9031 15769 -9016
rect 15969 -8846 16027 -8831
rect 15969 -8880 15981 -8846
rect 16015 -8880 16027 -8846
rect 15969 -8914 16027 -8880
rect 15969 -8948 15981 -8914
rect 16015 -8948 16027 -8914
rect 15969 -8982 16027 -8948
rect 15969 -9016 15981 -8982
rect 16015 -9016 16027 -8982
rect 15969 -9031 16027 -9016
rect 16227 -8846 16285 -8831
rect 16227 -8880 16239 -8846
rect 16273 -8880 16285 -8846
rect 16227 -8914 16285 -8880
rect 16227 -8948 16239 -8914
rect 16273 -8948 16285 -8914
rect 16227 -8982 16285 -8948
rect 16227 -9016 16239 -8982
rect 16273 -9016 16285 -8982
rect 16227 -9031 16285 -9016
rect 16485 -8846 16543 -8831
rect 16485 -8880 16497 -8846
rect 16531 -8880 16543 -8846
rect 16485 -8914 16543 -8880
rect 16485 -8948 16497 -8914
rect 16531 -8948 16543 -8914
rect 16485 -8982 16543 -8948
rect 16485 -9016 16497 -8982
rect 16531 -9016 16543 -8982
rect 16485 -9031 16543 -9016
rect 16679 -8846 16737 -8831
rect 16679 -8880 16691 -8846
rect 16725 -8880 16737 -8846
rect 16679 -8914 16737 -8880
rect 16679 -8948 16691 -8914
rect 16725 -8948 16737 -8914
rect 16679 -8982 16737 -8948
rect 16679 -9016 16691 -8982
rect 16725 -9016 16737 -8982
rect 16679 -9031 16737 -9016
rect 16937 -8846 16995 -8831
rect 16937 -8880 16949 -8846
rect 16983 -8880 16995 -8846
rect 16937 -8914 16995 -8880
rect 16937 -8948 16949 -8914
rect 16983 -8948 16995 -8914
rect 16937 -8982 16995 -8948
rect 16937 -9016 16949 -8982
rect 16983 -9016 16995 -8982
rect 16937 -9031 16995 -9016
rect 17195 -8846 17253 -8831
rect 17195 -8880 17207 -8846
rect 17241 -8880 17253 -8846
rect 17195 -8914 17253 -8880
rect 17195 -8948 17207 -8914
rect 17241 -8948 17253 -8914
rect 17195 -8982 17253 -8948
rect 17195 -9016 17207 -8982
rect 17241 -9016 17253 -8982
rect 17195 -9031 17253 -9016
rect 17453 -8846 17511 -8831
rect 17453 -8880 17465 -8846
rect 17499 -8880 17511 -8846
rect 17453 -8914 17511 -8880
rect 17453 -8948 17465 -8914
rect 17499 -8948 17511 -8914
rect 17453 -8982 17511 -8948
rect 17453 -9016 17465 -8982
rect 17499 -9016 17511 -8982
rect 17453 -9031 17511 -9016
rect 17711 -8846 17769 -8831
rect 17711 -8880 17723 -8846
rect 17757 -8880 17769 -8846
rect 17711 -8914 17769 -8880
rect 17711 -8948 17723 -8914
rect 17757 -8948 17769 -8914
rect 17711 -8982 17769 -8948
rect 17711 -9016 17723 -8982
rect 17757 -9016 17769 -8982
rect 17711 -9031 17769 -9016
rect 17905 -8846 17963 -8831
rect 17905 -8880 17917 -8846
rect 17951 -8880 17963 -8846
rect 17905 -8914 17963 -8880
rect 17905 -8948 17917 -8914
rect 17951 -8948 17963 -8914
rect 17905 -8982 17963 -8948
rect 17905 -9016 17917 -8982
rect 17951 -9016 17963 -8982
rect 17905 -9031 17963 -9016
rect 18163 -8846 18221 -8831
rect 18163 -8880 18175 -8846
rect 18209 -8880 18221 -8846
rect 18163 -8914 18221 -8880
rect 18163 -8948 18175 -8914
rect 18209 -8948 18221 -8914
rect 18163 -8982 18221 -8948
rect 18163 -9016 18175 -8982
rect 18209 -9016 18221 -8982
rect 18163 -9031 18221 -9016
<< pdiffc >>
rect 971 219 1005 253
rect 971 151 1005 185
rect 971 83 1005 117
rect 1229 219 1263 253
rect 1229 151 1263 185
rect 1229 83 1263 117
rect 1423 219 1457 253
rect 1423 151 1457 185
rect 1423 83 1457 117
rect 1681 219 1715 253
rect 1681 151 1715 185
rect 1681 83 1715 117
rect 1939 219 1973 253
rect 1939 151 1973 185
rect 1939 83 1973 117
rect 2197 219 2231 253
rect 2197 151 2231 185
rect 2197 83 2231 117
rect 2455 219 2489 253
rect 2455 151 2489 185
rect 2455 83 2489 117
rect 2649 219 2683 253
rect 2649 151 2683 185
rect 2649 83 2683 117
rect 2907 219 2941 253
rect 2907 151 2941 185
rect 2907 83 2941 117
rect 3165 219 3199 253
rect 3165 151 3199 185
rect 3165 83 3199 117
rect 3423 219 3457 253
rect 3423 151 3457 185
rect 3423 83 3457 117
rect 3617 219 3651 253
rect 3617 151 3651 185
rect 3617 83 3651 117
rect 3875 219 3909 253
rect 3875 151 3909 185
rect 3875 83 3909 117
rect 4133 219 4167 253
rect 4133 151 4167 185
rect 4133 83 4167 117
rect 4391 219 4425 253
rect 4391 151 4425 185
rect 4391 83 4425 117
rect 4649 219 4683 253
rect 4649 151 4683 185
rect 4649 83 4683 117
rect 4842 219 4876 253
rect 4842 151 4876 185
rect 4842 83 4876 117
rect 5100 219 5134 253
rect 5100 151 5134 185
rect 5100 83 5134 117
rect 5328 219 5362 253
rect 5328 151 5362 185
rect 5328 83 5362 117
rect 5586 219 5620 253
rect 5586 151 5620 185
rect 5586 83 5620 117
rect 5780 219 5814 253
rect 5780 151 5814 185
rect 5780 83 5814 117
rect 6038 219 6072 253
rect 6038 151 6072 185
rect 6038 83 6072 117
rect 6296 219 6330 253
rect 6296 151 6330 185
rect 6296 83 6330 117
rect 6554 219 6588 253
rect 6554 151 6588 185
rect 6554 83 6588 117
rect 6812 219 6846 253
rect 6812 151 6846 185
rect 6812 83 6846 117
rect 7006 219 7040 253
rect 7006 151 7040 185
rect 7006 83 7040 117
rect 7264 219 7298 253
rect 7264 151 7298 185
rect 7264 83 7298 117
rect 7522 219 7556 253
rect 7522 151 7556 185
rect 7522 83 7556 117
rect 7780 219 7814 253
rect 7780 151 7814 185
rect 7780 83 7814 117
rect 7974 219 8008 253
rect 7974 151 8008 185
rect 7974 83 8008 117
rect 8232 219 8266 253
rect 8232 151 8266 185
rect 8232 83 8266 117
rect 8490 219 8524 253
rect 8490 151 8524 185
rect 8490 83 8524 117
rect 8748 219 8782 253
rect 8748 151 8782 185
rect 8748 83 8782 117
rect 9006 219 9040 253
rect 9006 151 9040 185
rect 9006 83 9040 117
rect 9200 219 9234 253
rect 9200 151 9234 185
rect 9200 83 9234 117
rect 9458 219 9492 253
rect 9458 151 9492 185
rect 9458 83 9492 117
rect 9688 219 9722 253
rect 9688 151 9722 185
rect 9688 83 9722 117
rect 9946 219 9980 253
rect 9946 151 9980 185
rect 9946 83 9980 117
rect 10140 219 10174 253
rect 10140 151 10174 185
rect 10140 83 10174 117
rect 10398 219 10432 253
rect 10398 151 10432 185
rect 10398 83 10432 117
rect 10656 219 10690 253
rect 10656 151 10690 185
rect 10656 83 10690 117
rect 10914 219 10948 253
rect 10914 151 10948 185
rect 10914 83 10948 117
rect 11172 219 11206 253
rect 11172 151 11206 185
rect 11172 83 11206 117
rect 11366 219 11400 253
rect 11366 151 11400 185
rect 11366 83 11400 117
rect 11624 219 11658 253
rect 11624 151 11658 185
rect 11624 83 11658 117
rect 11882 219 11916 253
rect 11882 151 11916 185
rect 11882 83 11916 117
rect 12140 219 12174 253
rect 12140 151 12174 185
rect 12140 83 12174 117
rect 12334 219 12368 253
rect 12334 151 12368 185
rect 12334 83 12368 117
rect 12592 219 12626 253
rect 12592 151 12626 185
rect 12592 83 12626 117
rect 12850 219 12884 253
rect 12850 151 12884 185
rect 12850 83 12884 117
rect 13108 219 13142 253
rect 13108 151 13142 185
rect 13108 83 13142 117
rect 13366 219 13400 253
rect 13366 151 13400 185
rect 13366 83 13400 117
rect 13560 219 13594 253
rect 13560 151 13594 185
rect 13560 83 13594 117
rect 13818 219 13852 253
rect 13818 151 13852 185
rect 13818 83 13852 117
rect 14046 219 14080 253
rect 14046 151 14080 185
rect 14046 83 14080 117
rect 14304 219 14338 253
rect 14304 151 14338 185
rect 14304 83 14338 117
rect 14497 219 14531 253
rect 14497 151 14531 185
rect 14497 83 14531 117
rect 14755 219 14789 253
rect 14755 151 14789 185
rect 14755 83 14789 117
rect 15013 219 15047 253
rect 15013 151 15047 185
rect 15013 83 15047 117
rect 15271 219 15305 253
rect 15271 151 15305 185
rect 15271 83 15305 117
rect 15529 219 15563 253
rect 15529 151 15563 185
rect 15529 83 15563 117
rect 15723 219 15757 253
rect 15723 151 15757 185
rect 15723 83 15757 117
rect 15981 219 16015 253
rect 15981 151 16015 185
rect 15981 83 16015 117
rect 16239 219 16273 253
rect 16239 151 16273 185
rect 16239 83 16273 117
rect 16497 219 16531 253
rect 16497 151 16531 185
rect 16497 83 16531 117
rect 16691 219 16725 253
rect 16691 151 16725 185
rect 16691 83 16725 117
rect 16949 219 16983 253
rect 16949 151 16983 185
rect 16949 83 16983 117
rect 17207 219 17241 253
rect 17207 151 17241 185
rect 17207 83 17241 117
rect 17465 219 17499 253
rect 17465 151 17499 185
rect 17465 83 17499 117
rect 17723 219 17757 253
rect 17723 151 17757 185
rect 17723 83 17757 117
rect 17917 219 17951 253
rect 17917 151 17951 185
rect 17917 83 17951 117
rect 18175 219 18209 253
rect 18175 151 18209 185
rect 18175 83 18209 117
rect 971 -725 1005 -691
rect 971 -793 1005 -759
rect 971 -861 1005 -827
rect 1229 -725 1263 -691
rect 1229 -793 1263 -759
rect 1229 -861 1263 -827
rect 1423 -725 1457 -691
rect 1423 -793 1457 -759
rect 1423 -861 1457 -827
rect 1681 -725 1715 -691
rect 1681 -793 1715 -759
rect 1681 -861 1715 -827
rect 1939 -725 1973 -691
rect 1939 -793 1973 -759
rect 1939 -861 1973 -827
rect 2197 -725 2231 -691
rect 2197 -793 2231 -759
rect 2197 -861 2231 -827
rect 2455 -725 2489 -691
rect 2455 -793 2489 -759
rect 2455 -861 2489 -827
rect 2649 -725 2683 -691
rect 2649 -793 2683 -759
rect 2649 -861 2683 -827
rect 2907 -725 2941 -691
rect 2907 -793 2941 -759
rect 2907 -861 2941 -827
rect 3165 -725 3199 -691
rect 3165 -793 3199 -759
rect 3165 -861 3199 -827
rect 3423 -725 3457 -691
rect 3423 -793 3457 -759
rect 3423 -861 3457 -827
rect 3617 -725 3651 -691
rect 3617 -793 3651 -759
rect 3617 -861 3651 -827
rect 3875 -725 3909 -691
rect 3875 -793 3909 -759
rect 3875 -861 3909 -827
rect 4133 -725 4167 -691
rect 4133 -793 4167 -759
rect 4133 -861 4167 -827
rect 4391 -725 4425 -691
rect 4391 -793 4425 -759
rect 4391 -861 4425 -827
rect 4649 -725 4683 -691
rect 4649 -793 4683 -759
rect 4649 -861 4683 -827
rect 4842 -725 4876 -691
rect 4842 -793 4876 -759
rect 4842 -861 4876 -827
rect 5100 -725 5134 -691
rect 5100 -793 5134 -759
rect 5100 -861 5134 -827
rect 5328 -725 5362 -691
rect 5328 -793 5362 -759
rect 5328 -861 5362 -827
rect 5586 -725 5620 -691
rect 5586 -793 5620 -759
rect 5586 -861 5620 -827
rect 5780 -725 5814 -691
rect 5780 -793 5814 -759
rect 5780 -861 5814 -827
rect 6038 -725 6072 -691
rect 6038 -793 6072 -759
rect 6038 -861 6072 -827
rect 6296 -725 6330 -691
rect 6296 -793 6330 -759
rect 6296 -861 6330 -827
rect 6554 -725 6588 -691
rect 6554 -793 6588 -759
rect 6554 -861 6588 -827
rect 6812 -725 6846 -691
rect 6812 -793 6846 -759
rect 6812 -861 6846 -827
rect 7006 -725 7040 -691
rect 7006 -793 7040 -759
rect 7006 -861 7040 -827
rect 7264 -725 7298 -691
rect 7264 -793 7298 -759
rect 7264 -861 7298 -827
rect 7522 -725 7556 -691
rect 7522 -793 7556 -759
rect 7522 -861 7556 -827
rect 7780 -725 7814 -691
rect 7780 -793 7814 -759
rect 7780 -861 7814 -827
rect 7974 -725 8008 -691
rect 7974 -793 8008 -759
rect 7974 -861 8008 -827
rect 8232 -725 8266 -691
rect 8232 -793 8266 -759
rect 8232 -861 8266 -827
rect 8490 -725 8524 -691
rect 8490 -793 8524 -759
rect 8490 -861 8524 -827
rect 8748 -725 8782 -691
rect 8748 -793 8782 -759
rect 8748 -861 8782 -827
rect 9006 -725 9040 -691
rect 9006 -793 9040 -759
rect 9006 -861 9040 -827
rect 9200 -725 9234 -691
rect 9200 -793 9234 -759
rect 9200 -861 9234 -827
rect 9458 -725 9492 -691
rect 9458 -793 9492 -759
rect 9458 -861 9492 -827
rect 9688 -725 9722 -691
rect 9688 -793 9722 -759
rect 9688 -861 9722 -827
rect 9946 -725 9980 -691
rect 9946 -793 9980 -759
rect 9946 -861 9980 -827
rect 10140 -725 10174 -691
rect 10140 -793 10174 -759
rect 10140 -861 10174 -827
rect 10398 -725 10432 -691
rect 10398 -793 10432 -759
rect 10398 -861 10432 -827
rect 10656 -725 10690 -691
rect 10656 -793 10690 -759
rect 10656 -861 10690 -827
rect 10914 -725 10948 -691
rect 10914 -793 10948 -759
rect 10914 -861 10948 -827
rect 11172 -725 11206 -691
rect 11172 -793 11206 -759
rect 11172 -861 11206 -827
rect 11366 -725 11400 -691
rect 11366 -793 11400 -759
rect 11366 -861 11400 -827
rect 11624 -725 11658 -691
rect 11624 -793 11658 -759
rect 11624 -861 11658 -827
rect 11882 -725 11916 -691
rect 11882 -793 11916 -759
rect 11882 -861 11916 -827
rect 12140 -725 12174 -691
rect 12140 -793 12174 -759
rect 12140 -861 12174 -827
rect 12334 -725 12368 -691
rect 12334 -793 12368 -759
rect 12334 -861 12368 -827
rect 12592 -725 12626 -691
rect 12592 -793 12626 -759
rect 12592 -861 12626 -827
rect 12850 -725 12884 -691
rect 12850 -793 12884 -759
rect 12850 -861 12884 -827
rect 13108 -725 13142 -691
rect 13108 -793 13142 -759
rect 13108 -861 13142 -827
rect 13366 -725 13400 -691
rect 13366 -793 13400 -759
rect 13366 -861 13400 -827
rect 13560 -725 13594 -691
rect 13560 -793 13594 -759
rect 13560 -861 13594 -827
rect 13818 -725 13852 -691
rect 13818 -793 13852 -759
rect 13818 -861 13852 -827
rect 14046 -725 14080 -691
rect 14046 -793 14080 -759
rect 14046 -861 14080 -827
rect 14304 -725 14338 -691
rect 14304 -793 14338 -759
rect 14304 -861 14338 -827
rect 14497 -725 14531 -691
rect 14497 -793 14531 -759
rect 14497 -861 14531 -827
rect 14755 -725 14789 -691
rect 14755 -793 14789 -759
rect 14755 -861 14789 -827
rect 15013 -725 15047 -691
rect 15013 -793 15047 -759
rect 15013 -861 15047 -827
rect 15271 -725 15305 -691
rect 15271 -793 15305 -759
rect 15271 -861 15305 -827
rect 15529 -725 15563 -691
rect 15529 -793 15563 -759
rect 15529 -861 15563 -827
rect 15723 -725 15757 -691
rect 15723 -793 15757 -759
rect 15723 -861 15757 -827
rect 15981 -725 16015 -691
rect 15981 -793 16015 -759
rect 15981 -861 16015 -827
rect 16239 -725 16273 -691
rect 16239 -793 16273 -759
rect 16239 -861 16273 -827
rect 16497 -725 16531 -691
rect 16497 -793 16531 -759
rect 16497 -861 16531 -827
rect 16691 -725 16725 -691
rect 16691 -793 16725 -759
rect 16691 -861 16725 -827
rect 16949 -725 16983 -691
rect 16949 -793 16983 -759
rect 16949 -861 16983 -827
rect 17207 -725 17241 -691
rect 17207 -793 17241 -759
rect 17207 -861 17241 -827
rect 17465 -725 17499 -691
rect 17465 -793 17499 -759
rect 17465 -861 17499 -827
rect 17723 -725 17757 -691
rect 17723 -793 17757 -759
rect 17723 -861 17757 -827
rect 17917 -725 17951 -691
rect 17917 -793 17951 -759
rect 17917 -861 17951 -827
rect 18175 -725 18209 -691
rect 18175 -793 18209 -759
rect 18175 -861 18209 -827
rect 971 -1416 1005 -1382
rect 971 -1484 1005 -1450
rect 971 -1552 1005 -1518
rect 1229 -1416 1263 -1382
rect 1229 -1484 1263 -1450
rect 1229 -1552 1263 -1518
rect 1423 -1416 1457 -1382
rect 1423 -1484 1457 -1450
rect 1423 -1552 1457 -1518
rect 1681 -1416 1715 -1382
rect 1681 -1484 1715 -1450
rect 1681 -1552 1715 -1518
rect 1939 -1416 1973 -1382
rect 1939 -1484 1973 -1450
rect 1939 -1552 1973 -1518
rect 2197 -1416 2231 -1382
rect 2197 -1484 2231 -1450
rect 2197 -1552 2231 -1518
rect 2455 -1416 2489 -1382
rect 2455 -1484 2489 -1450
rect 2455 -1552 2489 -1518
rect 2649 -1416 2683 -1382
rect 2649 -1484 2683 -1450
rect 2649 -1552 2683 -1518
rect 2907 -1416 2941 -1382
rect 2907 -1484 2941 -1450
rect 2907 -1552 2941 -1518
rect 3165 -1416 3199 -1382
rect 3165 -1484 3199 -1450
rect 3165 -1552 3199 -1518
rect 3423 -1416 3457 -1382
rect 3423 -1484 3457 -1450
rect 3423 -1552 3457 -1518
rect 3617 -1416 3651 -1382
rect 3617 -1484 3651 -1450
rect 3617 -1552 3651 -1518
rect 3875 -1416 3909 -1382
rect 3875 -1484 3909 -1450
rect 3875 -1552 3909 -1518
rect 4133 -1416 4167 -1382
rect 4133 -1484 4167 -1450
rect 4133 -1552 4167 -1518
rect 4391 -1416 4425 -1382
rect 4391 -1484 4425 -1450
rect 4391 -1552 4425 -1518
rect 4649 -1416 4683 -1382
rect 4649 -1484 4683 -1450
rect 4649 -1552 4683 -1518
rect 4842 -1416 4876 -1382
rect 4842 -1484 4876 -1450
rect 4842 -1552 4876 -1518
rect 5100 -1416 5134 -1382
rect 5100 -1484 5134 -1450
rect 5100 -1552 5134 -1518
rect 5328 -1416 5362 -1382
rect 5328 -1484 5362 -1450
rect 5328 -1552 5362 -1518
rect 5586 -1416 5620 -1382
rect 5586 -1484 5620 -1450
rect 5586 -1552 5620 -1518
rect 5780 -1416 5814 -1382
rect 5780 -1484 5814 -1450
rect 5780 -1552 5814 -1518
rect 6038 -1416 6072 -1382
rect 6038 -1484 6072 -1450
rect 6038 -1552 6072 -1518
rect 6296 -1416 6330 -1382
rect 6296 -1484 6330 -1450
rect 6296 -1552 6330 -1518
rect 6554 -1416 6588 -1382
rect 6554 -1484 6588 -1450
rect 6554 -1552 6588 -1518
rect 6812 -1416 6846 -1382
rect 6812 -1484 6846 -1450
rect 6812 -1552 6846 -1518
rect 7006 -1416 7040 -1382
rect 7006 -1484 7040 -1450
rect 7006 -1552 7040 -1518
rect 7264 -1416 7298 -1382
rect 7264 -1484 7298 -1450
rect 7264 -1552 7298 -1518
rect 7522 -1416 7556 -1382
rect 7522 -1484 7556 -1450
rect 7522 -1552 7556 -1518
rect 7780 -1416 7814 -1382
rect 7780 -1484 7814 -1450
rect 7780 -1552 7814 -1518
rect 7974 -1416 8008 -1382
rect 7974 -1484 8008 -1450
rect 7974 -1552 8008 -1518
rect 8232 -1416 8266 -1382
rect 8232 -1484 8266 -1450
rect 8232 -1552 8266 -1518
rect 8490 -1416 8524 -1382
rect 8490 -1484 8524 -1450
rect 8490 -1552 8524 -1518
rect 8748 -1416 8782 -1382
rect 8748 -1484 8782 -1450
rect 8748 -1552 8782 -1518
rect 9006 -1416 9040 -1382
rect 9006 -1484 9040 -1450
rect 9006 -1552 9040 -1518
rect 9200 -1416 9234 -1382
rect 9200 -1484 9234 -1450
rect 9200 -1552 9234 -1518
rect 9458 -1416 9492 -1382
rect 9458 -1484 9492 -1450
rect 9458 -1552 9492 -1518
rect 9688 -1416 9722 -1382
rect 9688 -1484 9722 -1450
rect 9688 -1552 9722 -1518
rect 9946 -1416 9980 -1382
rect 9946 -1484 9980 -1450
rect 9946 -1552 9980 -1518
rect 10140 -1416 10174 -1382
rect 10140 -1484 10174 -1450
rect 10140 -1552 10174 -1518
rect 10398 -1416 10432 -1382
rect 10398 -1484 10432 -1450
rect 10398 -1552 10432 -1518
rect 10656 -1416 10690 -1382
rect 10656 -1484 10690 -1450
rect 10656 -1552 10690 -1518
rect 10914 -1416 10948 -1382
rect 10914 -1484 10948 -1450
rect 10914 -1552 10948 -1518
rect 11172 -1416 11206 -1382
rect 11172 -1484 11206 -1450
rect 11172 -1552 11206 -1518
rect 11366 -1416 11400 -1382
rect 11366 -1484 11400 -1450
rect 11366 -1552 11400 -1518
rect 11624 -1416 11658 -1382
rect 11624 -1484 11658 -1450
rect 11624 -1552 11658 -1518
rect 11882 -1416 11916 -1382
rect 11882 -1484 11916 -1450
rect 11882 -1552 11916 -1518
rect 12140 -1416 12174 -1382
rect 12140 -1484 12174 -1450
rect 12140 -1552 12174 -1518
rect 12334 -1416 12368 -1382
rect 12334 -1484 12368 -1450
rect 12334 -1552 12368 -1518
rect 12592 -1416 12626 -1382
rect 12592 -1484 12626 -1450
rect 12592 -1552 12626 -1518
rect 12850 -1416 12884 -1382
rect 12850 -1484 12884 -1450
rect 12850 -1552 12884 -1518
rect 13108 -1416 13142 -1382
rect 13108 -1484 13142 -1450
rect 13108 -1552 13142 -1518
rect 13366 -1416 13400 -1382
rect 13366 -1484 13400 -1450
rect 13366 -1552 13400 -1518
rect 13560 -1416 13594 -1382
rect 13560 -1484 13594 -1450
rect 13560 -1552 13594 -1518
rect 13818 -1416 13852 -1382
rect 13818 -1484 13852 -1450
rect 13818 -1552 13852 -1518
rect 14046 -1416 14080 -1382
rect 14046 -1484 14080 -1450
rect 14046 -1552 14080 -1518
rect 14304 -1416 14338 -1382
rect 14304 -1484 14338 -1450
rect 14304 -1552 14338 -1518
rect 14497 -1416 14531 -1382
rect 14497 -1484 14531 -1450
rect 14497 -1552 14531 -1518
rect 14755 -1416 14789 -1382
rect 14755 -1484 14789 -1450
rect 14755 -1552 14789 -1518
rect 15013 -1416 15047 -1382
rect 15013 -1484 15047 -1450
rect 15013 -1552 15047 -1518
rect 15271 -1416 15305 -1382
rect 15271 -1484 15305 -1450
rect 15271 -1552 15305 -1518
rect 15529 -1416 15563 -1382
rect 15529 -1484 15563 -1450
rect 15529 -1552 15563 -1518
rect 15723 -1416 15757 -1382
rect 15723 -1484 15757 -1450
rect 15723 -1552 15757 -1518
rect 15981 -1416 16015 -1382
rect 15981 -1484 16015 -1450
rect 15981 -1552 16015 -1518
rect 16239 -1416 16273 -1382
rect 16239 -1484 16273 -1450
rect 16239 -1552 16273 -1518
rect 16497 -1416 16531 -1382
rect 16497 -1484 16531 -1450
rect 16497 -1552 16531 -1518
rect 16691 -1416 16725 -1382
rect 16691 -1484 16725 -1450
rect 16691 -1552 16725 -1518
rect 16949 -1416 16983 -1382
rect 16949 -1484 16983 -1450
rect 16949 -1552 16983 -1518
rect 17207 -1416 17241 -1382
rect 17207 -1484 17241 -1450
rect 17207 -1552 17241 -1518
rect 17465 -1416 17499 -1382
rect 17465 -1484 17499 -1450
rect 17465 -1552 17499 -1518
rect 17723 -1416 17757 -1382
rect 17723 -1484 17757 -1450
rect 17723 -1552 17757 -1518
rect 17917 -1416 17951 -1382
rect 17917 -1484 17951 -1450
rect 17917 -1552 17951 -1518
rect 18175 -1416 18209 -1382
rect 18175 -1484 18209 -1450
rect 18175 -1552 18209 -1518
rect 971 -2372 1005 -2338
rect 971 -2440 1005 -2406
rect 971 -2508 1005 -2474
rect 1229 -2372 1263 -2338
rect 1229 -2440 1263 -2406
rect 1229 -2508 1263 -2474
rect 1423 -2372 1457 -2338
rect 1423 -2440 1457 -2406
rect 1423 -2508 1457 -2474
rect 1681 -2372 1715 -2338
rect 1681 -2440 1715 -2406
rect 1681 -2508 1715 -2474
rect 1939 -2372 1973 -2338
rect 1939 -2440 1973 -2406
rect 1939 -2508 1973 -2474
rect 2197 -2372 2231 -2338
rect 2197 -2440 2231 -2406
rect 2197 -2508 2231 -2474
rect 2455 -2372 2489 -2338
rect 2455 -2440 2489 -2406
rect 2455 -2508 2489 -2474
rect 2649 -2372 2683 -2338
rect 2649 -2440 2683 -2406
rect 2649 -2508 2683 -2474
rect 2907 -2372 2941 -2338
rect 2907 -2440 2941 -2406
rect 2907 -2508 2941 -2474
rect 3165 -2372 3199 -2338
rect 3165 -2440 3199 -2406
rect 3165 -2508 3199 -2474
rect 3423 -2372 3457 -2338
rect 3423 -2440 3457 -2406
rect 3423 -2508 3457 -2474
rect 3617 -2372 3651 -2338
rect 3617 -2440 3651 -2406
rect 3617 -2508 3651 -2474
rect 3875 -2372 3909 -2338
rect 3875 -2440 3909 -2406
rect 3875 -2508 3909 -2474
rect 4133 -2372 4167 -2338
rect 4133 -2440 4167 -2406
rect 4133 -2508 4167 -2474
rect 4391 -2372 4425 -2338
rect 4391 -2440 4425 -2406
rect 4391 -2508 4425 -2474
rect 4649 -2372 4683 -2338
rect 4649 -2440 4683 -2406
rect 4649 -2508 4683 -2474
rect 4842 -2372 4876 -2338
rect 4842 -2440 4876 -2406
rect 4842 -2508 4876 -2474
rect 5100 -2372 5134 -2338
rect 5100 -2440 5134 -2406
rect 5100 -2508 5134 -2474
rect 5328 -2372 5362 -2338
rect 5328 -2440 5362 -2406
rect 5328 -2508 5362 -2474
rect 5586 -2372 5620 -2338
rect 5586 -2440 5620 -2406
rect 5586 -2508 5620 -2474
rect 5780 -2372 5814 -2338
rect 5780 -2440 5814 -2406
rect 5780 -2508 5814 -2474
rect 6038 -2372 6072 -2338
rect 6038 -2440 6072 -2406
rect 6038 -2508 6072 -2474
rect 6296 -2372 6330 -2338
rect 6296 -2440 6330 -2406
rect 6296 -2508 6330 -2474
rect 6554 -2372 6588 -2338
rect 6554 -2440 6588 -2406
rect 6554 -2508 6588 -2474
rect 6812 -2372 6846 -2338
rect 6812 -2440 6846 -2406
rect 6812 -2508 6846 -2474
rect 7006 -2372 7040 -2338
rect 7006 -2440 7040 -2406
rect 7006 -2508 7040 -2474
rect 7264 -2372 7298 -2338
rect 7264 -2440 7298 -2406
rect 7264 -2508 7298 -2474
rect 7522 -2372 7556 -2338
rect 7522 -2440 7556 -2406
rect 7522 -2508 7556 -2474
rect 7780 -2372 7814 -2338
rect 7780 -2440 7814 -2406
rect 7780 -2508 7814 -2474
rect 7974 -2372 8008 -2338
rect 7974 -2440 8008 -2406
rect 7974 -2508 8008 -2474
rect 8232 -2372 8266 -2338
rect 8232 -2440 8266 -2406
rect 8232 -2508 8266 -2474
rect 8490 -2372 8524 -2338
rect 8490 -2440 8524 -2406
rect 8490 -2508 8524 -2474
rect 8748 -2372 8782 -2338
rect 8748 -2440 8782 -2406
rect 8748 -2508 8782 -2474
rect 9006 -2372 9040 -2338
rect 9006 -2440 9040 -2406
rect 9006 -2508 9040 -2474
rect 9200 -2372 9234 -2338
rect 9200 -2440 9234 -2406
rect 9200 -2508 9234 -2474
rect 9458 -2372 9492 -2338
rect 9458 -2440 9492 -2406
rect 9458 -2508 9492 -2474
rect 9688 -2372 9722 -2338
rect 9688 -2440 9722 -2406
rect 9688 -2508 9722 -2474
rect 9946 -2372 9980 -2338
rect 9946 -2440 9980 -2406
rect 9946 -2508 9980 -2474
rect 10140 -2372 10174 -2338
rect 10140 -2440 10174 -2406
rect 10140 -2508 10174 -2474
rect 10398 -2372 10432 -2338
rect 10398 -2440 10432 -2406
rect 10398 -2508 10432 -2474
rect 10656 -2372 10690 -2338
rect 10656 -2440 10690 -2406
rect 10656 -2508 10690 -2474
rect 10914 -2372 10948 -2338
rect 10914 -2440 10948 -2406
rect 10914 -2508 10948 -2474
rect 11172 -2372 11206 -2338
rect 11172 -2440 11206 -2406
rect 11172 -2508 11206 -2474
rect 11366 -2372 11400 -2338
rect 11366 -2440 11400 -2406
rect 11366 -2508 11400 -2474
rect 11624 -2372 11658 -2338
rect 11624 -2440 11658 -2406
rect 11624 -2508 11658 -2474
rect 11882 -2372 11916 -2338
rect 11882 -2440 11916 -2406
rect 11882 -2508 11916 -2474
rect 12140 -2372 12174 -2338
rect 12140 -2440 12174 -2406
rect 12140 -2508 12174 -2474
rect 12334 -2372 12368 -2338
rect 12334 -2440 12368 -2406
rect 12334 -2508 12368 -2474
rect 12592 -2372 12626 -2338
rect 12592 -2440 12626 -2406
rect 12592 -2508 12626 -2474
rect 12850 -2372 12884 -2338
rect 12850 -2440 12884 -2406
rect 12850 -2508 12884 -2474
rect 13108 -2372 13142 -2338
rect 13108 -2440 13142 -2406
rect 13108 -2508 13142 -2474
rect 13366 -2372 13400 -2338
rect 13366 -2440 13400 -2406
rect 13366 -2508 13400 -2474
rect 13560 -2372 13594 -2338
rect 13560 -2440 13594 -2406
rect 13560 -2508 13594 -2474
rect 13818 -2372 13852 -2338
rect 13818 -2440 13852 -2406
rect 13818 -2508 13852 -2474
rect 14046 -2372 14080 -2338
rect 14046 -2440 14080 -2406
rect 14046 -2508 14080 -2474
rect 14304 -2372 14338 -2338
rect 14304 -2440 14338 -2406
rect 14304 -2508 14338 -2474
rect 14497 -2372 14531 -2338
rect 14497 -2440 14531 -2406
rect 14497 -2508 14531 -2474
rect 14755 -2372 14789 -2338
rect 14755 -2440 14789 -2406
rect 14755 -2508 14789 -2474
rect 15013 -2372 15047 -2338
rect 15013 -2440 15047 -2406
rect 15013 -2508 15047 -2474
rect 15271 -2372 15305 -2338
rect 15271 -2440 15305 -2406
rect 15271 -2508 15305 -2474
rect 15529 -2372 15563 -2338
rect 15529 -2440 15563 -2406
rect 15529 -2508 15563 -2474
rect 15723 -2372 15757 -2338
rect 15723 -2440 15757 -2406
rect 15723 -2508 15757 -2474
rect 15981 -2372 16015 -2338
rect 15981 -2440 16015 -2406
rect 15981 -2508 16015 -2474
rect 16239 -2372 16273 -2338
rect 16239 -2440 16273 -2406
rect 16239 -2508 16273 -2474
rect 16497 -2372 16531 -2338
rect 16497 -2440 16531 -2406
rect 16497 -2508 16531 -2474
rect 16691 -2372 16725 -2338
rect 16691 -2440 16725 -2406
rect 16691 -2508 16725 -2474
rect 16949 -2372 16983 -2338
rect 16949 -2440 16983 -2406
rect 16949 -2508 16983 -2474
rect 17207 -2372 17241 -2338
rect 17207 -2440 17241 -2406
rect 17207 -2508 17241 -2474
rect 17465 -2372 17499 -2338
rect 17465 -2440 17499 -2406
rect 17465 -2508 17499 -2474
rect 17723 -2372 17757 -2338
rect 17723 -2440 17757 -2406
rect 17723 -2508 17757 -2474
rect 17917 -2372 17951 -2338
rect 17917 -2440 17951 -2406
rect 17917 -2508 17951 -2474
rect 18175 -2372 18209 -2338
rect 18175 -2440 18209 -2406
rect 18175 -2508 18209 -2474
rect 971 -3063 1005 -3029
rect 971 -3131 1005 -3097
rect 971 -3199 1005 -3165
rect 1229 -3063 1263 -3029
rect 1229 -3131 1263 -3097
rect 1229 -3199 1263 -3165
rect 1423 -3063 1457 -3029
rect 1423 -3131 1457 -3097
rect 1423 -3199 1457 -3165
rect 1681 -3063 1715 -3029
rect 1681 -3131 1715 -3097
rect 1681 -3199 1715 -3165
rect 1939 -3063 1973 -3029
rect 1939 -3131 1973 -3097
rect 1939 -3199 1973 -3165
rect 2197 -3063 2231 -3029
rect 2197 -3131 2231 -3097
rect 2197 -3199 2231 -3165
rect 2455 -3063 2489 -3029
rect 2455 -3131 2489 -3097
rect 2455 -3199 2489 -3165
rect 2649 -3063 2683 -3029
rect 2649 -3131 2683 -3097
rect 2649 -3199 2683 -3165
rect 2907 -3063 2941 -3029
rect 2907 -3131 2941 -3097
rect 2907 -3199 2941 -3165
rect 3165 -3063 3199 -3029
rect 3165 -3131 3199 -3097
rect 3165 -3199 3199 -3165
rect 3423 -3063 3457 -3029
rect 3423 -3131 3457 -3097
rect 3423 -3199 3457 -3165
rect 3617 -3063 3651 -3029
rect 3617 -3131 3651 -3097
rect 3617 -3199 3651 -3165
rect 3875 -3063 3909 -3029
rect 3875 -3131 3909 -3097
rect 3875 -3199 3909 -3165
rect 4133 -3063 4167 -3029
rect 4133 -3131 4167 -3097
rect 4133 -3199 4167 -3165
rect 4391 -3063 4425 -3029
rect 4391 -3131 4425 -3097
rect 4391 -3199 4425 -3165
rect 4649 -3063 4683 -3029
rect 4649 -3131 4683 -3097
rect 4649 -3199 4683 -3165
rect 4842 -3063 4876 -3029
rect 4842 -3131 4876 -3097
rect 4842 -3199 4876 -3165
rect 5100 -3063 5134 -3029
rect 5100 -3131 5134 -3097
rect 5100 -3199 5134 -3165
rect 5328 -3063 5362 -3029
rect 5328 -3131 5362 -3097
rect 5328 -3199 5362 -3165
rect 5586 -3063 5620 -3029
rect 5586 -3131 5620 -3097
rect 5586 -3199 5620 -3165
rect 5780 -3063 5814 -3029
rect 5780 -3131 5814 -3097
rect 5780 -3199 5814 -3165
rect 6038 -3063 6072 -3029
rect 6038 -3131 6072 -3097
rect 6038 -3199 6072 -3165
rect 6296 -3063 6330 -3029
rect 6296 -3131 6330 -3097
rect 6296 -3199 6330 -3165
rect 6554 -3063 6588 -3029
rect 6554 -3131 6588 -3097
rect 6554 -3199 6588 -3165
rect 6812 -3063 6846 -3029
rect 6812 -3131 6846 -3097
rect 6812 -3199 6846 -3165
rect 7006 -3063 7040 -3029
rect 7006 -3131 7040 -3097
rect 7006 -3199 7040 -3165
rect 7264 -3063 7298 -3029
rect 7264 -3131 7298 -3097
rect 7264 -3199 7298 -3165
rect 7522 -3063 7556 -3029
rect 7522 -3131 7556 -3097
rect 7522 -3199 7556 -3165
rect 7780 -3063 7814 -3029
rect 7780 -3131 7814 -3097
rect 7780 -3199 7814 -3165
rect 7974 -3063 8008 -3029
rect 7974 -3131 8008 -3097
rect 7974 -3199 8008 -3165
rect 8232 -3063 8266 -3029
rect 8232 -3131 8266 -3097
rect 8232 -3199 8266 -3165
rect 8490 -3063 8524 -3029
rect 8490 -3131 8524 -3097
rect 8490 -3199 8524 -3165
rect 8748 -3063 8782 -3029
rect 8748 -3131 8782 -3097
rect 8748 -3199 8782 -3165
rect 9006 -3063 9040 -3029
rect 9006 -3131 9040 -3097
rect 9006 -3199 9040 -3165
rect 9200 -3063 9234 -3029
rect 9200 -3131 9234 -3097
rect 9200 -3199 9234 -3165
rect 9458 -3063 9492 -3029
rect 9458 -3131 9492 -3097
rect 9458 -3199 9492 -3165
rect 9688 -3063 9722 -3029
rect 9688 -3131 9722 -3097
rect 9688 -3199 9722 -3165
rect 9946 -3063 9980 -3029
rect 9946 -3131 9980 -3097
rect 9946 -3199 9980 -3165
rect 10140 -3063 10174 -3029
rect 10140 -3131 10174 -3097
rect 10140 -3199 10174 -3165
rect 10398 -3063 10432 -3029
rect 10398 -3131 10432 -3097
rect 10398 -3199 10432 -3165
rect 10656 -3063 10690 -3029
rect 10656 -3131 10690 -3097
rect 10656 -3199 10690 -3165
rect 10914 -3063 10948 -3029
rect 10914 -3131 10948 -3097
rect 10914 -3199 10948 -3165
rect 11172 -3063 11206 -3029
rect 11172 -3131 11206 -3097
rect 11172 -3199 11206 -3165
rect 11366 -3063 11400 -3029
rect 11366 -3131 11400 -3097
rect 11366 -3199 11400 -3165
rect 11624 -3063 11658 -3029
rect 11624 -3131 11658 -3097
rect 11624 -3199 11658 -3165
rect 11882 -3063 11916 -3029
rect 11882 -3131 11916 -3097
rect 11882 -3199 11916 -3165
rect 12140 -3063 12174 -3029
rect 12140 -3131 12174 -3097
rect 12140 -3199 12174 -3165
rect 12334 -3063 12368 -3029
rect 12334 -3131 12368 -3097
rect 12334 -3199 12368 -3165
rect 12592 -3063 12626 -3029
rect 12592 -3131 12626 -3097
rect 12592 -3199 12626 -3165
rect 12850 -3063 12884 -3029
rect 12850 -3131 12884 -3097
rect 12850 -3199 12884 -3165
rect 13108 -3063 13142 -3029
rect 13108 -3131 13142 -3097
rect 13108 -3199 13142 -3165
rect 13366 -3063 13400 -3029
rect 13366 -3131 13400 -3097
rect 13366 -3199 13400 -3165
rect 13560 -3063 13594 -3029
rect 13560 -3131 13594 -3097
rect 13560 -3199 13594 -3165
rect 13818 -3063 13852 -3029
rect 13818 -3131 13852 -3097
rect 13818 -3199 13852 -3165
rect 14046 -3063 14080 -3029
rect 14046 -3131 14080 -3097
rect 14046 -3199 14080 -3165
rect 14304 -3063 14338 -3029
rect 14304 -3131 14338 -3097
rect 14304 -3199 14338 -3165
rect 14497 -3063 14531 -3029
rect 14497 -3131 14531 -3097
rect 14497 -3199 14531 -3165
rect 14755 -3063 14789 -3029
rect 14755 -3131 14789 -3097
rect 14755 -3199 14789 -3165
rect 15013 -3063 15047 -3029
rect 15013 -3131 15047 -3097
rect 15013 -3199 15047 -3165
rect 15271 -3063 15305 -3029
rect 15271 -3131 15305 -3097
rect 15271 -3199 15305 -3165
rect 15529 -3063 15563 -3029
rect 15529 -3131 15563 -3097
rect 15529 -3199 15563 -3165
rect 15723 -3063 15757 -3029
rect 15723 -3131 15757 -3097
rect 15723 -3199 15757 -3165
rect 15981 -3063 16015 -3029
rect 15981 -3131 16015 -3097
rect 15981 -3199 16015 -3165
rect 16239 -3063 16273 -3029
rect 16239 -3131 16273 -3097
rect 16239 -3199 16273 -3165
rect 16497 -3063 16531 -3029
rect 16497 -3131 16531 -3097
rect 16497 -3199 16531 -3165
rect 16691 -3063 16725 -3029
rect 16691 -3131 16725 -3097
rect 16691 -3199 16725 -3165
rect 16949 -3063 16983 -3029
rect 16949 -3131 16983 -3097
rect 16949 -3199 16983 -3165
rect 17207 -3063 17241 -3029
rect 17207 -3131 17241 -3097
rect 17207 -3199 17241 -3165
rect 17465 -3063 17499 -3029
rect 17465 -3131 17499 -3097
rect 17465 -3199 17499 -3165
rect 17723 -3063 17757 -3029
rect 17723 -3131 17757 -3097
rect 17723 -3199 17757 -3165
rect 17917 -3063 17951 -3029
rect 17917 -3131 17951 -3097
rect 17917 -3199 17951 -3165
rect 18175 -3063 18209 -3029
rect 18175 -3131 18209 -3097
rect 18175 -3199 18209 -3165
rect 971 -4053 1005 -4019
rect 971 -4121 1005 -4087
rect 971 -4189 1005 -4155
rect 1229 -4053 1263 -4019
rect 1229 -4121 1263 -4087
rect 1229 -4189 1263 -4155
rect 1423 -4053 1457 -4019
rect 1423 -4121 1457 -4087
rect 1423 -4189 1457 -4155
rect 1681 -4053 1715 -4019
rect 1681 -4121 1715 -4087
rect 1681 -4189 1715 -4155
rect 1939 -4053 1973 -4019
rect 1939 -4121 1973 -4087
rect 1939 -4189 1973 -4155
rect 2197 -4053 2231 -4019
rect 2197 -4121 2231 -4087
rect 2197 -4189 2231 -4155
rect 2455 -4053 2489 -4019
rect 2455 -4121 2489 -4087
rect 2455 -4189 2489 -4155
rect 2649 -4053 2683 -4019
rect 2649 -4121 2683 -4087
rect 2649 -4189 2683 -4155
rect 2907 -4053 2941 -4019
rect 2907 -4121 2941 -4087
rect 2907 -4189 2941 -4155
rect 3165 -4053 3199 -4019
rect 3165 -4121 3199 -4087
rect 3165 -4189 3199 -4155
rect 3423 -4053 3457 -4019
rect 3423 -4121 3457 -4087
rect 3423 -4189 3457 -4155
rect 3617 -4053 3651 -4019
rect 3617 -4121 3651 -4087
rect 3617 -4189 3651 -4155
rect 3875 -4053 3909 -4019
rect 3875 -4121 3909 -4087
rect 3875 -4189 3909 -4155
rect 4133 -4053 4167 -4019
rect 4133 -4121 4167 -4087
rect 4133 -4189 4167 -4155
rect 4391 -4053 4425 -4019
rect 4391 -4121 4425 -4087
rect 4391 -4189 4425 -4155
rect 4649 -4053 4683 -4019
rect 4649 -4121 4683 -4087
rect 4649 -4189 4683 -4155
rect 4842 -4053 4876 -4019
rect 4842 -4121 4876 -4087
rect 4842 -4189 4876 -4155
rect 5100 -4053 5134 -4019
rect 5100 -4121 5134 -4087
rect 5100 -4189 5134 -4155
rect 5328 -4053 5362 -4019
rect 5328 -4121 5362 -4087
rect 5328 -4189 5362 -4155
rect 5586 -4053 5620 -4019
rect 5586 -4121 5620 -4087
rect 5586 -4189 5620 -4155
rect 5780 -4053 5814 -4019
rect 5780 -4121 5814 -4087
rect 5780 -4189 5814 -4155
rect 6038 -4053 6072 -4019
rect 6038 -4121 6072 -4087
rect 6038 -4189 6072 -4155
rect 6296 -4053 6330 -4019
rect 6296 -4121 6330 -4087
rect 6296 -4189 6330 -4155
rect 6554 -4053 6588 -4019
rect 6554 -4121 6588 -4087
rect 6554 -4189 6588 -4155
rect 6812 -4053 6846 -4019
rect 6812 -4121 6846 -4087
rect 6812 -4189 6846 -4155
rect 7006 -4053 7040 -4019
rect 7006 -4121 7040 -4087
rect 7006 -4189 7040 -4155
rect 7264 -4053 7298 -4019
rect 7264 -4121 7298 -4087
rect 7264 -4189 7298 -4155
rect 7522 -4053 7556 -4019
rect 7522 -4121 7556 -4087
rect 7522 -4189 7556 -4155
rect 7780 -4053 7814 -4019
rect 7780 -4121 7814 -4087
rect 7780 -4189 7814 -4155
rect 7974 -4053 8008 -4019
rect 7974 -4121 8008 -4087
rect 7974 -4189 8008 -4155
rect 8232 -4053 8266 -4019
rect 8232 -4121 8266 -4087
rect 8232 -4189 8266 -4155
rect 8490 -4053 8524 -4019
rect 8490 -4121 8524 -4087
rect 8490 -4189 8524 -4155
rect 8748 -4053 8782 -4019
rect 8748 -4121 8782 -4087
rect 8748 -4189 8782 -4155
rect 9006 -4053 9040 -4019
rect 9006 -4121 9040 -4087
rect 9006 -4189 9040 -4155
rect 9200 -4053 9234 -4019
rect 9200 -4121 9234 -4087
rect 9200 -4189 9234 -4155
rect 9458 -4053 9492 -4019
rect 9458 -4121 9492 -4087
rect 9458 -4189 9492 -4155
rect 9688 -4053 9722 -4019
rect 9688 -4121 9722 -4087
rect 9688 -4189 9722 -4155
rect 9946 -4053 9980 -4019
rect 9946 -4121 9980 -4087
rect 9946 -4189 9980 -4155
rect 10140 -4053 10174 -4019
rect 10140 -4121 10174 -4087
rect 10140 -4189 10174 -4155
rect 10398 -4053 10432 -4019
rect 10398 -4121 10432 -4087
rect 10398 -4189 10432 -4155
rect 10656 -4053 10690 -4019
rect 10656 -4121 10690 -4087
rect 10656 -4189 10690 -4155
rect 10914 -4053 10948 -4019
rect 10914 -4121 10948 -4087
rect 10914 -4189 10948 -4155
rect 11172 -4053 11206 -4019
rect 11172 -4121 11206 -4087
rect 11172 -4189 11206 -4155
rect 11366 -4053 11400 -4019
rect 11366 -4121 11400 -4087
rect 11366 -4189 11400 -4155
rect 11624 -4053 11658 -4019
rect 11624 -4121 11658 -4087
rect 11624 -4189 11658 -4155
rect 11882 -4053 11916 -4019
rect 11882 -4121 11916 -4087
rect 11882 -4189 11916 -4155
rect 12140 -4053 12174 -4019
rect 12140 -4121 12174 -4087
rect 12140 -4189 12174 -4155
rect 12334 -4053 12368 -4019
rect 12334 -4121 12368 -4087
rect 12334 -4189 12368 -4155
rect 12592 -4053 12626 -4019
rect 12592 -4121 12626 -4087
rect 12592 -4189 12626 -4155
rect 12850 -4053 12884 -4019
rect 12850 -4121 12884 -4087
rect 12850 -4189 12884 -4155
rect 13108 -4053 13142 -4019
rect 13108 -4121 13142 -4087
rect 13108 -4189 13142 -4155
rect 13366 -4053 13400 -4019
rect 13366 -4121 13400 -4087
rect 13366 -4189 13400 -4155
rect 13560 -4053 13594 -4019
rect 13560 -4121 13594 -4087
rect 13560 -4189 13594 -4155
rect 13818 -4053 13852 -4019
rect 13818 -4121 13852 -4087
rect 13818 -4189 13852 -4155
rect 14046 -4053 14080 -4019
rect 14046 -4121 14080 -4087
rect 14046 -4189 14080 -4155
rect 14304 -4053 14338 -4019
rect 14304 -4121 14338 -4087
rect 14304 -4189 14338 -4155
rect 14497 -4053 14531 -4019
rect 14497 -4121 14531 -4087
rect 14497 -4189 14531 -4155
rect 14755 -4053 14789 -4019
rect 14755 -4121 14789 -4087
rect 14755 -4189 14789 -4155
rect 15013 -4053 15047 -4019
rect 15013 -4121 15047 -4087
rect 15013 -4189 15047 -4155
rect 15271 -4053 15305 -4019
rect 15271 -4121 15305 -4087
rect 15271 -4189 15305 -4155
rect 15529 -4053 15563 -4019
rect 15529 -4121 15563 -4087
rect 15529 -4189 15563 -4155
rect 15723 -4053 15757 -4019
rect 15723 -4121 15757 -4087
rect 15723 -4189 15757 -4155
rect 15981 -4053 16015 -4019
rect 15981 -4121 16015 -4087
rect 15981 -4189 16015 -4155
rect 16239 -4053 16273 -4019
rect 16239 -4121 16273 -4087
rect 16239 -4189 16273 -4155
rect 16497 -4053 16531 -4019
rect 16497 -4121 16531 -4087
rect 16497 -4189 16531 -4155
rect 16691 -4053 16725 -4019
rect 16691 -4121 16725 -4087
rect 16691 -4189 16725 -4155
rect 16949 -4053 16983 -4019
rect 16949 -4121 16983 -4087
rect 16949 -4189 16983 -4155
rect 17207 -4053 17241 -4019
rect 17207 -4121 17241 -4087
rect 17207 -4189 17241 -4155
rect 17465 -4053 17499 -4019
rect 17465 -4121 17499 -4087
rect 17465 -4189 17499 -4155
rect 17723 -4053 17757 -4019
rect 17723 -4121 17757 -4087
rect 17723 -4189 17757 -4155
rect 17917 -4053 17951 -4019
rect 17917 -4121 17951 -4087
rect 17917 -4189 17951 -4155
rect 18175 -4053 18209 -4019
rect 18175 -4121 18209 -4087
rect 18175 -4189 18209 -4155
rect 971 -4609 1005 -4575
rect 971 -4677 1005 -4643
rect 971 -4745 1005 -4711
rect 1229 -4609 1263 -4575
rect 1229 -4677 1263 -4643
rect 1229 -4745 1263 -4711
rect 1423 -4609 1457 -4575
rect 1423 -4677 1457 -4643
rect 1423 -4745 1457 -4711
rect 1681 -4609 1715 -4575
rect 1681 -4677 1715 -4643
rect 1681 -4745 1715 -4711
rect 1939 -4609 1973 -4575
rect 1939 -4677 1973 -4643
rect 1939 -4745 1973 -4711
rect 2197 -4609 2231 -4575
rect 2197 -4677 2231 -4643
rect 2197 -4745 2231 -4711
rect 2455 -4609 2489 -4575
rect 2455 -4677 2489 -4643
rect 2455 -4745 2489 -4711
rect 2649 -4609 2683 -4575
rect 2649 -4677 2683 -4643
rect 2649 -4745 2683 -4711
rect 2907 -4609 2941 -4575
rect 2907 -4677 2941 -4643
rect 2907 -4745 2941 -4711
rect 3165 -4609 3199 -4575
rect 3165 -4677 3199 -4643
rect 3165 -4745 3199 -4711
rect 3423 -4609 3457 -4575
rect 3423 -4677 3457 -4643
rect 3423 -4745 3457 -4711
rect 3617 -4609 3651 -4575
rect 3617 -4677 3651 -4643
rect 3617 -4745 3651 -4711
rect 3875 -4609 3909 -4575
rect 3875 -4677 3909 -4643
rect 3875 -4745 3909 -4711
rect 4133 -4609 4167 -4575
rect 4133 -4677 4167 -4643
rect 4133 -4745 4167 -4711
rect 4391 -4609 4425 -4575
rect 4391 -4677 4425 -4643
rect 4391 -4745 4425 -4711
rect 4649 -4609 4683 -4575
rect 4649 -4677 4683 -4643
rect 4649 -4745 4683 -4711
rect 4842 -4609 4876 -4575
rect 4842 -4677 4876 -4643
rect 4842 -4745 4876 -4711
rect 5100 -4609 5134 -4575
rect 5100 -4677 5134 -4643
rect 5100 -4745 5134 -4711
rect 5328 -4609 5362 -4575
rect 5328 -4677 5362 -4643
rect 5328 -4745 5362 -4711
rect 5586 -4609 5620 -4575
rect 5586 -4677 5620 -4643
rect 5586 -4745 5620 -4711
rect 5780 -4609 5814 -4575
rect 5780 -4677 5814 -4643
rect 5780 -4745 5814 -4711
rect 6038 -4609 6072 -4575
rect 6038 -4677 6072 -4643
rect 6038 -4745 6072 -4711
rect 6296 -4609 6330 -4575
rect 6296 -4677 6330 -4643
rect 6296 -4745 6330 -4711
rect 6554 -4609 6588 -4575
rect 6554 -4677 6588 -4643
rect 6554 -4745 6588 -4711
rect 6812 -4609 6846 -4575
rect 6812 -4677 6846 -4643
rect 6812 -4745 6846 -4711
rect 7006 -4609 7040 -4575
rect 7006 -4677 7040 -4643
rect 7006 -4745 7040 -4711
rect 7264 -4609 7298 -4575
rect 7264 -4677 7298 -4643
rect 7264 -4745 7298 -4711
rect 7522 -4609 7556 -4575
rect 7522 -4677 7556 -4643
rect 7522 -4745 7556 -4711
rect 7780 -4609 7814 -4575
rect 7780 -4677 7814 -4643
rect 7780 -4745 7814 -4711
rect 7974 -4609 8008 -4575
rect 7974 -4677 8008 -4643
rect 7974 -4745 8008 -4711
rect 8232 -4609 8266 -4575
rect 8232 -4677 8266 -4643
rect 8232 -4745 8266 -4711
rect 8490 -4609 8524 -4575
rect 8490 -4677 8524 -4643
rect 8490 -4745 8524 -4711
rect 8748 -4609 8782 -4575
rect 8748 -4677 8782 -4643
rect 8748 -4745 8782 -4711
rect 9006 -4609 9040 -4575
rect 9006 -4677 9040 -4643
rect 9006 -4745 9040 -4711
rect 9200 -4609 9234 -4575
rect 9200 -4677 9234 -4643
rect 9200 -4745 9234 -4711
rect 9458 -4609 9492 -4575
rect 9458 -4677 9492 -4643
rect 9458 -4745 9492 -4711
rect 9688 -4609 9722 -4575
rect 9688 -4677 9722 -4643
rect 9688 -4745 9722 -4711
rect 9946 -4609 9980 -4575
rect 9946 -4677 9980 -4643
rect 9946 -4745 9980 -4711
rect 10140 -4609 10174 -4575
rect 10140 -4677 10174 -4643
rect 10140 -4745 10174 -4711
rect 10398 -4609 10432 -4575
rect 10398 -4677 10432 -4643
rect 10398 -4745 10432 -4711
rect 10656 -4609 10690 -4575
rect 10656 -4677 10690 -4643
rect 10656 -4745 10690 -4711
rect 10914 -4609 10948 -4575
rect 10914 -4677 10948 -4643
rect 10914 -4745 10948 -4711
rect 11172 -4609 11206 -4575
rect 11172 -4677 11206 -4643
rect 11172 -4745 11206 -4711
rect 11366 -4609 11400 -4575
rect 11366 -4677 11400 -4643
rect 11366 -4745 11400 -4711
rect 11624 -4609 11658 -4575
rect 11624 -4677 11658 -4643
rect 11624 -4745 11658 -4711
rect 11882 -4609 11916 -4575
rect 11882 -4677 11916 -4643
rect 11882 -4745 11916 -4711
rect 12140 -4609 12174 -4575
rect 12140 -4677 12174 -4643
rect 12140 -4745 12174 -4711
rect 12334 -4609 12368 -4575
rect 12334 -4677 12368 -4643
rect 12334 -4745 12368 -4711
rect 12592 -4609 12626 -4575
rect 12592 -4677 12626 -4643
rect 12592 -4745 12626 -4711
rect 12850 -4609 12884 -4575
rect 12850 -4677 12884 -4643
rect 12850 -4745 12884 -4711
rect 13108 -4609 13142 -4575
rect 13108 -4677 13142 -4643
rect 13108 -4745 13142 -4711
rect 13366 -4609 13400 -4575
rect 13366 -4677 13400 -4643
rect 13366 -4745 13400 -4711
rect 13560 -4609 13594 -4575
rect 13560 -4677 13594 -4643
rect 13560 -4745 13594 -4711
rect 13818 -4609 13852 -4575
rect 13818 -4677 13852 -4643
rect 13818 -4745 13852 -4711
rect 14046 -4609 14080 -4575
rect 14046 -4677 14080 -4643
rect 14046 -4745 14080 -4711
rect 14304 -4609 14338 -4575
rect 14304 -4677 14338 -4643
rect 14304 -4745 14338 -4711
rect 14497 -4609 14531 -4575
rect 14497 -4677 14531 -4643
rect 14497 -4745 14531 -4711
rect 14755 -4609 14789 -4575
rect 14755 -4677 14789 -4643
rect 14755 -4745 14789 -4711
rect 15013 -4609 15047 -4575
rect 15013 -4677 15047 -4643
rect 15013 -4745 15047 -4711
rect 15271 -4609 15305 -4575
rect 15271 -4677 15305 -4643
rect 15271 -4745 15305 -4711
rect 15529 -4609 15563 -4575
rect 15529 -4677 15563 -4643
rect 15529 -4745 15563 -4711
rect 15723 -4609 15757 -4575
rect 15723 -4677 15757 -4643
rect 15723 -4745 15757 -4711
rect 15981 -4609 16015 -4575
rect 15981 -4677 16015 -4643
rect 15981 -4745 16015 -4711
rect 16239 -4609 16273 -4575
rect 16239 -4677 16273 -4643
rect 16239 -4745 16273 -4711
rect 16497 -4609 16531 -4575
rect 16497 -4677 16531 -4643
rect 16497 -4745 16531 -4711
rect 16691 -4609 16725 -4575
rect 16691 -4677 16725 -4643
rect 16691 -4745 16725 -4711
rect 16949 -4609 16983 -4575
rect 16949 -4677 16983 -4643
rect 16949 -4745 16983 -4711
rect 17207 -4609 17241 -4575
rect 17207 -4677 17241 -4643
rect 17207 -4745 17241 -4711
rect 17465 -4609 17499 -4575
rect 17465 -4677 17499 -4643
rect 17465 -4745 17499 -4711
rect 17723 -4609 17757 -4575
rect 17723 -4677 17757 -4643
rect 17723 -4745 17757 -4711
rect 17917 -4609 17951 -4575
rect 17917 -4677 17951 -4643
rect 17917 -4745 17951 -4711
rect 18175 -4609 18209 -4575
rect 18175 -4677 18209 -4643
rect 18175 -4745 18209 -4711
rect 971 -5599 1005 -5565
rect 971 -5667 1005 -5633
rect 971 -5735 1005 -5701
rect 1229 -5599 1263 -5565
rect 1229 -5667 1263 -5633
rect 1229 -5735 1263 -5701
rect 1423 -5599 1457 -5565
rect 1423 -5667 1457 -5633
rect 1423 -5735 1457 -5701
rect 1681 -5599 1715 -5565
rect 1681 -5667 1715 -5633
rect 1681 -5735 1715 -5701
rect 1939 -5599 1973 -5565
rect 1939 -5667 1973 -5633
rect 1939 -5735 1973 -5701
rect 2197 -5599 2231 -5565
rect 2197 -5667 2231 -5633
rect 2197 -5735 2231 -5701
rect 2455 -5599 2489 -5565
rect 2455 -5667 2489 -5633
rect 2455 -5735 2489 -5701
rect 2649 -5599 2683 -5565
rect 2649 -5667 2683 -5633
rect 2649 -5735 2683 -5701
rect 2907 -5599 2941 -5565
rect 2907 -5667 2941 -5633
rect 2907 -5735 2941 -5701
rect 3165 -5599 3199 -5565
rect 3165 -5667 3199 -5633
rect 3165 -5735 3199 -5701
rect 3423 -5599 3457 -5565
rect 3423 -5667 3457 -5633
rect 3423 -5735 3457 -5701
rect 3617 -5599 3651 -5565
rect 3617 -5667 3651 -5633
rect 3617 -5735 3651 -5701
rect 3875 -5599 3909 -5565
rect 3875 -5667 3909 -5633
rect 3875 -5735 3909 -5701
rect 4133 -5599 4167 -5565
rect 4133 -5667 4167 -5633
rect 4133 -5735 4167 -5701
rect 4391 -5599 4425 -5565
rect 4391 -5667 4425 -5633
rect 4391 -5735 4425 -5701
rect 4649 -5599 4683 -5565
rect 4649 -5667 4683 -5633
rect 4649 -5735 4683 -5701
rect 4842 -5599 4876 -5565
rect 4842 -5667 4876 -5633
rect 4842 -5735 4876 -5701
rect 5100 -5599 5134 -5565
rect 5100 -5667 5134 -5633
rect 5100 -5735 5134 -5701
rect 5328 -5599 5362 -5565
rect 5328 -5667 5362 -5633
rect 5328 -5735 5362 -5701
rect 5586 -5599 5620 -5565
rect 5586 -5667 5620 -5633
rect 5586 -5735 5620 -5701
rect 5780 -5599 5814 -5565
rect 5780 -5667 5814 -5633
rect 5780 -5735 5814 -5701
rect 6038 -5599 6072 -5565
rect 6038 -5667 6072 -5633
rect 6038 -5735 6072 -5701
rect 6296 -5599 6330 -5565
rect 6296 -5667 6330 -5633
rect 6296 -5735 6330 -5701
rect 6554 -5599 6588 -5565
rect 6554 -5667 6588 -5633
rect 6554 -5735 6588 -5701
rect 6812 -5599 6846 -5565
rect 6812 -5667 6846 -5633
rect 6812 -5735 6846 -5701
rect 7006 -5599 7040 -5565
rect 7006 -5667 7040 -5633
rect 7006 -5735 7040 -5701
rect 7264 -5599 7298 -5565
rect 7264 -5667 7298 -5633
rect 7264 -5735 7298 -5701
rect 7522 -5599 7556 -5565
rect 7522 -5667 7556 -5633
rect 7522 -5735 7556 -5701
rect 7780 -5599 7814 -5565
rect 7780 -5667 7814 -5633
rect 7780 -5735 7814 -5701
rect 7974 -5599 8008 -5565
rect 7974 -5667 8008 -5633
rect 7974 -5735 8008 -5701
rect 8232 -5599 8266 -5565
rect 8232 -5667 8266 -5633
rect 8232 -5735 8266 -5701
rect 8490 -5599 8524 -5565
rect 8490 -5667 8524 -5633
rect 8490 -5735 8524 -5701
rect 8748 -5599 8782 -5565
rect 8748 -5667 8782 -5633
rect 8748 -5735 8782 -5701
rect 9006 -5599 9040 -5565
rect 9006 -5667 9040 -5633
rect 9006 -5735 9040 -5701
rect 9200 -5599 9234 -5565
rect 9200 -5667 9234 -5633
rect 9200 -5735 9234 -5701
rect 9458 -5599 9492 -5565
rect 9458 -5667 9492 -5633
rect 9458 -5735 9492 -5701
rect 9688 -5599 9722 -5565
rect 9688 -5667 9722 -5633
rect 9688 -5735 9722 -5701
rect 9946 -5599 9980 -5565
rect 9946 -5667 9980 -5633
rect 9946 -5735 9980 -5701
rect 10140 -5599 10174 -5565
rect 10140 -5667 10174 -5633
rect 10140 -5735 10174 -5701
rect 10398 -5599 10432 -5565
rect 10398 -5667 10432 -5633
rect 10398 -5735 10432 -5701
rect 10656 -5599 10690 -5565
rect 10656 -5667 10690 -5633
rect 10656 -5735 10690 -5701
rect 10914 -5599 10948 -5565
rect 10914 -5667 10948 -5633
rect 10914 -5735 10948 -5701
rect 11172 -5599 11206 -5565
rect 11172 -5667 11206 -5633
rect 11172 -5735 11206 -5701
rect 11366 -5599 11400 -5565
rect 11366 -5667 11400 -5633
rect 11366 -5735 11400 -5701
rect 11624 -5599 11658 -5565
rect 11624 -5667 11658 -5633
rect 11624 -5735 11658 -5701
rect 11882 -5599 11916 -5565
rect 11882 -5667 11916 -5633
rect 11882 -5735 11916 -5701
rect 12140 -5599 12174 -5565
rect 12140 -5667 12174 -5633
rect 12140 -5735 12174 -5701
rect 12334 -5599 12368 -5565
rect 12334 -5667 12368 -5633
rect 12334 -5735 12368 -5701
rect 12592 -5599 12626 -5565
rect 12592 -5667 12626 -5633
rect 12592 -5735 12626 -5701
rect 12850 -5599 12884 -5565
rect 12850 -5667 12884 -5633
rect 12850 -5735 12884 -5701
rect 13108 -5599 13142 -5565
rect 13108 -5667 13142 -5633
rect 13108 -5735 13142 -5701
rect 13366 -5599 13400 -5565
rect 13366 -5667 13400 -5633
rect 13366 -5735 13400 -5701
rect 13560 -5599 13594 -5565
rect 13560 -5667 13594 -5633
rect 13560 -5735 13594 -5701
rect 13818 -5599 13852 -5565
rect 13818 -5667 13852 -5633
rect 13818 -5735 13852 -5701
rect 14046 -5599 14080 -5565
rect 14046 -5667 14080 -5633
rect 14046 -5735 14080 -5701
rect 14304 -5599 14338 -5565
rect 14304 -5667 14338 -5633
rect 14304 -5735 14338 -5701
rect 14497 -5599 14531 -5565
rect 14497 -5667 14531 -5633
rect 14497 -5735 14531 -5701
rect 14755 -5599 14789 -5565
rect 14755 -5667 14789 -5633
rect 14755 -5735 14789 -5701
rect 15013 -5599 15047 -5565
rect 15013 -5667 15047 -5633
rect 15013 -5735 15047 -5701
rect 15271 -5599 15305 -5565
rect 15271 -5667 15305 -5633
rect 15271 -5735 15305 -5701
rect 15529 -5599 15563 -5565
rect 15529 -5667 15563 -5633
rect 15529 -5735 15563 -5701
rect 15723 -5599 15757 -5565
rect 15723 -5667 15757 -5633
rect 15723 -5735 15757 -5701
rect 15981 -5599 16015 -5565
rect 15981 -5667 16015 -5633
rect 15981 -5735 16015 -5701
rect 16239 -5599 16273 -5565
rect 16239 -5667 16273 -5633
rect 16239 -5735 16273 -5701
rect 16497 -5599 16531 -5565
rect 16497 -5667 16531 -5633
rect 16497 -5735 16531 -5701
rect 16691 -5599 16725 -5565
rect 16691 -5667 16725 -5633
rect 16691 -5735 16725 -5701
rect 16949 -5599 16983 -5565
rect 16949 -5667 16983 -5633
rect 16949 -5735 16983 -5701
rect 17207 -5599 17241 -5565
rect 17207 -5667 17241 -5633
rect 17207 -5735 17241 -5701
rect 17465 -5599 17499 -5565
rect 17465 -5667 17499 -5633
rect 17465 -5735 17499 -5701
rect 17723 -5599 17757 -5565
rect 17723 -5667 17757 -5633
rect 17723 -5735 17757 -5701
rect 17917 -5599 17951 -5565
rect 17917 -5667 17951 -5633
rect 17917 -5735 17951 -5701
rect 18175 -5599 18209 -5565
rect 18175 -5667 18209 -5633
rect 18175 -5735 18209 -5701
rect 971 -6289 1005 -6255
rect 971 -6357 1005 -6323
rect 971 -6425 1005 -6391
rect 1229 -6289 1263 -6255
rect 1229 -6357 1263 -6323
rect 1229 -6425 1263 -6391
rect 1423 -6289 1457 -6255
rect 1423 -6357 1457 -6323
rect 1423 -6425 1457 -6391
rect 1681 -6289 1715 -6255
rect 1681 -6357 1715 -6323
rect 1681 -6425 1715 -6391
rect 1939 -6289 1973 -6255
rect 1939 -6357 1973 -6323
rect 1939 -6425 1973 -6391
rect 2197 -6289 2231 -6255
rect 2197 -6357 2231 -6323
rect 2197 -6425 2231 -6391
rect 2455 -6289 2489 -6255
rect 2455 -6357 2489 -6323
rect 2455 -6425 2489 -6391
rect 2649 -6289 2683 -6255
rect 2649 -6357 2683 -6323
rect 2649 -6425 2683 -6391
rect 2907 -6289 2941 -6255
rect 2907 -6357 2941 -6323
rect 2907 -6425 2941 -6391
rect 3165 -6289 3199 -6255
rect 3165 -6357 3199 -6323
rect 3165 -6425 3199 -6391
rect 3423 -6289 3457 -6255
rect 3423 -6357 3457 -6323
rect 3423 -6425 3457 -6391
rect 3617 -6289 3651 -6255
rect 3617 -6357 3651 -6323
rect 3617 -6425 3651 -6391
rect 3875 -6289 3909 -6255
rect 3875 -6357 3909 -6323
rect 3875 -6425 3909 -6391
rect 4133 -6289 4167 -6255
rect 4133 -6357 4167 -6323
rect 4133 -6425 4167 -6391
rect 4391 -6289 4425 -6255
rect 4391 -6357 4425 -6323
rect 4391 -6425 4425 -6391
rect 4649 -6289 4683 -6255
rect 4649 -6357 4683 -6323
rect 4649 -6425 4683 -6391
rect 4842 -6289 4876 -6255
rect 4842 -6357 4876 -6323
rect 4842 -6425 4876 -6391
rect 5100 -6289 5134 -6255
rect 5100 -6357 5134 -6323
rect 5100 -6425 5134 -6391
rect 5328 -6289 5362 -6255
rect 5328 -6357 5362 -6323
rect 5328 -6425 5362 -6391
rect 5586 -6289 5620 -6255
rect 5586 -6357 5620 -6323
rect 5586 -6425 5620 -6391
rect 5780 -6289 5814 -6255
rect 5780 -6357 5814 -6323
rect 5780 -6425 5814 -6391
rect 6038 -6289 6072 -6255
rect 6038 -6357 6072 -6323
rect 6038 -6425 6072 -6391
rect 6296 -6289 6330 -6255
rect 6296 -6357 6330 -6323
rect 6296 -6425 6330 -6391
rect 6554 -6289 6588 -6255
rect 6554 -6357 6588 -6323
rect 6554 -6425 6588 -6391
rect 6812 -6289 6846 -6255
rect 6812 -6357 6846 -6323
rect 6812 -6425 6846 -6391
rect 7006 -6289 7040 -6255
rect 7006 -6357 7040 -6323
rect 7006 -6425 7040 -6391
rect 7264 -6289 7298 -6255
rect 7264 -6357 7298 -6323
rect 7264 -6425 7298 -6391
rect 7522 -6289 7556 -6255
rect 7522 -6357 7556 -6323
rect 7522 -6425 7556 -6391
rect 7780 -6289 7814 -6255
rect 7780 -6357 7814 -6323
rect 7780 -6425 7814 -6391
rect 7974 -6289 8008 -6255
rect 7974 -6357 8008 -6323
rect 7974 -6425 8008 -6391
rect 8232 -6289 8266 -6255
rect 8232 -6357 8266 -6323
rect 8232 -6425 8266 -6391
rect 8490 -6289 8524 -6255
rect 8490 -6357 8524 -6323
rect 8490 -6425 8524 -6391
rect 8748 -6289 8782 -6255
rect 8748 -6357 8782 -6323
rect 8748 -6425 8782 -6391
rect 9006 -6289 9040 -6255
rect 9006 -6357 9040 -6323
rect 9006 -6425 9040 -6391
rect 9200 -6289 9234 -6255
rect 9200 -6357 9234 -6323
rect 9200 -6425 9234 -6391
rect 9458 -6289 9492 -6255
rect 9458 -6357 9492 -6323
rect 9458 -6425 9492 -6391
rect 9688 -6289 9722 -6255
rect 9688 -6357 9722 -6323
rect 9688 -6425 9722 -6391
rect 9946 -6289 9980 -6255
rect 9946 -6357 9980 -6323
rect 9946 -6425 9980 -6391
rect 10140 -6289 10174 -6255
rect 10140 -6357 10174 -6323
rect 10140 -6425 10174 -6391
rect 10398 -6289 10432 -6255
rect 10398 -6357 10432 -6323
rect 10398 -6425 10432 -6391
rect 10656 -6289 10690 -6255
rect 10656 -6357 10690 -6323
rect 10656 -6425 10690 -6391
rect 10914 -6289 10948 -6255
rect 10914 -6357 10948 -6323
rect 10914 -6425 10948 -6391
rect 11172 -6289 11206 -6255
rect 11172 -6357 11206 -6323
rect 11172 -6425 11206 -6391
rect 11366 -6289 11400 -6255
rect 11366 -6357 11400 -6323
rect 11366 -6425 11400 -6391
rect 11624 -6289 11658 -6255
rect 11624 -6357 11658 -6323
rect 11624 -6425 11658 -6391
rect 11882 -6289 11916 -6255
rect 11882 -6357 11916 -6323
rect 11882 -6425 11916 -6391
rect 12140 -6289 12174 -6255
rect 12140 -6357 12174 -6323
rect 12140 -6425 12174 -6391
rect 12334 -6289 12368 -6255
rect 12334 -6357 12368 -6323
rect 12334 -6425 12368 -6391
rect 12592 -6289 12626 -6255
rect 12592 -6357 12626 -6323
rect 12592 -6425 12626 -6391
rect 12850 -6289 12884 -6255
rect 12850 -6357 12884 -6323
rect 12850 -6425 12884 -6391
rect 13108 -6289 13142 -6255
rect 13108 -6357 13142 -6323
rect 13108 -6425 13142 -6391
rect 13366 -6289 13400 -6255
rect 13366 -6357 13400 -6323
rect 13366 -6425 13400 -6391
rect 13560 -6289 13594 -6255
rect 13560 -6357 13594 -6323
rect 13560 -6425 13594 -6391
rect 13818 -6289 13852 -6255
rect 13818 -6357 13852 -6323
rect 13818 -6425 13852 -6391
rect 14046 -6289 14080 -6255
rect 14046 -6357 14080 -6323
rect 14046 -6425 14080 -6391
rect 14304 -6289 14338 -6255
rect 14304 -6357 14338 -6323
rect 14304 -6425 14338 -6391
rect 14497 -6289 14531 -6255
rect 14497 -6357 14531 -6323
rect 14497 -6425 14531 -6391
rect 14755 -6289 14789 -6255
rect 14755 -6357 14789 -6323
rect 14755 -6425 14789 -6391
rect 15013 -6289 15047 -6255
rect 15013 -6357 15047 -6323
rect 15013 -6425 15047 -6391
rect 15271 -6289 15305 -6255
rect 15271 -6357 15305 -6323
rect 15271 -6425 15305 -6391
rect 15529 -6289 15563 -6255
rect 15529 -6357 15563 -6323
rect 15529 -6425 15563 -6391
rect 15723 -6289 15757 -6255
rect 15723 -6357 15757 -6323
rect 15723 -6425 15757 -6391
rect 15981 -6289 16015 -6255
rect 15981 -6357 16015 -6323
rect 15981 -6425 16015 -6391
rect 16239 -6289 16273 -6255
rect 16239 -6357 16273 -6323
rect 16239 -6425 16273 -6391
rect 16497 -6289 16531 -6255
rect 16497 -6357 16531 -6323
rect 16497 -6425 16531 -6391
rect 16691 -6289 16725 -6255
rect 16691 -6357 16725 -6323
rect 16691 -6425 16725 -6391
rect 16949 -6289 16983 -6255
rect 16949 -6357 16983 -6323
rect 16949 -6425 16983 -6391
rect 17207 -6289 17241 -6255
rect 17207 -6357 17241 -6323
rect 17207 -6425 17241 -6391
rect 17465 -6289 17499 -6255
rect 17465 -6357 17499 -6323
rect 17465 -6425 17499 -6391
rect 17723 -6289 17757 -6255
rect 17723 -6357 17757 -6323
rect 17723 -6425 17757 -6391
rect 17917 -6289 17951 -6255
rect 17917 -6357 17951 -6323
rect 17917 -6425 17951 -6391
rect 18175 -6289 18209 -6255
rect 18175 -6357 18209 -6323
rect 18175 -6425 18209 -6391
rect 971 -7246 1005 -7212
rect 971 -7314 1005 -7280
rect 971 -7382 1005 -7348
rect 1229 -7246 1263 -7212
rect 1229 -7314 1263 -7280
rect 1229 -7382 1263 -7348
rect 1423 -7246 1457 -7212
rect 1423 -7314 1457 -7280
rect 1423 -7382 1457 -7348
rect 1681 -7246 1715 -7212
rect 1681 -7314 1715 -7280
rect 1681 -7382 1715 -7348
rect 1939 -7246 1973 -7212
rect 1939 -7314 1973 -7280
rect 1939 -7382 1973 -7348
rect 2197 -7246 2231 -7212
rect 2197 -7314 2231 -7280
rect 2197 -7382 2231 -7348
rect 2455 -7246 2489 -7212
rect 2455 -7314 2489 -7280
rect 2455 -7382 2489 -7348
rect 2649 -7246 2683 -7212
rect 2649 -7314 2683 -7280
rect 2649 -7382 2683 -7348
rect 2907 -7246 2941 -7212
rect 2907 -7314 2941 -7280
rect 2907 -7382 2941 -7348
rect 3165 -7246 3199 -7212
rect 3165 -7314 3199 -7280
rect 3165 -7382 3199 -7348
rect 3423 -7246 3457 -7212
rect 3423 -7314 3457 -7280
rect 3423 -7382 3457 -7348
rect 3617 -7246 3651 -7212
rect 3617 -7314 3651 -7280
rect 3617 -7382 3651 -7348
rect 3875 -7246 3909 -7212
rect 3875 -7314 3909 -7280
rect 3875 -7382 3909 -7348
rect 4133 -7246 4167 -7212
rect 4133 -7314 4167 -7280
rect 4133 -7382 4167 -7348
rect 4391 -7246 4425 -7212
rect 4391 -7314 4425 -7280
rect 4391 -7382 4425 -7348
rect 4649 -7246 4683 -7212
rect 4649 -7314 4683 -7280
rect 4649 -7382 4683 -7348
rect 4842 -7246 4876 -7212
rect 4842 -7314 4876 -7280
rect 4842 -7382 4876 -7348
rect 5100 -7246 5134 -7212
rect 5100 -7314 5134 -7280
rect 5100 -7382 5134 -7348
rect 5328 -7246 5362 -7212
rect 5328 -7314 5362 -7280
rect 5328 -7382 5362 -7348
rect 5586 -7246 5620 -7212
rect 5586 -7314 5620 -7280
rect 5586 -7382 5620 -7348
rect 5780 -7246 5814 -7212
rect 5780 -7314 5814 -7280
rect 5780 -7382 5814 -7348
rect 6038 -7246 6072 -7212
rect 6038 -7314 6072 -7280
rect 6038 -7382 6072 -7348
rect 6296 -7246 6330 -7212
rect 6296 -7314 6330 -7280
rect 6296 -7382 6330 -7348
rect 6554 -7246 6588 -7212
rect 6554 -7314 6588 -7280
rect 6554 -7382 6588 -7348
rect 6812 -7246 6846 -7212
rect 6812 -7314 6846 -7280
rect 6812 -7382 6846 -7348
rect 7006 -7246 7040 -7212
rect 7006 -7314 7040 -7280
rect 7006 -7382 7040 -7348
rect 7264 -7246 7298 -7212
rect 7264 -7314 7298 -7280
rect 7264 -7382 7298 -7348
rect 7522 -7246 7556 -7212
rect 7522 -7314 7556 -7280
rect 7522 -7382 7556 -7348
rect 7780 -7246 7814 -7212
rect 7780 -7314 7814 -7280
rect 7780 -7382 7814 -7348
rect 7974 -7246 8008 -7212
rect 7974 -7314 8008 -7280
rect 7974 -7382 8008 -7348
rect 8232 -7246 8266 -7212
rect 8232 -7314 8266 -7280
rect 8232 -7382 8266 -7348
rect 8490 -7246 8524 -7212
rect 8490 -7314 8524 -7280
rect 8490 -7382 8524 -7348
rect 8748 -7246 8782 -7212
rect 8748 -7314 8782 -7280
rect 8748 -7382 8782 -7348
rect 9006 -7246 9040 -7212
rect 9006 -7314 9040 -7280
rect 9006 -7382 9040 -7348
rect 9200 -7246 9234 -7212
rect 9200 -7314 9234 -7280
rect 9200 -7382 9234 -7348
rect 9458 -7246 9492 -7212
rect 9458 -7314 9492 -7280
rect 9458 -7382 9492 -7348
rect 9688 -7246 9722 -7212
rect 9688 -7314 9722 -7280
rect 9688 -7382 9722 -7348
rect 9946 -7246 9980 -7212
rect 9946 -7314 9980 -7280
rect 9946 -7382 9980 -7348
rect 10140 -7246 10174 -7212
rect 10140 -7314 10174 -7280
rect 10140 -7382 10174 -7348
rect 10398 -7246 10432 -7212
rect 10398 -7314 10432 -7280
rect 10398 -7382 10432 -7348
rect 10656 -7246 10690 -7212
rect 10656 -7314 10690 -7280
rect 10656 -7382 10690 -7348
rect 10914 -7246 10948 -7212
rect 10914 -7314 10948 -7280
rect 10914 -7382 10948 -7348
rect 11172 -7246 11206 -7212
rect 11172 -7314 11206 -7280
rect 11172 -7382 11206 -7348
rect 11366 -7246 11400 -7212
rect 11366 -7314 11400 -7280
rect 11366 -7382 11400 -7348
rect 11624 -7246 11658 -7212
rect 11624 -7314 11658 -7280
rect 11624 -7382 11658 -7348
rect 11882 -7246 11916 -7212
rect 11882 -7314 11916 -7280
rect 11882 -7382 11916 -7348
rect 12140 -7246 12174 -7212
rect 12140 -7314 12174 -7280
rect 12140 -7382 12174 -7348
rect 12334 -7246 12368 -7212
rect 12334 -7314 12368 -7280
rect 12334 -7382 12368 -7348
rect 12592 -7246 12626 -7212
rect 12592 -7314 12626 -7280
rect 12592 -7382 12626 -7348
rect 12850 -7246 12884 -7212
rect 12850 -7314 12884 -7280
rect 12850 -7382 12884 -7348
rect 13108 -7246 13142 -7212
rect 13108 -7314 13142 -7280
rect 13108 -7382 13142 -7348
rect 13366 -7246 13400 -7212
rect 13366 -7314 13400 -7280
rect 13366 -7382 13400 -7348
rect 13560 -7246 13594 -7212
rect 13560 -7314 13594 -7280
rect 13560 -7382 13594 -7348
rect 13818 -7246 13852 -7212
rect 13818 -7314 13852 -7280
rect 13818 -7382 13852 -7348
rect 14046 -7246 14080 -7212
rect 14046 -7314 14080 -7280
rect 14046 -7382 14080 -7348
rect 14304 -7246 14338 -7212
rect 14304 -7314 14338 -7280
rect 14304 -7382 14338 -7348
rect 14497 -7246 14531 -7212
rect 14497 -7314 14531 -7280
rect 14497 -7382 14531 -7348
rect 14755 -7246 14789 -7212
rect 14755 -7314 14789 -7280
rect 14755 -7382 14789 -7348
rect 15013 -7246 15047 -7212
rect 15013 -7314 15047 -7280
rect 15013 -7382 15047 -7348
rect 15271 -7246 15305 -7212
rect 15271 -7314 15305 -7280
rect 15271 -7382 15305 -7348
rect 15529 -7246 15563 -7212
rect 15529 -7314 15563 -7280
rect 15529 -7382 15563 -7348
rect 15723 -7246 15757 -7212
rect 15723 -7314 15757 -7280
rect 15723 -7382 15757 -7348
rect 15981 -7246 16015 -7212
rect 15981 -7314 16015 -7280
rect 15981 -7382 16015 -7348
rect 16239 -7246 16273 -7212
rect 16239 -7314 16273 -7280
rect 16239 -7382 16273 -7348
rect 16497 -7246 16531 -7212
rect 16497 -7314 16531 -7280
rect 16497 -7382 16531 -7348
rect 16691 -7246 16725 -7212
rect 16691 -7314 16725 -7280
rect 16691 -7382 16725 -7348
rect 16949 -7246 16983 -7212
rect 16949 -7314 16983 -7280
rect 16949 -7382 16983 -7348
rect 17207 -7246 17241 -7212
rect 17207 -7314 17241 -7280
rect 17207 -7382 17241 -7348
rect 17465 -7246 17499 -7212
rect 17465 -7314 17499 -7280
rect 17465 -7382 17499 -7348
rect 17723 -7246 17757 -7212
rect 17723 -7314 17757 -7280
rect 17723 -7382 17757 -7348
rect 17917 -7246 17951 -7212
rect 17917 -7314 17951 -7280
rect 17917 -7382 17951 -7348
rect 18175 -7246 18209 -7212
rect 18175 -7314 18209 -7280
rect 18175 -7382 18209 -7348
rect 971 -7936 1005 -7902
rect 971 -8004 1005 -7970
rect 971 -8072 1005 -8038
rect 1229 -7936 1263 -7902
rect 1229 -8004 1263 -7970
rect 1229 -8072 1263 -8038
rect 1423 -7936 1457 -7902
rect 1423 -8004 1457 -7970
rect 1423 -8072 1457 -8038
rect 1681 -7936 1715 -7902
rect 1681 -8004 1715 -7970
rect 1681 -8072 1715 -8038
rect 1939 -7936 1973 -7902
rect 1939 -8004 1973 -7970
rect 1939 -8072 1973 -8038
rect 2197 -7936 2231 -7902
rect 2197 -8004 2231 -7970
rect 2197 -8072 2231 -8038
rect 2455 -7936 2489 -7902
rect 2455 -8004 2489 -7970
rect 2455 -8072 2489 -8038
rect 2649 -7936 2683 -7902
rect 2649 -8004 2683 -7970
rect 2649 -8072 2683 -8038
rect 2907 -7936 2941 -7902
rect 2907 -8004 2941 -7970
rect 2907 -8072 2941 -8038
rect 3165 -7936 3199 -7902
rect 3165 -8004 3199 -7970
rect 3165 -8072 3199 -8038
rect 3423 -7936 3457 -7902
rect 3423 -8004 3457 -7970
rect 3423 -8072 3457 -8038
rect 3617 -7936 3651 -7902
rect 3617 -8004 3651 -7970
rect 3617 -8072 3651 -8038
rect 3875 -7936 3909 -7902
rect 3875 -8004 3909 -7970
rect 3875 -8072 3909 -8038
rect 4133 -7936 4167 -7902
rect 4133 -8004 4167 -7970
rect 4133 -8072 4167 -8038
rect 4391 -7936 4425 -7902
rect 4391 -8004 4425 -7970
rect 4391 -8072 4425 -8038
rect 4649 -7936 4683 -7902
rect 4649 -8004 4683 -7970
rect 4649 -8072 4683 -8038
rect 4842 -7936 4876 -7902
rect 4842 -8004 4876 -7970
rect 4842 -8072 4876 -8038
rect 5100 -7936 5134 -7902
rect 5100 -8004 5134 -7970
rect 5100 -8072 5134 -8038
rect 5328 -7936 5362 -7902
rect 5328 -8004 5362 -7970
rect 5328 -8072 5362 -8038
rect 5586 -7936 5620 -7902
rect 5586 -8004 5620 -7970
rect 5586 -8072 5620 -8038
rect 5780 -7936 5814 -7902
rect 5780 -8004 5814 -7970
rect 5780 -8072 5814 -8038
rect 6038 -7936 6072 -7902
rect 6038 -8004 6072 -7970
rect 6038 -8072 6072 -8038
rect 6296 -7936 6330 -7902
rect 6296 -8004 6330 -7970
rect 6296 -8072 6330 -8038
rect 6554 -7936 6588 -7902
rect 6554 -8004 6588 -7970
rect 6554 -8072 6588 -8038
rect 6812 -7936 6846 -7902
rect 6812 -8004 6846 -7970
rect 6812 -8072 6846 -8038
rect 7006 -7936 7040 -7902
rect 7006 -8004 7040 -7970
rect 7006 -8072 7040 -8038
rect 7264 -7936 7298 -7902
rect 7264 -8004 7298 -7970
rect 7264 -8072 7298 -8038
rect 7522 -7936 7556 -7902
rect 7522 -8004 7556 -7970
rect 7522 -8072 7556 -8038
rect 7780 -7936 7814 -7902
rect 7780 -8004 7814 -7970
rect 7780 -8072 7814 -8038
rect 7974 -7936 8008 -7902
rect 7974 -8004 8008 -7970
rect 7974 -8072 8008 -8038
rect 8232 -7936 8266 -7902
rect 8232 -8004 8266 -7970
rect 8232 -8072 8266 -8038
rect 8490 -7936 8524 -7902
rect 8490 -8004 8524 -7970
rect 8490 -8072 8524 -8038
rect 8748 -7936 8782 -7902
rect 8748 -8004 8782 -7970
rect 8748 -8072 8782 -8038
rect 9006 -7936 9040 -7902
rect 9006 -8004 9040 -7970
rect 9006 -8072 9040 -8038
rect 9200 -7936 9234 -7902
rect 9200 -8004 9234 -7970
rect 9200 -8072 9234 -8038
rect 9458 -7936 9492 -7902
rect 9458 -8004 9492 -7970
rect 9458 -8072 9492 -8038
rect 9688 -7936 9722 -7902
rect 9688 -8004 9722 -7970
rect 9688 -8072 9722 -8038
rect 9946 -7936 9980 -7902
rect 9946 -8004 9980 -7970
rect 9946 -8072 9980 -8038
rect 10140 -7936 10174 -7902
rect 10140 -8004 10174 -7970
rect 10140 -8072 10174 -8038
rect 10398 -7936 10432 -7902
rect 10398 -8004 10432 -7970
rect 10398 -8072 10432 -8038
rect 10656 -7936 10690 -7902
rect 10656 -8004 10690 -7970
rect 10656 -8072 10690 -8038
rect 10914 -7936 10948 -7902
rect 10914 -8004 10948 -7970
rect 10914 -8072 10948 -8038
rect 11172 -7936 11206 -7902
rect 11172 -8004 11206 -7970
rect 11172 -8072 11206 -8038
rect 11366 -7936 11400 -7902
rect 11366 -8004 11400 -7970
rect 11366 -8072 11400 -8038
rect 11624 -7936 11658 -7902
rect 11624 -8004 11658 -7970
rect 11624 -8072 11658 -8038
rect 11882 -7936 11916 -7902
rect 11882 -8004 11916 -7970
rect 11882 -8072 11916 -8038
rect 12140 -7936 12174 -7902
rect 12140 -8004 12174 -7970
rect 12140 -8072 12174 -8038
rect 12334 -7936 12368 -7902
rect 12334 -8004 12368 -7970
rect 12334 -8072 12368 -8038
rect 12592 -7936 12626 -7902
rect 12592 -8004 12626 -7970
rect 12592 -8072 12626 -8038
rect 12850 -7936 12884 -7902
rect 12850 -8004 12884 -7970
rect 12850 -8072 12884 -8038
rect 13108 -7936 13142 -7902
rect 13108 -8004 13142 -7970
rect 13108 -8072 13142 -8038
rect 13366 -7936 13400 -7902
rect 13366 -8004 13400 -7970
rect 13366 -8072 13400 -8038
rect 13560 -7936 13594 -7902
rect 13560 -8004 13594 -7970
rect 13560 -8072 13594 -8038
rect 13818 -7936 13852 -7902
rect 13818 -8004 13852 -7970
rect 13818 -8072 13852 -8038
rect 14046 -7936 14080 -7902
rect 14046 -8004 14080 -7970
rect 14046 -8072 14080 -8038
rect 14304 -7936 14338 -7902
rect 14304 -8004 14338 -7970
rect 14304 -8072 14338 -8038
rect 14497 -7936 14531 -7902
rect 14497 -8004 14531 -7970
rect 14497 -8072 14531 -8038
rect 14755 -7936 14789 -7902
rect 14755 -8004 14789 -7970
rect 14755 -8072 14789 -8038
rect 15013 -7936 15047 -7902
rect 15013 -8004 15047 -7970
rect 15013 -8072 15047 -8038
rect 15271 -7936 15305 -7902
rect 15271 -8004 15305 -7970
rect 15271 -8072 15305 -8038
rect 15529 -7936 15563 -7902
rect 15529 -8004 15563 -7970
rect 15529 -8072 15563 -8038
rect 15723 -7936 15757 -7902
rect 15723 -8004 15757 -7970
rect 15723 -8072 15757 -8038
rect 15981 -7936 16015 -7902
rect 15981 -8004 16015 -7970
rect 15981 -8072 16015 -8038
rect 16239 -7936 16273 -7902
rect 16239 -8004 16273 -7970
rect 16239 -8072 16273 -8038
rect 16497 -7936 16531 -7902
rect 16497 -8004 16531 -7970
rect 16497 -8072 16531 -8038
rect 16691 -7936 16725 -7902
rect 16691 -8004 16725 -7970
rect 16691 -8072 16725 -8038
rect 16949 -7936 16983 -7902
rect 16949 -8004 16983 -7970
rect 16949 -8072 16983 -8038
rect 17207 -7936 17241 -7902
rect 17207 -8004 17241 -7970
rect 17207 -8072 17241 -8038
rect 17465 -7936 17499 -7902
rect 17465 -8004 17499 -7970
rect 17465 -8072 17499 -8038
rect 17723 -7936 17757 -7902
rect 17723 -8004 17757 -7970
rect 17723 -8072 17757 -8038
rect 17917 -7936 17951 -7902
rect 17917 -8004 17951 -7970
rect 17917 -8072 17951 -8038
rect 18175 -7936 18209 -7902
rect 18175 -8004 18209 -7970
rect 18175 -8072 18209 -8038
rect 971 -8880 1005 -8846
rect 971 -8948 1005 -8914
rect 971 -9016 1005 -8982
rect 1229 -8880 1263 -8846
rect 1229 -8948 1263 -8914
rect 1229 -9016 1263 -8982
rect 1423 -8880 1457 -8846
rect 1423 -8948 1457 -8914
rect 1423 -9016 1457 -8982
rect 1681 -8880 1715 -8846
rect 1681 -8948 1715 -8914
rect 1681 -9016 1715 -8982
rect 1939 -8880 1973 -8846
rect 1939 -8948 1973 -8914
rect 1939 -9016 1973 -8982
rect 2197 -8880 2231 -8846
rect 2197 -8948 2231 -8914
rect 2197 -9016 2231 -8982
rect 2455 -8880 2489 -8846
rect 2455 -8948 2489 -8914
rect 2455 -9016 2489 -8982
rect 2649 -8880 2683 -8846
rect 2649 -8948 2683 -8914
rect 2649 -9016 2683 -8982
rect 2907 -8880 2941 -8846
rect 2907 -8948 2941 -8914
rect 2907 -9016 2941 -8982
rect 3165 -8880 3199 -8846
rect 3165 -8948 3199 -8914
rect 3165 -9016 3199 -8982
rect 3423 -8880 3457 -8846
rect 3423 -8948 3457 -8914
rect 3423 -9016 3457 -8982
rect 3617 -8880 3651 -8846
rect 3617 -8948 3651 -8914
rect 3617 -9016 3651 -8982
rect 3875 -8880 3909 -8846
rect 3875 -8948 3909 -8914
rect 3875 -9016 3909 -8982
rect 4133 -8880 4167 -8846
rect 4133 -8948 4167 -8914
rect 4133 -9016 4167 -8982
rect 4391 -8880 4425 -8846
rect 4391 -8948 4425 -8914
rect 4391 -9016 4425 -8982
rect 4649 -8880 4683 -8846
rect 4649 -8948 4683 -8914
rect 4649 -9016 4683 -8982
rect 4842 -8880 4876 -8846
rect 4842 -8948 4876 -8914
rect 4842 -9016 4876 -8982
rect 5100 -8880 5134 -8846
rect 5100 -8948 5134 -8914
rect 5100 -9016 5134 -8982
rect 5328 -8880 5362 -8846
rect 5328 -8948 5362 -8914
rect 5328 -9016 5362 -8982
rect 5586 -8880 5620 -8846
rect 5586 -8948 5620 -8914
rect 5586 -9016 5620 -8982
rect 5780 -8880 5814 -8846
rect 5780 -8948 5814 -8914
rect 5780 -9016 5814 -8982
rect 6038 -8880 6072 -8846
rect 6038 -8948 6072 -8914
rect 6038 -9016 6072 -8982
rect 6296 -8880 6330 -8846
rect 6296 -8948 6330 -8914
rect 6296 -9016 6330 -8982
rect 6554 -8880 6588 -8846
rect 6554 -8948 6588 -8914
rect 6554 -9016 6588 -8982
rect 6812 -8880 6846 -8846
rect 6812 -8948 6846 -8914
rect 6812 -9016 6846 -8982
rect 7006 -8880 7040 -8846
rect 7006 -8948 7040 -8914
rect 7006 -9016 7040 -8982
rect 7264 -8880 7298 -8846
rect 7264 -8948 7298 -8914
rect 7264 -9016 7298 -8982
rect 7522 -8880 7556 -8846
rect 7522 -8948 7556 -8914
rect 7522 -9016 7556 -8982
rect 7780 -8880 7814 -8846
rect 7780 -8948 7814 -8914
rect 7780 -9016 7814 -8982
rect 7974 -8880 8008 -8846
rect 7974 -8948 8008 -8914
rect 7974 -9016 8008 -8982
rect 8232 -8880 8266 -8846
rect 8232 -8948 8266 -8914
rect 8232 -9016 8266 -8982
rect 8490 -8880 8524 -8846
rect 8490 -8948 8524 -8914
rect 8490 -9016 8524 -8982
rect 8748 -8880 8782 -8846
rect 8748 -8948 8782 -8914
rect 8748 -9016 8782 -8982
rect 9006 -8880 9040 -8846
rect 9006 -8948 9040 -8914
rect 9006 -9016 9040 -8982
rect 9200 -8880 9234 -8846
rect 9200 -8948 9234 -8914
rect 9200 -9016 9234 -8982
rect 9458 -8880 9492 -8846
rect 9458 -8948 9492 -8914
rect 9458 -9016 9492 -8982
rect 9688 -8880 9722 -8846
rect 9688 -8948 9722 -8914
rect 9688 -9016 9722 -8982
rect 9946 -8880 9980 -8846
rect 9946 -8948 9980 -8914
rect 9946 -9016 9980 -8982
rect 10140 -8880 10174 -8846
rect 10140 -8948 10174 -8914
rect 10140 -9016 10174 -8982
rect 10398 -8880 10432 -8846
rect 10398 -8948 10432 -8914
rect 10398 -9016 10432 -8982
rect 10656 -8880 10690 -8846
rect 10656 -8948 10690 -8914
rect 10656 -9016 10690 -8982
rect 10914 -8880 10948 -8846
rect 10914 -8948 10948 -8914
rect 10914 -9016 10948 -8982
rect 11172 -8880 11206 -8846
rect 11172 -8948 11206 -8914
rect 11172 -9016 11206 -8982
rect 11366 -8880 11400 -8846
rect 11366 -8948 11400 -8914
rect 11366 -9016 11400 -8982
rect 11624 -8880 11658 -8846
rect 11624 -8948 11658 -8914
rect 11624 -9016 11658 -8982
rect 11882 -8880 11916 -8846
rect 11882 -8948 11916 -8914
rect 11882 -9016 11916 -8982
rect 12140 -8880 12174 -8846
rect 12140 -8948 12174 -8914
rect 12140 -9016 12174 -8982
rect 12334 -8880 12368 -8846
rect 12334 -8948 12368 -8914
rect 12334 -9016 12368 -8982
rect 12592 -8880 12626 -8846
rect 12592 -8948 12626 -8914
rect 12592 -9016 12626 -8982
rect 12850 -8880 12884 -8846
rect 12850 -8948 12884 -8914
rect 12850 -9016 12884 -8982
rect 13108 -8880 13142 -8846
rect 13108 -8948 13142 -8914
rect 13108 -9016 13142 -8982
rect 13366 -8880 13400 -8846
rect 13366 -8948 13400 -8914
rect 13366 -9016 13400 -8982
rect 13560 -8880 13594 -8846
rect 13560 -8948 13594 -8914
rect 13560 -9016 13594 -8982
rect 13818 -8880 13852 -8846
rect 13818 -8948 13852 -8914
rect 13818 -9016 13852 -8982
rect 14046 -8880 14080 -8846
rect 14046 -8948 14080 -8914
rect 14046 -9016 14080 -8982
rect 14304 -8880 14338 -8846
rect 14304 -8948 14338 -8914
rect 14304 -9016 14338 -8982
rect 14497 -8880 14531 -8846
rect 14497 -8948 14531 -8914
rect 14497 -9016 14531 -8982
rect 14755 -8880 14789 -8846
rect 14755 -8948 14789 -8914
rect 14755 -9016 14789 -8982
rect 15013 -8880 15047 -8846
rect 15013 -8948 15047 -8914
rect 15013 -9016 15047 -8982
rect 15271 -8880 15305 -8846
rect 15271 -8948 15305 -8914
rect 15271 -9016 15305 -8982
rect 15529 -8880 15563 -8846
rect 15529 -8948 15563 -8914
rect 15529 -9016 15563 -8982
rect 15723 -8880 15757 -8846
rect 15723 -8948 15757 -8914
rect 15723 -9016 15757 -8982
rect 15981 -8880 16015 -8846
rect 15981 -8948 16015 -8914
rect 15981 -9016 16015 -8982
rect 16239 -8880 16273 -8846
rect 16239 -8948 16273 -8914
rect 16239 -9016 16273 -8982
rect 16497 -8880 16531 -8846
rect 16497 -8948 16531 -8914
rect 16497 -9016 16531 -8982
rect 16691 -8880 16725 -8846
rect 16691 -8948 16725 -8914
rect 16691 -9016 16725 -8982
rect 16949 -8880 16983 -8846
rect 16949 -8948 16983 -8914
rect 16949 -9016 16983 -8982
rect 17207 -8880 17241 -8846
rect 17207 -8948 17241 -8914
rect 17207 -9016 17241 -8982
rect 17465 -8880 17499 -8846
rect 17465 -8948 17499 -8914
rect 17465 -9016 17499 -8982
rect 17723 -8880 17757 -8846
rect 17723 -8948 17757 -8914
rect 17723 -9016 17757 -8982
rect 17917 -8880 17951 -8846
rect 17917 -8948 17951 -8914
rect 17917 -9016 17951 -8982
rect 18175 -8880 18209 -8846
rect 18175 -8948 18209 -8914
rect 18175 -9016 18209 -8982
<< nsubdiff >>
rect 856 429 977 463
rect 1011 429 1045 463
rect 1079 429 1113 463
rect 1147 429 1181 463
rect 1215 429 1249 463
rect 1283 429 1317 463
rect 1351 429 1385 463
rect 1419 429 1453 463
rect 1487 429 1521 463
rect 1555 429 1589 463
rect 1623 429 1657 463
rect 1691 429 1725 463
rect 1759 429 1793 463
rect 1827 429 1861 463
rect 1895 429 1929 463
rect 1963 429 1997 463
rect 2031 429 2065 463
rect 2099 429 2133 463
rect 2167 429 2201 463
rect 2235 429 2269 463
rect 2303 429 2337 463
rect 2371 429 2405 463
rect 2439 429 2473 463
rect 2507 429 2541 463
rect 2575 429 2609 463
rect 2643 429 2677 463
rect 2711 429 2745 463
rect 2779 429 2813 463
rect 2847 429 2881 463
rect 2915 429 2949 463
rect 2983 429 3017 463
rect 3051 429 3085 463
rect 3119 429 3153 463
rect 3187 429 3221 463
rect 3255 429 3289 463
rect 3323 429 3357 463
rect 3391 429 3425 463
rect 3459 429 3493 463
rect 3527 429 3561 463
rect 3595 429 3629 463
rect 3663 429 3697 463
rect 3731 429 3765 463
rect 3799 429 3833 463
rect 3867 429 3901 463
rect 3935 429 3969 463
rect 4003 429 4037 463
rect 4071 429 4105 463
rect 4139 429 4173 463
rect 4207 429 4241 463
rect 4275 429 4309 463
rect 4343 429 4377 463
rect 4411 429 4445 463
rect 4479 429 4513 463
rect 4547 429 4581 463
rect 4615 429 4649 463
rect 4683 429 4717 463
rect 4751 429 4785 463
rect 4819 429 4853 463
rect 4887 429 4921 463
rect 4955 429 4989 463
rect 5023 429 5057 463
rect 5091 429 5372 463
rect 5406 429 5440 463
rect 5474 429 5508 463
rect 5542 429 5576 463
rect 5610 429 5644 463
rect 5678 429 5712 463
rect 5746 429 5780 463
rect 5814 429 5848 463
rect 5882 429 5916 463
rect 5950 429 5984 463
rect 6018 429 6052 463
rect 6086 429 6120 463
rect 6154 429 6188 463
rect 6222 429 6256 463
rect 6290 429 6324 463
rect 6358 429 6392 463
rect 6426 429 6460 463
rect 6494 429 6528 463
rect 6562 429 6596 463
rect 6630 429 6664 463
rect 6698 429 6732 463
rect 6766 429 6800 463
rect 6834 429 6868 463
rect 6902 429 6936 463
rect 6970 429 7004 463
rect 7038 429 7072 463
rect 7106 429 7140 463
rect 7174 429 7208 463
rect 7242 429 7276 463
rect 7310 429 7344 463
rect 7378 429 7412 463
rect 7446 429 7480 463
rect 7514 429 7548 463
rect 7582 429 7616 463
rect 7650 429 7684 463
rect 7718 429 7752 463
rect 7786 429 7820 463
rect 7854 429 7888 463
rect 7922 429 7956 463
rect 7990 429 8024 463
rect 8058 429 8092 463
rect 8126 429 8160 463
rect 8194 429 8228 463
rect 8262 429 8296 463
rect 8330 429 8364 463
rect 8398 429 8432 463
rect 8466 429 8500 463
rect 8534 429 8568 463
rect 8602 429 8636 463
rect 8670 429 8704 463
rect 8738 429 8772 463
rect 8806 429 8840 463
rect 8874 429 8908 463
rect 8942 429 8976 463
rect 9010 429 9044 463
rect 9078 429 9112 463
rect 9146 429 9180 463
rect 9214 429 9248 463
rect 9282 429 9316 463
rect 9350 429 9384 463
rect 9418 429 9452 463
rect 9486 429 9694 463
rect 9728 429 9762 463
rect 9796 429 9830 463
rect 9864 429 9898 463
rect 9932 429 9966 463
rect 10000 429 10034 463
rect 10068 429 10102 463
rect 10136 429 10170 463
rect 10204 429 10238 463
rect 10272 429 10306 463
rect 10340 429 10374 463
rect 10408 429 10442 463
rect 10476 429 10510 463
rect 10544 429 10578 463
rect 10612 429 10646 463
rect 10680 429 10714 463
rect 10748 429 10782 463
rect 10816 429 10850 463
rect 10884 429 10918 463
rect 10952 429 10986 463
rect 11020 429 11054 463
rect 11088 429 11122 463
rect 11156 429 11190 463
rect 11224 429 11258 463
rect 11292 429 11326 463
rect 11360 429 11394 463
rect 11428 429 11462 463
rect 11496 429 11530 463
rect 11564 429 11598 463
rect 11632 429 11666 463
rect 11700 429 11734 463
rect 11768 429 11802 463
rect 11836 429 11870 463
rect 11904 429 11938 463
rect 11972 429 12006 463
rect 12040 429 12074 463
rect 12108 429 12142 463
rect 12176 429 12210 463
rect 12244 429 12278 463
rect 12312 429 12346 463
rect 12380 429 12414 463
rect 12448 429 12482 463
rect 12516 429 12550 463
rect 12584 429 12618 463
rect 12652 429 12686 463
rect 12720 429 12754 463
rect 12788 429 12822 463
rect 12856 429 12890 463
rect 12924 429 12958 463
rect 12992 429 13026 463
rect 13060 429 13094 463
rect 13128 429 13162 463
rect 13196 429 13230 463
rect 13264 429 13298 463
rect 13332 429 13366 463
rect 13400 429 13434 463
rect 13468 429 13502 463
rect 13536 429 13570 463
rect 13604 429 13638 463
rect 13672 429 13706 463
rect 13740 429 13774 463
rect 13808 429 14089 463
rect 14123 429 14157 463
rect 14191 429 14225 463
rect 14259 429 14293 463
rect 14327 429 14361 463
rect 14395 429 14429 463
rect 14463 429 14497 463
rect 14531 429 14565 463
rect 14599 429 14633 463
rect 14667 429 14701 463
rect 14735 429 14769 463
rect 14803 429 14837 463
rect 14871 429 14905 463
rect 14939 429 14973 463
rect 15007 429 15041 463
rect 15075 429 15109 463
rect 15143 429 15177 463
rect 15211 429 15245 463
rect 15279 429 15313 463
rect 15347 429 15381 463
rect 15415 429 15449 463
rect 15483 429 15517 463
rect 15551 429 15585 463
rect 15619 429 15653 463
rect 15687 429 15721 463
rect 15755 429 15789 463
rect 15823 429 15857 463
rect 15891 429 15925 463
rect 15959 429 15993 463
rect 16027 429 16061 463
rect 16095 429 16129 463
rect 16163 429 16197 463
rect 16231 429 16265 463
rect 16299 429 16333 463
rect 16367 429 16401 463
rect 16435 429 16469 463
rect 16503 429 16537 463
rect 16571 429 16605 463
rect 16639 429 16673 463
rect 16707 429 16741 463
rect 16775 429 16809 463
rect 16843 429 16877 463
rect 16911 429 16945 463
rect 16979 429 17013 463
rect 17047 429 17081 463
rect 17115 429 17149 463
rect 17183 429 17217 463
rect 17251 429 17285 463
rect 17319 429 17353 463
rect 17387 429 17421 463
rect 17455 429 17489 463
rect 17523 429 17557 463
rect 17591 429 17625 463
rect 17659 429 17693 463
rect 17727 429 17761 463
rect 17795 429 17829 463
rect 17863 429 17897 463
rect 17931 429 17965 463
rect 17999 429 18033 463
rect 18067 429 18101 463
rect 18135 429 18169 463
rect 18203 429 18324 463
rect 856 250 890 429
rect 856 182 890 216
rect 856 114 890 148
rect 856 46 890 80
rect 5214 250 5248 429
rect 5214 182 5248 216
rect 5214 114 5248 148
rect 5214 46 5248 80
rect 9573 250 9607 429
rect 9573 182 9607 216
rect 9573 114 9607 148
rect 856 -22 890 12
rect 856 -90 890 -56
rect 856 -158 890 -124
rect 856 -226 890 -192
rect 856 -294 890 -260
rect 9573 46 9607 80
rect 13932 250 13966 429
rect 13932 182 13966 216
rect 13932 114 13966 148
rect 5214 -22 5248 12
rect 5214 -90 5248 -56
rect 5214 -158 5248 -124
rect 5214 -226 5248 -192
rect 5214 -294 5248 -260
rect 13932 46 13966 80
rect 18290 250 18324 429
rect 18290 182 18324 216
rect 18290 114 18324 148
rect 9573 -22 9607 12
rect 9573 -90 9607 -56
rect 9573 -158 9607 -124
rect 9573 -226 9607 -192
rect 9573 -294 9607 -260
rect 18290 46 18324 80
rect 13932 -22 13966 12
rect 13932 -90 13966 -56
rect 13932 -158 13966 -124
rect 13932 -226 13966 -192
rect 13932 -294 13966 -260
rect 18290 -22 18324 12
rect 18290 -90 18324 -56
rect 18290 -158 18324 -124
rect 18290 -226 18324 -192
rect 18290 -294 18324 -260
rect 856 -362 977 -328
rect 1011 -362 1045 -328
rect 1079 -362 1113 -328
rect 1147 -362 1181 -328
rect 1215 -362 1249 -328
rect 1283 -362 1317 -328
rect 1351 -362 1385 -328
rect 1419 -362 1453 -328
rect 1487 -362 1521 -328
rect 1555 -362 1589 -328
rect 1623 -362 1657 -328
rect 1691 -362 1725 -328
rect 1759 -362 1793 -328
rect 1827 -362 1861 -328
rect 1895 -362 1929 -328
rect 1963 -362 1997 -328
rect 2031 -362 2065 -328
rect 2099 -362 2133 -328
rect 2167 -362 2201 -328
rect 2235 -362 2269 -328
rect 2303 -362 2337 -328
rect 2371 -362 2405 -328
rect 2439 -362 2473 -328
rect 2507 -362 2541 -328
rect 2575 -362 2609 -328
rect 2643 -362 2677 -328
rect 2711 -362 2745 -328
rect 2779 -362 2813 -328
rect 2847 -362 2881 -328
rect 2915 -362 2949 -328
rect 2983 -362 3017 -328
rect 3051 -362 3085 -328
rect 3119 -362 3153 -328
rect 3187 -362 3221 -328
rect 3255 -362 3289 -328
rect 3323 -362 3357 -328
rect 3391 -362 3425 -328
rect 3459 -362 3493 -328
rect 3527 -362 3561 -328
rect 3595 -362 3629 -328
rect 3663 -362 3697 -328
rect 3731 -362 3765 -328
rect 3799 -362 3833 -328
rect 3867 -362 3901 -328
rect 3935 -362 3969 -328
rect 4003 -362 4037 -328
rect 4071 -362 4105 -328
rect 4139 -362 4173 -328
rect 4207 -362 4241 -328
rect 4275 -362 4309 -328
rect 4343 -362 4377 -328
rect 4411 -362 4445 -328
rect 4479 -362 4513 -328
rect 4547 -362 4581 -328
rect 4615 -362 4649 -328
rect 4683 -362 4717 -328
rect 4751 -362 4785 -328
rect 4819 -362 4853 -328
rect 4887 -362 4921 -328
rect 4955 -362 4989 -328
rect 5023 -362 5057 -328
rect 5091 -362 5372 -328
rect 5406 -362 5440 -328
rect 5474 -362 5508 -328
rect 5542 -362 5576 -328
rect 5610 -362 5644 -328
rect 5678 -362 5712 -328
rect 5746 -362 5780 -328
rect 5814 -362 5848 -328
rect 5882 -362 5916 -328
rect 5950 -362 5984 -328
rect 6018 -362 6052 -328
rect 6086 -362 6120 -328
rect 6154 -362 6188 -328
rect 6222 -362 6256 -328
rect 6290 -362 6324 -328
rect 6358 -362 6392 -328
rect 6426 -362 6460 -328
rect 6494 -362 6528 -328
rect 6562 -362 6596 -328
rect 6630 -362 6664 -328
rect 6698 -362 6732 -328
rect 6766 -362 6800 -328
rect 6834 -362 6868 -328
rect 6902 -362 6936 -328
rect 6970 -362 7004 -328
rect 7038 -362 7072 -328
rect 7106 -362 7140 -328
rect 7174 -362 7208 -328
rect 7242 -362 7276 -328
rect 7310 -362 7344 -328
rect 7378 -362 7412 -328
rect 7446 -362 7480 -328
rect 7514 -362 7548 -328
rect 7582 -362 7616 -328
rect 7650 -362 7684 -328
rect 7718 -362 7752 -328
rect 7786 -362 7820 -328
rect 7854 -362 7888 -328
rect 7922 -362 7956 -328
rect 7990 -362 8024 -328
rect 8058 -362 8092 -328
rect 8126 -362 8160 -328
rect 8194 -362 8228 -328
rect 8262 -362 8296 -328
rect 8330 -362 8364 -328
rect 8398 -362 8432 -328
rect 8466 -362 8500 -328
rect 8534 -362 8568 -328
rect 8602 -362 8636 -328
rect 8670 -362 8704 -328
rect 8738 -362 8772 -328
rect 8806 -362 8840 -328
rect 8874 -362 8908 -328
rect 8942 -362 8976 -328
rect 9010 -362 9044 -328
rect 9078 -362 9112 -328
rect 9146 -362 9180 -328
rect 9214 -362 9248 -328
rect 9282 -362 9316 -328
rect 9350 -362 9384 -328
rect 9418 -362 9452 -328
rect 9486 -362 9694 -328
rect 9728 -362 9762 -328
rect 9796 -362 9830 -328
rect 9864 -362 9898 -328
rect 9932 -362 9966 -328
rect 10000 -362 10034 -328
rect 10068 -362 10102 -328
rect 10136 -362 10170 -328
rect 10204 -362 10238 -328
rect 10272 -362 10306 -328
rect 10340 -362 10374 -328
rect 10408 -362 10442 -328
rect 10476 -362 10510 -328
rect 10544 -362 10578 -328
rect 10612 -362 10646 -328
rect 10680 -362 10714 -328
rect 10748 -362 10782 -328
rect 10816 -362 10850 -328
rect 10884 -362 10918 -328
rect 10952 -362 10986 -328
rect 11020 -362 11054 -328
rect 11088 -362 11122 -328
rect 11156 -362 11190 -328
rect 11224 -362 11258 -328
rect 11292 -362 11326 -328
rect 11360 -362 11394 -328
rect 11428 -362 11462 -328
rect 11496 -362 11530 -328
rect 11564 -362 11598 -328
rect 11632 -362 11666 -328
rect 11700 -362 11734 -328
rect 11768 -362 11802 -328
rect 11836 -362 11870 -328
rect 11904 -362 11938 -328
rect 11972 -362 12006 -328
rect 12040 -362 12074 -328
rect 12108 -362 12142 -328
rect 12176 -362 12210 -328
rect 12244 -362 12278 -328
rect 12312 -362 12346 -328
rect 12380 -362 12414 -328
rect 12448 -362 12482 -328
rect 12516 -362 12550 -328
rect 12584 -362 12618 -328
rect 12652 -362 12686 -328
rect 12720 -362 12754 -328
rect 12788 -362 12822 -328
rect 12856 -362 12890 -328
rect 12924 -362 12958 -328
rect 12992 -362 13026 -328
rect 13060 -362 13094 -328
rect 13128 -362 13162 -328
rect 13196 -362 13230 -328
rect 13264 -362 13298 -328
rect 13332 -362 13366 -328
rect 13400 -362 13434 -328
rect 13468 -362 13502 -328
rect 13536 -362 13570 -328
rect 13604 -362 13638 -328
rect 13672 -362 13706 -328
rect 13740 -362 13774 -328
rect 13808 -362 14089 -328
rect 14123 -362 14157 -328
rect 14191 -362 14225 -328
rect 14259 -362 14293 -328
rect 14327 -362 14361 -328
rect 14395 -362 14429 -328
rect 14463 -362 14497 -328
rect 14531 -362 14565 -328
rect 14599 -362 14633 -328
rect 14667 -362 14701 -328
rect 14735 -362 14769 -328
rect 14803 -362 14837 -328
rect 14871 -362 14905 -328
rect 14939 -362 14973 -328
rect 15007 -362 15041 -328
rect 15075 -362 15109 -328
rect 15143 -362 15177 -328
rect 15211 -362 15245 -328
rect 15279 -362 15313 -328
rect 15347 -362 15381 -328
rect 15415 -362 15449 -328
rect 15483 -362 15517 -328
rect 15551 -362 15585 -328
rect 15619 -362 15653 -328
rect 15687 -362 15721 -328
rect 15755 -362 15789 -328
rect 15823 -362 15857 -328
rect 15891 -362 15925 -328
rect 15959 -362 15993 -328
rect 16027 -362 16061 -328
rect 16095 -362 16129 -328
rect 16163 -362 16197 -328
rect 16231 -362 16265 -328
rect 16299 -362 16333 -328
rect 16367 -362 16401 -328
rect 16435 -362 16469 -328
rect 16503 -362 16537 -328
rect 16571 -362 16605 -328
rect 16639 -362 16673 -328
rect 16707 -362 16741 -328
rect 16775 -362 16809 -328
rect 16843 -362 16877 -328
rect 16911 -362 16945 -328
rect 16979 -362 17013 -328
rect 17047 -362 17081 -328
rect 17115 -362 17149 -328
rect 17183 -362 17217 -328
rect 17251 -362 17285 -328
rect 17319 -362 17353 -328
rect 17387 -362 17421 -328
rect 17455 -362 17489 -328
rect 17523 -362 17557 -328
rect 17591 -362 17625 -328
rect 17659 -362 17693 -328
rect 17727 -362 17761 -328
rect 17795 -362 17829 -328
rect 17863 -362 17897 -328
rect 17931 -362 17965 -328
rect 17999 -362 18033 -328
rect 18067 -362 18101 -328
rect 18135 -362 18169 -328
rect 18203 -362 18324 -328
rect 856 -430 890 -396
rect 856 -498 890 -464
rect 856 -566 890 -532
rect 856 -634 890 -600
rect 5214 -430 5248 -396
rect 5214 -498 5248 -464
rect 5214 -566 5248 -532
rect 5214 -634 5248 -600
rect 856 -702 890 -668
rect 9573 -430 9607 -396
rect 9573 -498 9607 -464
rect 9573 -566 9607 -532
rect 9573 -634 9607 -600
rect 856 -770 890 -736
rect 856 -838 890 -804
rect 856 -906 890 -872
rect 5214 -702 5248 -668
rect 13932 -430 13966 -396
rect 13932 -498 13966 -464
rect 13932 -566 13966 -532
rect 13932 -634 13966 -600
rect 5214 -770 5248 -736
rect 5214 -838 5248 -804
rect 856 -974 890 -940
rect 5214 -906 5248 -872
rect 9573 -702 9607 -668
rect 18290 -430 18324 -396
rect 18290 -498 18324 -464
rect 18290 -566 18324 -532
rect 18290 -634 18324 -600
rect 9573 -770 9607 -736
rect 9573 -838 9607 -804
rect 856 -1042 890 -1008
rect 856 -1110 890 -1076
rect 856 -1178 890 -1144
rect 856 -1246 890 -1212
rect 5214 -974 5248 -940
rect 9573 -906 9607 -872
rect 13932 -702 13966 -668
rect 13932 -770 13966 -736
rect 13932 -838 13966 -804
rect 5214 -1042 5248 -1008
rect 5214 -1110 5248 -1076
rect 5214 -1178 5248 -1144
rect 5214 -1246 5248 -1212
rect 856 -1314 890 -1280
rect 856 -1382 890 -1348
rect 9573 -974 9607 -940
rect 13932 -906 13966 -872
rect 18290 -702 18324 -668
rect 18290 -770 18324 -736
rect 18290 -838 18324 -804
rect 9573 -1042 9607 -1008
rect 9573 -1110 9607 -1076
rect 9573 -1178 9607 -1144
rect 9573 -1246 9607 -1212
rect 5214 -1314 5248 -1280
rect 856 -1450 890 -1416
rect 856 -1518 890 -1484
rect 856 -1586 890 -1552
rect 5214 -1382 5248 -1348
rect 13932 -974 13966 -940
rect 18290 -906 18324 -872
rect 13932 -1042 13966 -1008
rect 13932 -1110 13966 -1076
rect 13932 -1178 13966 -1144
rect 13932 -1246 13966 -1212
rect 9573 -1314 9607 -1280
rect 5214 -1450 5248 -1416
rect 5214 -1518 5248 -1484
rect 5214 -1586 5248 -1552
rect 9573 -1382 9607 -1348
rect 18290 -974 18324 -940
rect 18290 -1042 18324 -1008
rect 18290 -1110 18324 -1076
rect 18290 -1178 18324 -1144
rect 18290 -1246 18324 -1212
rect 13932 -1314 13966 -1280
rect 9573 -1450 9607 -1416
rect 9573 -1518 9607 -1484
rect 856 -1654 890 -1620
rect 856 -1722 890 -1688
rect 856 -1790 890 -1756
rect 856 -1926 890 -1824
rect 9573 -1586 9607 -1552
rect 13932 -1382 13966 -1348
rect 18290 -1314 18324 -1280
rect 13932 -1450 13966 -1416
rect 13932 -1518 13966 -1484
rect 5214 -1654 5248 -1620
rect 5214 -1722 5248 -1688
rect 5214 -1790 5248 -1756
rect 5214 -1926 5248 -1824
rect 13932 -1586 13966 -1552
rect 18290 -1382 18324 -1348
rect 18290 -1450 18324 -1416
rect 18290 -1518 18324 -1484
rect 9573 -1654 9607 -1620
rect 9573 -1722 9607 -1688
rect 9573 -1790 9607 -1756
rect 9573 -1926 9607 -1824
rect 18290 -1586 18324 -1552
rect 13932 -1654 13966 -1620
rect 13932 -1722 13966 -1688
rect 13932 -1790 13966 -1756
rect 13932 -1926 13966 -1824
rect 18290 -1654 18324 -1620
rect 18290 -1722 18324 -1688
rect 18290 -1790 18324 -1756
rect 18290 -1926 18324 -1824
rect 856 -1960 977 -1926
rect 1011 -1960 1045 -1926
rect 1079 -1960 1113 -1926
rect 1147 -1960 1181 -1926
rect 1215 -1960 1249 -1926
rect 1283 -1960 1317 -1926
rect 1351 -1960 1385 -1926
rect 1419 -1960 1453 -1926
rect 1487 -1960 1521 -1926
rect 1555 -1960 1589 -1926
rect 1623 -1960 1657 -1926
rect 1691 -1960 1725 -1926
rect 1759 -1960 1793 -1926
rect 1827 -1960 1861 -1926
rect 1895 -1960 1929 -1926
rect 1963 -1960 1997 -1926
rect 2031 -1960 2065 -1926
rect 2099 -1960 2133 -1926
rect 2167 -1960 2201 -1926
rect 2235 -1960 2269 -1926
rect 2303 -1960 2337 -1926
rect 2371 -1960 2405 -1926
rect 2439 -1960 2473 -1926
rect 2507 -1960 2541 -1926
rect 2575 -1960 2609 -1926
rect 2643 -1960 2677 -1926
rect 2711 -1960 2745 -1926
rect 2779 -1960 2813 -1926
rect 2847 -1960 2881 -1926
rect 2915 -1960 2949 -1926
rect 2983 -1960 3017 -1926
rect 3051 -1960 3085 -1926
rect 3119 -1960 3153 -1926
rect 3187 -1960 3221 -1926
rect 3255 -1960 3289 -1926
rect 3323 -1960 3357 -1926
rect 3391 -1960 3425 -1926
rect 3459 -1960 3493 -1926
rect 3527 -1960 3561 -1926
rect 3595 -1960 3629 -1926
rect 3663 -1960 3697 -1926
rect 3731 -1960 3765 -1926
rect 3799 -1960 3833 -1926
rect 3867 -1960 3901 -1926
rect 3935 -1960 3969 -1926
rect 4003 -1960 4037 -1926
rect 4071 -1960 4105 -1926
rect 4139 -1960 4173 -1926
rect 4207 -1960 4241 -1926
rect 4275 -1960 4309 -1926
rect 4343 -1960 4377 -1926
rect 4411 -1960 4445 -1926
rect 4479 -1960 4513 -1926
rect 4547 -1960 4581 -1926
rect 4615 -1960 4649 -1926
rect 4683 -1960 4717 -1926
rect 4751 -1960 4785 -1926
rect 4819 -1960 4853 -1926
rect 4887 -1960 4921 -1926
rect 4955 -1960 4989 -1926
rect 5023 -1960 5057 -1926
rect 5091 -1960 5372 -1926
rect 5406 -1960 5440 -1926
rect 5474 -1960 5508 -1926
rect 5542 -1960 5576 -1926
rect 5610 -1960 5644 -1926
rect 5678 -1960 5712 -1926
rect 5746 -1960 5780 -1926
rect 5814 -1960 5848 -1926
rect 5882 -1960 5916 -1926
rect 5950 -1960 5984 -1926
rect 6018 -1960 6052 -1926
rect 6086 -1960 6120 -1926
rect 6154 -1960 6188 -1926
rect 6222 -1960 6256 -1926
rect 6290 -1960 6324 -1926
rect 6358 -1960 6392 -1926
rect 6426 -1960 6460 -1926
rect 6494 -1960 6528 -1926
rect 6562 -1960 6596 -1926
rect 6630 -1960 6664 -1926
rect 6698 -1960 6732 -1926
rect 6766 -1960 6800 -1926
rect 6834 -1960 6868 -1926
rect 6902 -1960 6936 -1926
rect 6970 -1960 7004 -1926
rect 7038 -1960 7072 -1926
rect 7106 -1960 7140 -1926
rect 7174 -1960 7208 -1926
rect 7242 -1960 7276 -1926
rect 7310 -1960 7344 -1926
rect 7378 -1960 7412 -1926
rect 7446 -1960 7480 -1926
rect 7514 -1960 7548 -1926
rect 7582 -1960 7616 -1926
rect 7650 -1960 7684 -1926
rect 7718 -1960 7752 -1926
rect 7786 -1960 7820 -1926
rect 7854 -1960 7888 -1926
rect 7922 -1960 7956 -1926
rect 7990 -1960 8024 -1926
rect 8058 -1960 8092 -1926
rect 8126 -1960 8160 -1926
rect 8194 -1960 8228 -1926
rect 8262 -1960 8296 -1926
rect 8330 -1960 8364 -1926
rect 8398 -1960 8432 -1926
rect 8466 -1960 8500 -1926
rect 8534 -1960 8568 -1926
rect 8602 -1960 8636 -1926
rect 8670 -1960 8704 -1926
rect 8738 -1960 8772 -1926
rect 8806 -1960 8840 -1926
rect 8874 -1960 8908 -1926
rect 8942 -1960 8976 -1926
rect 9010 -1960 9044 -1926
rect 9078 -1960 9112 -1926
rect 9146 -1960 9180 -1926
rect 9214 -1960 9248 -1926
rect 9282 -1960 9316 -1926
rect 9350 -1960 9384 -1926
rect 9418 -1960 9452 -1926
rect 9486 -1960 9694 -1926
rect 9728 -1960 9762 -1926
rect 9796 -1960 9830 -1926
rect 9864 -1960 9898 -1926
rect 9932 -1960 9966 -1926
rect 10000 -1960 10034 -1926
rect 10068 -1960 10102 -1926
rect 10136 -1960 10170 -1926
rect 10204 -1960 10238 -1926
rect 10272 -1960 10306 -1926
rect 10340 -1960 10374 -1926
rect 10408 -1960 10442 -1926
rect 10476 -1960 10510 -1926
rect 10544 -1960 10578 -1926
rect 10612 -1960 10646 -1926
rect 10680 -1960 10714 -1926
rect 10748 -1960 10782 -1926
rect 10816 -1960 10850 -1926
rect 10884 -1960 10918 -1926
rect 10952 -1960 10986 -1926
rect 11020 -1960 11054 -1926
rect 11088 -1960 11122 -1926
rect 11156 -1960 11190 -1926
rect 11224 -1960 11258 -1926
rect 11292 -1960 11326 -1926
rect 11360 -1960 11394 -1926
rect 11428 -1960 11462 -1926
rect 11496 -1960 11530 -1926
rect 11564 -1960 11598 -1926
rect 11632 -1960 11666 -1926
rect 11700 -1960 11734 -1926
rect 11768 -1960 11802 -1926
rect 11836 -1960 11870 -1926
rect 11904 -1960 11938 -1926
rect 11972 -1960 12006 -1926
rect 12040 -1960 12074 -1926
rect 12108 -1960 12142 -1926
rect 12176 -1960 12210 -1926
rect 12244 -1960 12278 -1926
rect 12312 -1960 12346 -1926
rect 12380 -1960 12414 -1926
rect 12448 -1960 12482 -1926
rect 12516 -1960 12550 -1926
rect 12584 -1960 12618 -1926
rect 12652 -1960 12686 -1926
rect 12720 -1960 12754 -1926
rect 12788 -1960 12822 -1926
rect 12856 -1960 12890 -1926
rect 12924 -1960 12958 -1926
rect 12992 -1960 13026 -1926
rect 13060 -1960 13094 -1926
rect 13128 -1960 13162 -1926
rect 13196 -1960 13230 -1926
rect 13264 -1960 13298 -1926
rect 13332 -1960 13366 -1926
rect 13400 -1960 13434 -1926
rect 13468 -1960 13502 -1926
rect 13536 -1960 13570 -1926
rect 13604 -1960 13638 -1926
rect 13672 -1960 13706 -1926
rect 13740 -1960 13774 -1926
rect 13808 -1960 14089 -1926
rect 14123 -1960 14157 -1926
rect 14191 -1960 14225 -1926
rect 14259 -1960 14293 -1926
rect 14327 -1960 14361 -1926
rect 14395 -1960 14429 -1926
rect 14463 -1960 14497 -1926
rect 14531 -1960 14565 -1926
rect 14599 -1960 14633 -1926
rect 14667 -1960 14701 -1926
rect 14735 -1960 14769 -1926
rect 14803 -1960 14837 -1926
rect 14871 -1960 14905 -1926
rect 14939 -1960 14973 -1926
rect 15007 -1960 15041 -1926
rect 15075 -1960 15109 -1926
rect 15143 -1960 15177 -1926
rect 15211 -1960 15245 -1926
rect 15279 -1960 15313 -1926
rect 15347 -1960 15381 -1926
rect 15415 -1960 15449 -1926
rect 15483 -1960 15517 -1926
rect 15551 -1960 15585 -1926
rect 15619 -1960 15653 -1926
rect 15687 -1960 15721 -1926
rect 15755 -1960 15789 -1926
rect 15823 -1960 15857 -1926
rect 15891 -1960 15925 -1926
rect 15959 -1960 15993 -1926
rect 16027 -1960 16061 -1926
rect 16095 -1960 16129 -1926
rect 16163 -1960 16197 -1926
rect 16231 -1960 16265 -1926
rect 16299 -1960 16333 -1926
rect 16367 -1960 16401 -1926
rect 16435 -1960 16469 -1926
rect 16503 -1960 16537 -1926
rect 16571 -1960 16605 -1926
rect 16639 -1960 16673 -1926
rect 16707 -1960 16741 -1926
rect 16775 -1960 16809 -1926
rect 16843 -1960 16877 -1926
rect 16911 -1960 16945 -1926
rect 16979 -1960 17013 -1926
rect 17047 -1960 17081 -1926
rect 17115 -1960 17149 -1926
rect 17183 -1960 17217 -1926
rect 17251 -1960 17285 -1926
rect 17319 -1960 17353 -1926
rect 17387 -1960 17421 -1926
rect 17455 -1960 17489 -1926
rect 17523 -1960 17557 -1926
rect 17591 -1960 17625 -1926
rect 17659 -1960 17693 -1926
rect 17727 -1960 17761 -1926
rect 17795 -1960 17829 -1926
rect 17863 -1960 17897 -1926
rect 17931 -1960 17965 -1926
rect 17999 -1960 18033 -1926
rect 18067 -1960 18101 -1926
rect 18135 -1960 18169 -1926
rect 18203 -1960 18324 -1926
rect 856 -2062 890 -1960
rect 856 -2130 890 -2096
rect 856 -2198 890 -2164
rect 856 -2266 890 -2232
rect 5214 -2062 5248 -1960
rect 5214 -2130 5248 -2096
rect 5214 -2198 5248 -2164
rect 5214 -2266 5248 -2232
rect 856 -2334 890 -2300
rect 9573 -2062 9607 -1960
rect 9573 -2130 9607 -2096
rect 9573 -2198 9607 -2164
rect 9573 -2266 9607 -2232
rect 856 -2402 890 -2368
rect 856 -2470 890 -2436
rect 856 -2538 890 -2504
rect 5214 -2334 5248 -2300
rect 13932 -2062 13966 -1960
rect 13932 -2130 13966 -2096
rect 13932 -2198 13966 -2164
rect 13932 -2266 13966 -2232
rect 5214 -2402 5248 -2368
rect 5214 -2470 5248 -2436
rect 856 -2606 890 -2572
rect 5214 -2538 5248 -2504
rect 9573 -2334 9607 -2300
rect 18290 -2062 18324 -1960
rect 18290 -2130 18324 -2096
rect 18290 -2198 18324 -2164
rect 18290 -2266 18324 -2232
rect 9573 -2402 9607 -2368
rect 9573 -2470 9607 -2436
rect 5214 -2606 5248 -2572
rect 856 -2674 890 -2640
rect 856 -2742 890 -2708
rect 856 -2810 890 -2776
rect 856 -2878 890 -2844
rect 856 -2946 890 -2912
rect 9573 -2538 9607 -2504
rect 13932 -2334 13966 -2300
rect 13932 -2402 13966 -2368
rect 13932 -2470 13966 -2436
rect 9573 -2606 9607 -2572
rect 5214 -2674 5248 -2640
rect 5214 -2742 5248 -2708
rect 5214 -2810 5248 -2776
rect 5214 -2878 5248 -2844
rect 856 -3014 890 -2980
rect 5214 -2946 5248 -2912
rect 13932 -2538 13966 -2504
rect 18290 -2334 18324 -2300
rect 18290 -2402 18324 -2368
rect 18290 -2470 18324 -2436
rect 13932 -2606 13966 -2572
rect 9573 -2674 9607 -2640
rect 9573 -2742 9607 -2708
rect 9573 -2810 9607 -2776
rect 9573 -2878 9607 -2844
rect 5214 -3014 5248 -2980
rect 9573 -2946 9607 -2912
rect 18290 -2538 18324 -2504
rect 18290 -2606 18324 -2572
rect 13932 -2674 13966 -2640
rect 13932 -2742 13966 -2708
rect 13932 -2810 13966 -2776
rect 13932 -2878 13966 -2844
rect 9573 -3014 9607 -2980
rect 13932 -2946 13966 -2912
rect 18290 -2674 18324 -2640
rect 18290 -2742 18324 -2708
rect 18290 -2810 18324 -2776
rect 18290 -2878 18324 -2844
rect 13932 -3014 13966 -2980
rect 18290 -2946 18324 -2912
rect 18290 -3014 18324 -2980
rect 856 -3082 890 -3048
rect 856 -3150 890 -3116
rect 856 -3218 890 -3184
rect 5214 -3082 5248 -3048
rect 5214 -3150 5248 -3116
rect 5214 -3218 5248 -3184
rect 9573 -3082 9607 -3048
rect 9573 -3150 9607 -3116
rect 856 -3286 890 -3252
rect 856 -3354 890 -3320
rect 856 -3422 890 -3388
rect 856 -3490 890 -3456
rect 856 -3558 890 -3524
rect 9573 -3218 9607 -3184
rect 13932 -3082 13966 -3048
rect 13932 -3150 13966 -3116
rect 5214 -3286 5248 -3252
rect 5214 -3354 5248 -3320
rect 5214 -3422 5248 -3388
rect 5214 -3490 5248 -3456
rect 5214 -3558 5248 -3524
rect 13932 -3218 13966 -3184
rect 18290 -3082 18324 -3048
rect 18290 -3150 18324 -3116
rect 9573 -3286 9607 -3252
rect 9573 -3354 9607 -3320
rect 9573 -3422 9607 -3388
rect 9573 -3490 9607 -3456
rect 9573 -3558 9607 -3524
rect 18290 -3218 18324 -3184
rect 13932 -3286 13966 -3252
rect 13932 -3354 13966 -3320
rect 13932 -3422 13966 -3388
rect 13932 -3490 13966 -3456
rect 13932 -3558 13966 -3524
rect 18290 -3286 18324 -3252
rect 18290 -3354 18324 -3320
rect 18290 -3422 18324 -3388
rect 18290 -3490 18324 -3456
rect 18290 -3558 18324 -3524
rect 856 -3626 977 -3592
rect 1011 -3626 1045 -3592
rect 1079 -3626 1113 -3592
rect 1147 -3626 1181 -3592
rect 1215 -3626 1249 -3592
rect 1283 -3626 1317 -3592
rect 1351 -3626 1385 -3592
rect 1419 -3626 1453 -3592
rect 1487 -3626 1521 -3592
rect 1555 -3626 1589 -3592
rect 1623 -3626 1657 -3592
rect 1691 -3626 1725 -3592
rect 1759 -3626 1793 -3592
rect 1827 -3626 1861 -3592
rect 1895 -3626 1929 -3592
rect 1963 -3626 1997 -3592
rect 2031 -3626 2065 -3592
rect 2099 -3626 2133 -3592
rect 2167 -3626 2201 -3592
rect 2235 -3626 2269 -3592
rect 2303 -3626 2337 -3592
rect 2371 -3626 2405 -3592
rect 2439 -3626 2473 -3592
rect 2507 -3626 2541 -3592
rect 2575 -3626 2609 -3592
rect 2643 -3626 2677 -3592
rect 2711 -3626 2745 -3592
rect 2779 -3626 2813 -3592
rect 2847 -3626 2881 -3592
rect 2915 -3626 2949 -3592
rect 2983 -3626 3017 -3592
rect 3051 -3626 3085 -3592
rect 3119 -3626 3153 -3592
rect 3187 -3626 3221 -3592
rect 3255 -3626 3289 -3592
rect 3323 -3626 3357 -3592
rect 3391 -3626 3425 -3592
rect 3459 -3626 3493 -3592
rect 3527 -3626 3561 -3592
rect 3595 -3626 3629 -3592
rect 3663 -3626 3697 -3592
rect 3731 -3626 3765 -3592
rect 3799 -3626 3833 -3592
rect 3867 -3626 3901 -3592
rect 3935 -3626 3969 -3592
rect 4003 -3626 4037 -3592
rect 4071 -3626 4105 -3592
rect 4139 -3626 4173 -3592
rect 4207 -3626 4241 -3592
rect 4275 -3626 4309 -3592
rect 4343 -3626 4377 -3592
rect 4411 -3626 4445 -3592
rect 4479 -3626 4513 -3592
rect 4547 -3626 4581 -3592
rect 4615 -3626 4649 -3592
rect 4683 -3626 4717 -3592
rect 4751 -3626 4785 -3592
rect 4819 -3626 4853 -3592
rect 4887 -3626 4921 -3592
rect 4955 -3626 4989 -3592
rect 5023 -3626 5057 -3592
rect 5091 -3626 5372 -3592
rect 5406 -3626 5440 -3592
rect 5474 -3626 5508 -3592
rect 5542 -3626 5576 -3592
rect 5610 -3626 5644 -3592
rect 5678 -3626 5712 -3592
rect 5746 -3626 5780 -3592
rect 5814 -3626 5848 -3592
rect 5882 -3626 5916 -3592
rect 5950 -3626 5984 -3592
rect 6018 -3626 6052 -3592
rect 6086 -3626 6120 -3592
rect 6154 -3626 6188 -3592
rect 6222 -3626 6256 -3592
rect 6290 -3626 6324 -3592
rect 6358 -3626 6392 -3592
rect 6426 -3626 6460 -3592
rect 6494 -3626 6528 -3592
rect 6562 -3626 6596 -3592
rect 6630 -3626 6664 -3592
rect 6698 -3626 6732 -3592
rect 6766 -3626 6800 -3592
rect 6834 -3626 6868 -3592
rect 6902 -3626 6936 -3592
rect 6970 -3626 7004 -3592
rect 7038 -3626 7072 -3592
rect 7106 -3626 7140 -3592
rect 7174 -3626 7208 -3592
rect 7242 -3626 7276 -3592
rect 7310 -3626 7344 -3592
rect 7378 -3626 7412 -3592
rect 7446 -3626 7480 -3592
rect 7514 -3626 7548 -3592
rect 7582 -3626 7616 -3592
rect 7650 -3626 7684 -3592
rect 7718 -3626 7752 -3592
rect 7786 -3626 7820 -3592
rect 7854 -3626 7888 -3592
rect 7922 -3626 7956 -3592
rect 7990 -3626 8024 -3592
rect 8058 -3626 8092 -3592
rect 8126 -3626 8160 -3592
rect 8194 -3626 8228 -3592
rect 8262 -3626 8296 -3592
rect 8330 -3626 8364 -3592
rect 8398 -3626 8432 -3592
rect 8466 -3626 8500 -3592
rect 8534 -3626 8568 -3592
rect 8602 -3626 8636 -3592
rect 8670 -3626 8704 -3592
rect 8738 -3626 8772 -3592
rect 8806 -3626 8840 -3592
rect 8874 -3626 8908 -3592
rect 8942 -3626 8976 -3592
rect 9010 -3626 9044 -3592
rect 9078 -3626 9112 -3592
rect 9146 -3626 9180 -3592
rect 9214 -3626 9248 -3592
rect 9282 -3626 9316 -3592
rect 9350 -3626 9384 -3592
rect 9418 -3626 9452 -3592
rect 9486 -3626 9694 -3592
rect 9728 -3626 9762 -3592
rect 9796 -3626 9830 -3592
rect 9864 -3626 9898 -3592
rect 9932 -3626 9966 -3592
rect 10000 -3626 10034 -3592
rect 10068 -3626 10102 -3592
rect 10136 -3626 10170 -3592
rect 10204 -3626 10238 -3592
rect 10272 -3626 10306 -3592
rect 10340 -3626 10374 -3592
rect 10408 -3626 10442 -3592
rect 10476 -3626 10510 -3592
rect 10544 -3626 10578 -3592
rect 10612 -3626 10646 -3592
rect 10680 -3626 10714 -3592
rect 10748 -3626 10782 -3592
rect 10816 -3626 10850 -3592
rect 10884 -3626 10918 -3592
rect 10952 -3626 10986 -3592
rect 11020 -3626 11054 -3592
rect 11088 -3626 11122 -3592
rect 11156 -3626 11190 -3592
rect 11224 -3626 11258 -3592
rect 11292 -3626 11326 -3592
rect 11360 -3626 11394 -3592
rect 11428 -3626 11462 -3592
rect 11496 -3626 11530 -3592
rect 11564 -3626 11598 -3592
rect 11632 -3626 11666 -3592
rect 11700 -3626 11734 -3592
rect 11768 -3626 11802 -3592
rect 11836 -3626 11870 -3592
rect 11904 -3626 11938 -3592
rect 11972 -3626 12006 -3592
rect 12040 -3626 12074 -3592
rect 12108 -3626 12142 -3592
rect 12176 -3626 12210 -3592
rect 12244 -3626 12278 -3592
rect 12312 -3626 12346 -3592
rect 12380 -3626 12414 -3592
rect 12448 -3626 12482 -3592
rect 12516 -3626 12550 -3592
rect 12584 -3626 12618 -3592
rect 12652 -3626 12686 -3592
rect 12720 -3626 12754 -3592
rect 12788 -3626 12822 -3592
rect 12856 -3626 12890 -3592
rect 12924 -3626 12958 -3592
rect 12992 -3626 13026 -3592
rect 13060 -3626 13094 -3592
rect 13128 -3626 13162 -3592
rect 13196 -3626 13230 -3592
rect 13264 -3626 13298 -3592
rect 13332 -3626 13366 -3592
rect 13400 -3626 13434 -3592
rect 13468 -3626 13502 -3592
rect 13536 -3626 13570 -3592
rect 13604 -3626 13638 -3592
rect 13672 -3626 13706 -3592
rect 13740 -3626 13774 -3592
rect 13808 -3626 14089 -3592
rect 14123 -3626 14157 -3592
rect 14191 -3626 14225 -3592
rect 14259 -3626 14293 -3592
rect 14327 -3626 14361 -3592
rect 14395 -3626 14429 -3592
rect 14463 -3626 14497 -3592
rect 14531 -3626 14565 -3592
rect 14599 -3626 14633 -3592
rect 14667 -3626 14701 -3592
rect 14735 -3626 14769 -3592
rect 14803 -3626 14837 -3592
rect 14871 -3626 14905 -3592
rect 14939 -3626 14973 -3592
rect 15007 -3626 15041 -3592
rect 15075 -3626 15109 -3592
rect 15143 -3626 15177 -3592
rect 15211 -3626 15245 -3592
rect 15279 -3626 15313 -3592
rect 15347 -3626 15381 -3592
rect 15415 -3626 15449 -3592
rect 15483 -3626 15517 -3592
rect 15551 -3626 15585 -3592
rect 15619 -3626 15653 -3592
rect 15687 -3626 15721 -3592
rect 15755 -3626 15789 -3592
rect 15823 -3626 15857 -3592
rect 15891 -3626 15925 -3592
rect 15959 -3626 15993 -3592
rect 16027 -3626 16061 -3592
rect 16095 -3626 16129 -3592
rect 16163 -3626 16197 -3592
rect 16231 -3626 16265 -3592
rect 16299 -3626 16333 -3592
rect 16367 -3626 16401 -3592
rect 16435 -3626 16469 -3592
rect 16503 -3626 16537 -3592
rect 16571 -3626 16605 -3592
rect 16639 -3626 16673 -3592
rect 16707 -3626 16741 -3592
rect 16775 -3626 16809 -3592
rect 16843 -3626 16877 -3592
rect 16911 -3626 16945 -3592
rect 16979 -3626 17013 -3592
rect 17047 -3626 17081 -3592
rect 17115 -3626 17149 -3592
rect 17183 -3626 17217 -3592
rect 17251 -3626 17285 -3592
rect 17319 -3626 17353 -3592
rect 17387 -3626 17421 -3592
rect 17455 -3626 17489 -3592
rect 17523 -3626 17557 -3592
rect 17591 -3626 17625 -3592
rect 17659 -3626 17693 -3592
rect 17727 -3626 17761 -3592
rect 17795 -3626 17829 -3592
rect 17863 -3626 17897 -3592
rect 17931 -3626 17965 -3592
rect 17999 -3626 18033 -3592
rect 18067 -3626 18101 -3592
rect 18135 -3626 18169 -3592
rect 18203 -3626 18324 -3592
rect 856 -3694 890 -3660
rect 856 -3762 890 -3728
rect 856 -3830 890 -3796
rect 856 -3898 890 -3864
rect 856 -3966 890 -3932
rect 5214 -3694 5248 -3660
rect 5214 -3762 5248 -3728
rect 5214 -3830 5248 -3796
rect 5214 -3898 5248 -3864
rect 5214 -3966 5248 -3932
rect 856 -4034 890 -4000
rect 9573 -3694 9607 -3660
rect 9573 -3762 9607 -3728
rect 9573 -3830 9607 -3796
rect 9573 -3898 9607 -3864
rect 9573 -3966 9607 -3932
rect 856 -4102 890 -4068
rect 856 -4365 890 -4136
rect 5214 -4034 5248 -4000
rect 13932 -3694 13966 -3660
rect 13932 -3762 13966 -3728
rect 13932 -3830 13966 -3796
rect 13932 -3898 13966 -3864
rect 13932 -3966 13966 -3932
rect 5214 -4102 5248 -4068
rect 5214 -4365 5248 -4136
rect 9573 -4034 9607 -4000
rect 18290 -3694 18324 -3660
rect 18290 -3762 18324 -3728
rect 18290 -3830 18324 -3796
rect 18290 -3898 18324 -3864
rect 18290 -3966 18324 -3932
rect 9573 -4102 9607 -4068
rect 9573 -4365 9607 -4136
rect 13932 -4034 13966 -4000
rect 13932 -4102 13966 -4068
rect 13932 -4365 13966 -4136
rect 18290 -4034 18324 -4000
rect 18290 -4102 18324 -4068
rect 18290 -4365 18324 -4136
rect 856 -4399 977 -4365
rect 1011 -4399 1045 -4365
rect 1079 -4399 1113 -4365
rect 1147 -4399 1181 -4365
rect 1215 -4399 1249 -4365
rect 1283 -4399 1317 -4365
rect 1351 -4399 1385 -4365
rect 1419 -4399 1453 -4365
rect 1487 -4399 1521 -4365
rect 1555 -4399 1589 -4365
rect 1623 -4399 1657 -4365
rect 1691 -4399 1725 -4365
rect 1759 -4399 1793 -4365
rect 1827 -4399 1861 -4365
rect 1895 -4399 1929 -4365
rect 1963 -4399 1997 -4365
rect 2031 -4399 2065 -4365
rect 2099 -4399 2133 -4365
rect 2167 -4399 2201 -4365
rect 2235 -4399 2269 -4365
rect 2303 -4399 2337 -4365
rect 2371 -4399 2405 -4365
rect 2439 -4399 2473 -4365
rect 2507 -4399 2541 -4365
rect 2575 -4399 2609 -4365
rect 2643 -4399 2677 -4365
rect 2711 -4399 2745 -4365
rect 2779 -4399 2813 -4365
rect 2847 -4399 2881 -4365
rect 2915 -4399 2949 -4365
rect 2983 -4399 3017 -4365
rect 3051 -4399 3085 -4365
rect 3119 -4399 3153 -4365
rect 3187 -4399 3221 -4365
rect 3255 -4399 3289 -4365
rect 3323 -4399 3357 -4365
rect 3391 -4399 3425 -4365
rect 3459 -4399 3493 -4365
rect 3527 -4399 3561 -4365
rect 3595 -4399 3629 -4365
rect 3663 -4399 3697 -4365
rect 3731 -4399 3765 -4365
rect 3799 -4399 3833 -4365
rect 3867 -4399 3901 -4365
rect 3935 -4399 3969 -4365
rect 4003 -4399 4037 -4365
rect 4071 -4399 4105 -4365
rect 4139 -4399 4173 -4365
rect 4207 -4399 4241 -4365
rect 4275 -4399 4309 -4365
rect 4343 -4399 4377 -4365
rect 4411 -4399 4445 -4365
rect 4479 -4399 4513 -4365
rect 4547 -4399 4581 -4365
rect 4615 -4399 4649 -4365
rect 4683 -4399 4717 -4365
rect 4751 -4399 4785 -4365
rect 4819 -4399 4853 -4365
rect 4887 -4399 4921 -4365
rect 4955 -4399 4989 -4365
rect 5023 -4399 5057 -4365
rect 5091 -4399 5372 -4365
rect 5406 -4399 5440 -4365
rect 5474 -4399 5508 -4365
rect 5542 -4399 5576 -4365
rect 5610 -4399 5644 -4365
rect 5678 -4399 5712 -4365
rect 5746 -4399 5780 -4365
rect 5814 -4399 5848 -4365
rect 5882 -4399 5916 -4365
rect 5950 -4399 5984 -4365
rect 6018 -4399 6052 -4365
rect 6086 -4399 6120 -4365
rect 6154 -4399 6188 -4365
rect 6222 -4399 6256 -4365
rect 6290 -4399 6324 -4365
rect 6358 -4399 6392 -4365
rect 6426 -4399 6460 -4365
rect 6494 -4399 6528 -4365
rect 6562 -4399 6596 -4365
rect 6630 -4399 6664 -4365
rect 6698 -4399 6732 -4365
rect 6766 -4399 6800 -4365
rect 6834 -4399 6868 -4365
rect 6902 -4399 6936 -4365
rect 6970 -4399 7004 -4365
rect 7038 -4399 7072 -4365
rect 7106 -4399 7140 -4365
rect 7174 -4399 7208 -4365
rect 7242 -4399 7276 -4365
rect 7310 -4399 7344 -4365
rect 7378 -4399 7412 -4365
rect 7446 -4399 7480 -4365
rect 7514 -4399 7548 -4365
rect 7582 -4399 7616 -4365
rect 7650 -4399 7684 -4365
rect 7718 -4399 7752 -4365
rect 7786 -4399 7820 -4365
rect 7854 -4399 7888 -4365
rect 7922 -4399 7956 -4365
rect 7990 -4399 8024 -4365
rect 8058 -4399 8092 -4365
rect 8126 -4399 8160 -4365
rect 8194 -4399 8228 -4365
rect 8262 -4399 8296 -4365
rect 8330 -4399 8364 -4365
rect 8398 -4399 8432 -4365
rect 8466 -4399 8500 -4365
rect 8534 -4399 8568 -4365
rect 8602 -4399 8636 -4365
rect 8670 -4399 8704 -4365
rect 8738 -4399 8772 -4365
rect 8806 -4399 8840 -4365
rect 8874 -4399 8908 -4365
rect 8942 -4399 8976 -4365
rect 9010 -4399 9044 -4365
rect 9078 -4399 9112 -4365
rect 9146 -4399 9180 -4365
rect 9214 -4399 9248 -4365
rect 9282 -4399 9316 -4365
rect 9350 -4399 9384 -4365
rect 9418 -4399 9452 -4365
rect 9486 -4399 9694 -4365
rect 9728 -4399 9762 -4365
rect 9796 -4399 9830 -4365
rect 9864 -4399 9898 -4365
rect 9932 -4399 9966 -4365
rect 10000 -4399 10034 -4365
rect 10068 -4399 10102 -4365
rect 10136 -4399 10170 -4365
rect 10204 -4399 10238 -4365
rect 10272 -4399 10306 -4365
rect 10340 -4399 10374 -4365
rect 10408 -4399 10442 -4365
rect 10476 -4399 10510 -4365
rect 10544 -4399 10578 -4365
rect 10612 -4399 10646 -4365
rect 10680 -4399 10714 -4365
rect 10748 -4399 10782 -4365
rect 10816 -4399 10850 -4365
rect 10884 -4399 10918 -4365
rect 10952 -4399 10986 -4365
rect 11020 -4399 11054 -4365
rect 11088 -4399 11122 -4365
rect 11156 -4399 11190 -4365
rect 11224 -4399 11258 -4365
rect 11292 -4399 11326 -4365
rect 11360 -4399 11394 -4365
rect 11428 -4399 11462 -4365
rect 11496 -4399 11530 -4365
rect 11564 -4399 11598 -4365
rect 11632 -4399 11666 -4365
rect 11700 -4399 11734 -4365
rect 11768 -4399 11802 -4365
rect 11836 -4399 11870 -4365
rect 11904 -4399 11938 -4365
rect 11972 -4399 12006 -4365
rect 12040 -4399 12074 -4365
rect 12108 -4399 12142 -4365
rect 12176 -4399 12210 -4365
rect 12244 -4399 12278 -4365
rect 12312 -4399 12346 -4365
rect 12380 -4399 12414 -4365
rect 12448 -4399 12482 -4365
rect 12516 -4399 12550 -4365
rect 12584 -4399 12618 -4365
rect 12652 -4399 12686 -4365
rect 12720 -4399 12754 -4365
rect 12788 -4399 12822 -4365
rect 12856 -4399 12890 -4365
rect 12924 -4399 12958 -4365
rect 12992 -4399 13026 -4365
rect 13060 -4399 13094 -4365
rect 13128 -4399 13162 -4365
rect 13196 -4399 13230 -4365
rect 13264 -4399 13298 -4365
rect 13332 -4399 13366 -4365
rect 13400 -4399 13434 -4365
rect 13468 -4399 13502 -4365
rect 13536 -4399 13570 -4365
rect 13604 -4399 13638 -4365
rect 13672 -4399 13706 -4365
rect 13740 -4399 13774 -4365
rect 13808 -4399 14089 -4365
rect 14123 -4399 14157 -4365
rect 14191 -4399 14225 -4365
rect 14259 -4399 14293 -4365
rect 14327 -4399 14361 -4365
rect 14395 -4399 14429 -4365
rect 14463 -4399 14497 -4365
rect 14531 -4399 14565 -4365
rect 14599 -4399 14633 -4365
rect 14667 -4399 14701 -4365
rect 14735 -4399 14769 -4365
rect 14803 -4399 14837 -4365
rect 14871 -4399 14905 -4365
rect 14939 -4399 14973 -4365
rect 15007 -4399 15041 -4365
rect 15075 -4399 15109 -4365
rect 15143 -4399 15177 -4365
rect 15211 -4399 15245 -4365
rect 15279 -4399 15313 -4365
rect 15347 -4399 15381 -4365
rect 15415 -4399 15449 -4365
rect 15483 -4399 15517 -4365
rect 15551 -4399 15585 -4365
rect 15619 -4399 15653 -4365
rect 15687 -4399 15721 -4365
rect 15755 -4399 15789 -4365
rect 15823 -4399 15857 -4365
rect 15891 -4399 15925 -4365
rect 15959 -4399 15993 -4365
rect 16027 -4399 16061 -4365
rect 16095 -4399 16129 -4365
rect 16163 -4399 16197 -4365
rect 16231 -4399 16265 -4365
rect 16299 -4399 16333 -4365
rect 16367 -4399 16401 -4365
rect 16435 -4399 16469 -4365
rect 16503 -4399 16537 -4365
rect 16571 -4399 16605 -4365
rect 16639 -4399 16673 -4365
rect 16707 -4399 16741 -4365
rect 16775 -4399 16809 -4365
rect 16843 -4399 16877 -4365
rect 16911 -4399 16945 -4365
rect 16979 -4399 17013 -4365
rect 17047 -4399 17081 -4365
rect 17115 -4399 17149 -4365
rect 17183 -4399 17217 -4365
rect 17251 -4399 17285 -4365
rect 17319 -4399 17353 -4365
rect 17387 -4399 17421 -4365
rect 17455 -4399 17489 -4365
rect 17523 -4399 17557 -4365
rect 17591 -4399 17625 -4365
rect 17659 -4399 17693 -4365
rect 17727 -4399 17761 -4365
rect 17795 -4399 17829 -4365
rect 17863 -4399 17897 -4365
rect 17931 -4399 17965 -4365
rect 17999 -4399 18033 -4365
rect 18067 -4399 18101 -4365
rect 18135 -4399 18169 -4365
rect 18203 -4399 18324 -4365
rect 856 -4628 890 -4399
rect 856 -4696 890 -4662
rect 856 -4764 890 -4730
rect 5214 -4628 5248 -4399
rect 5214 -4696 5248 -4662
rect 5214 -4764 5248 -4730
rect 9573 -4628 9607 -4399
rect 9573 -4696 9607 -4662
rect 856 -4832 890 -4798
rect 856 -4900 890 -4866
rect 856 -4968 890 -4934
rect 856 -5036 890 -5002
rect 856 -5104 890 -5070
rect 9573 -4764 9607 -4730
rect 13932 -4628 13966 -4399
rect 13932 -4696 13966 -4662
rect 5214 -4832 5248 -4798
rect 5214 -4900 5248 -4866
rect 5214 -4968 5248 -4934
rect 5214 -5036 5248 -5002
rect 5214 -5104 5248 -5070
rect 13932 -4764 13966 -4730
rect 18290 -4628 18324 -4399
rect 18290 -4696 18324 -4662
rect 9573 -4832 9607 -4798
rect 9573 -4900 9607 -4866
rect 9573 -4968 9607 -4934
rect 9573 -5036 9607 -5002
rect 9573 -5104 9607 -5070
rect 18290 -4764 18324 -4730
rect 13932 -4832 13966 -4798
rect 13932 -4900 13966 -4866
rect 13932 -4968 13966 -4934
rect 13932 -5036 13966 -5002
rect 13932 -5104 13966 -5070
rect 18290 -4832 18324 -4798
rect 18290 -4900 18324 -4866
rect 18290 -4968 18324 -4934
rect 18290 -5036 18324 -5002
rect 18290 -5104 18324 -5070
rect 856 -5172 977 -5138
rect 1011 -5172 1045 -5138
rect 1079 -5172 1113 -5138
rect 1147 -5172 1181 -5138
rect 1215 -5172 1249 -5138
rect 1283 -5172 1317 -5138
rect 1351 -5172 1385 -5138
rect 1419 -5172 1453 -5138
rect 1487 -5172 1521 -5138
rect 1555 -5172 1589 -5138
rect 1623 -5172 1657 -5138
rect 1691 -5172 1725 -5138
rect 1759 -5172 1793 -5138
rect 1827 -5172 1861 -5138
rect 1895 -5172 1929 -5138
rect 1963 -5172 1997 -5138
rect 2031 -5172 2065 -5138
rect 2099 -5172 2133 -5138
rect 2167 -5172 2201 -5138
rect 2235 -5172 2269 -5138
rect 2303 -5172 2337 -5138
rect 2371 -5172 2405 -5138
rect 2439 -5172 2473 -5138
rect 2507 -5172 2541 -5138
rect 2575 -5172 2609 -5138
rect 2643 -5172 2677 -5138
rect 2711 -5172 2745 -5138
rect 2779 -5172 2813 -5138
rect 2847 -5172 2881 -5138
rect 2915 -5172 2949 -5138
rect 2983 -5172 3017 -5138
rect 3051 -5172 3085 -5138
rect 3119 -5172 3153 -5138
rect 3187 -5172 3221 -5138
rect 3255 -5172 3289 -5138
rect 3323 -5172 3357 -5138
rect 3391 -5172 3425 -5138
rect 3459 -5172 3493 -5138
rect 3527 -5172 3561 -5138
rect 3595 -5172 3629 -5138
rect 3663 -5172 3697 -5138
rect 3731 -5172 3765 -5138
rect 3799 -5172 3833 -5138
rect 3867 -5172 3901 -5138
rect 3935 -5172 3969 -5138
rect 4003 -5172 4037 -5138
rect 4071 -5172 4105 -5138
rect 4139 -5172 4173 -5138
rect 4207 -5172 4241 -5138
rect 4275 -5172 4309 -5138
rect 4343 -5172 4377 -5138
rect 4411 -5172 4445 -5138
rect 4479 -5172 4513 -5138
rect 4547 -5172 4581 -5138
rect 4615 -5172 4649 -5138
rect 4683 -5172 4717 -5138
rect 4751 -5172 4785 -5138
rect 4819 -5172 4853 -5138
rect 4887 -5172 4921 -5138
rect 4955 -5172 4989 -5138
rect 5023 -5172 5057 -5138
rect 5091 -5172 5372 -5138
rect 5406 -5172 5440 -5138
rect 5474 -5172 5508 -5138
rect 5542 -5172 5576 -5138
rect 5610 -5172 5644 -5138
rect 5678 -5172 5712 -5138
rect 5746 -5172 5780 -5138
rect 5814 -5172 5848 -5138
rect 5882 -5172 5916 -5138
rect 5950 -5172 5984 -5138
rect 6018 -5172 6052 -5138
rect 6086 -5172 6120 -5138
rect 6154 -5172 6188 -5138
rect 6222 -5172 6256 -5138
rect 6290 -5172 6324 -5138
rect 6358 -5172 6392 -5138
rect 6426 -5172 6460 -5138
rect 6494 -5172 6528 -5138
rect 6562 -5172 6596 -5138
rect 6630 -5172 6664 -5138
rect 6698 -5172 6732 -5138
rect 6766 -5172 6800 -5138
rect 6834 -5172 6868 -5138
rect 6902 -5172 6936 -5138
rect 6970 -5172 7004 -5138
rect 7038 -5172 7072 -5138
rect 7106 -5172 7140 -5138
rect 7174 -5172 7208 -5138
rect 7242 -5172 7276 -5138
rect 7310 -5172 7344 -5138
rect 7378 -5172 7412 -5138
rect 7446 -5172 7480 -5138
rect 7514 -5172 7548 -5138
rect 7582 -5172 7616 -5138
rect 7650 -5172 7684 -5138
rect 7718 -5172 7752 -5138
rect 7786 -5172 7820 -5138
rect 7854 -5172 7888 -5138
rect 7922 -5172 7956 -5138
rect 7990 -5172 8024 -5138
rect 8058 -5172 8092 -5138
rect 8126 -5172 8160 -5138
rect 8194 -5172 8228 -5138
rect 8262 -5172 8296 -5138
rect 8330 -5172 8364 -5138
rect 8398 -5172 8432 -5138
rect 8466 -5172 8500 -5138
rect 8534 -5172 8568 -5138
rect 8602 -5172 8636 -5138
rect 8670 -5172 8704 -5138
rect 8738 -5172 8772 -5138
rect 8806 -5172 8840 -5138
rect 8874 -5172 8908 -5138
rect 8942 -5172 8976 -5138
rect 9010 -5172 9044 -5138
rect 9078 -5172 9112 -5138
rect 9146 -5172 9180 -5138
rect 9214 -5172 9248 -5138
rect 9282 -5172 9316 -5138
rect 9350 -5172 9384 -5138
rect 9418 -5172 9452 -5138
rect 9486 -5172 9694 -5138
rect 9728 -5172 9762 -5138
rect 9796 -5172 9830 -5138
rect 9864 -5172 9898 -5138
rect 9932 -5172 9966 -5138
rect 10000 -5172 10034 -5138
rect 10068 -5172 10102 -5138
rect 10136 -5172 10170 -5138
rect 10204 -5172 10238 -5138
rect 10272 -5172 10306 -5138
rect 10340 -5172 10374 -5138
rect 10408 -5172 10442 -5138
rect 10476 -5172 10510 -5138
rect 10544 -5172 10578 -5138
rect 10612 -5172 10646 -5138
rect 10680 -5172 10714 -5138
rect 10748 -5172 10782 -5138
rect 10816 -5172 10850 -5138
rect 10884 -5172 10918 -5138
rect 10952 -5172 10986 -5138
rect 11020 -5172 11054 -5138
rect 11088 -5172 11122 -5138
rect 11156 -5172 11190 -5138
rect 11224 -5172 11258 -5138
rect 11292 -5172 11326 -5138
rect 11360 -5172 11394 -5138
rect 11428 -5172 11462 -5138
rect 11496 -5172 11530 -5138
rect 11564 -5172 11598 -5138
rect 11632 -5172 11666 -5138
rect 11700 -5172 11734 -5138
rect 11768 -5172 11802 -5138
rect 11836 -5172 11870 -5138
rect 11904 -5172 11938 -5138
rect 11972 -5172 12006 -5138
rect 12040 -5172 12074 -5138
rect 12108 -5172 12142 -5138
rect 12176 -5172 12210 -5138
rect 12244 -5172 12278 -5138
rect 12312 -5172 12346 -5138
rect 12380 -5172 12414 -5138
rect 12448 -5172 12482 -5138
rect 12516 -5172 12550 -5138
rect 12584 -5172 12618 -5138
rect 12652 -5172 12686 -5138
rect 12720 -5172 12754 -5138
rect 12788 -5172 12822 -5138
rect 12856 -5172 12890 -5138
rect 12924 -5172 12958 -5138
rect 12992 -5172 13026 -5138
rect 13060 -5172 13094 -5138
rect 13128 -5172 13162 -5138
rect 13196 -5172 13230 -5138
rect 13264 -5172 13298 -5138
rect 13332 -5172 13366 -5138
rect 13400 -5172 13434 -5138
rect 13468 -5172 13502 -5138
rect 13536 -5172 13570 -5138
rect 13604 -5172 13638 -5138
rect 13672 -5172 13706 -5138
rect 13740 -5172 13774 -5138
rect 13808 -5172 14089 -5138
rect 14123 -5172 14157 -5138
rect 14191 -5172 14225 -5138
rect 14259 -5172 14293 -5138
rect 14327 -5172 14361 -5138
rect 14395 -5172 14429 -5138
rect 14463 -5172 14497 -5138
rect 14531 -5172 14565 -5138
rect 14599 -5172 14633 -5138
rect 14667 -5172 14701 -5138
rect 14735 -5172 14769 -5138
rect 14803 -5172 14837 -5138
rect 14871 -5172 14905 -5138
rect 14939 -5172 14973 -5138
rect 15007 -5172 15041 -5138
rect 15075 -5172 15109 -5138
rect 15143 -5172 15177 -5138
rect 15211 -5172 15245 -5138
rect 15279 -5172 15313 -5138
rect 15347 -5172 15381 -5138
rect 15415 -5172 15449 -5138
rect 15483 -5172 15517 -5138
rect 15551 -5172 15585 -5138
rect 15619 -5172 15653 -5138
rect 15687 -5172 15721 -5138
rect 15755 -5172 15789 -5138
rect 15823 -5172 15857 -5138
rect 15891 -5172 15925 -5138
rect 15959 -5172 15993 -5138
rect 16027 -5172 16061 -5138
rect 16095 -5172 16129 -5138
rect 16163 -5172 16197 -5138
rect 16231 -5172 16265 -5138
rect 16299 -5172 16333 -5138
rect 16367 -5172 16401 -5138
rect 16435 -5172 16469 -5138
rect 16503 -5172 16537 -5138
rect 16571 -5172 16605 -5138
rect 16639 -5172 16673 -5138
rect 16707 -5172 16741 -5138
rect 16775 -5172 16809 -5138
rect 16843 -5172 16877 -5138
rect 16911 -5172 16945 -5138
rect 16979 -5172 17013 -5138
rect 17047 -5172 17081 -5138
rect 17115 -5172 17149 -5138
rect 17183 -5172 17217 -5138
rect 17251 -5172 17285 -5138
rect 17319 -5172 17353 -5138
rect 17387 -5172 17421 -5138
rect 17455 -5172 17489 -5138
rect 17523 -5172 17557 -5138
rect 17591 -5172 17625 -5138
rect 17659 -5172 17693 -5138
rect 17727 -5172 17761 -5138
rect 17795 -5172 17829 -5138
rect 17863 -5172 17897 -5138
rect 17931 -5172 17965 -5138
rect 17999 -5172 18033 -5138
rect 18067 -5172 18101 -5138
rect 18135 -5172 18169 -5138
rect 18203 -5172 18324 -5138
rect 856 -5240 890 -5206
rect 856 -5308 890 -5274
rect 856 -5376 890 -5342
rect 856 -5444 890 -5410
rect 856 -5512 890 -5478
rect 5214 -5240 5248 -5206
rect 5214 -5308 5248 -5274
rect 5214 -5376 5248 -5342
rect 5214 -5444 5248 -5410
rect 5214 -5512 5248 -5478
rect 856 -5580 890 -5546
rect 9573 -5240 9607 -5206
rect 9573 -5308 9607 -5274
rect 9573 -5376 9607 -5342
rect 9573 -5444 9607 -5410
rect 9573 -5512 9607 -5478
rect 856 -5648 890 -5614
rect 856 -5716 890 -5682
rect 5214 -5580 5248 -5546
rect 13932 -5240 13966 -5206
rect 13932 -5308 13966 -5274
rect 13932 -5376 13966 -5342
rect 13932 -5444 13966 -5410
rect 13932 -5512 13966 -5478
rect 5214 -5648 5248 -5614
rect 5214 -5716 5248 -5682
rect 9573 -5580 9607 -5546
rect 18290 -5240 18324 -5206
rect 18290 -5308 18324 -5274
rect 18290 -5376 18324 -5342
rect 18290 -5444 18324 -5410
rect 18290 -5512 18324 -5478
rect 9573 -5648 9607 -5614
rect 9573 -5716 9607 -5682
rect 13932 -5580 13966 -5546
rect 13932 -5648 13966 -5614
rect 13932 -5716 13966 -5682
rect 18290 -5580 18324 -5546
rect 18290 -5648 18324 -5614
rect 18290 -5716 18324 -5682
rect 856 -5784 890 -5750
rect 856 -5852 890 -5818
rect 5214 -5784 5248 -5750
rect 856 -5920 890 -5886
rect 856 -5988 890 -5954
rect 856 -6056 890 -6022
rect 856 -6124 890 -6090
rect 5214 -5852 5248 -5818
rect 9573 -5784 9607 -5750
rect 5214 -5920 5248 -5886
rect 5214 -5988 5248 -5954
rect 5214 -6056 5248 -6022
rect 5214 -6124 5248 -6090
rect 856 -6192 890 -6158
rect 856 -6260 890 -6226
rect 9573 -5852 9607 -5818
rect 13932 -5784 13966 -5750
rect 9573 -5920 9607 -5886
rect 9573 -5988 9607 -5954
rect 9573 -6056 9607 -6022
rect 9573 -6124 9607 -6090
rect 5214 -6192 5248 -6158
rect 856 -6328 890 -6294
rect 856 -6396 890 -6362
rect 856 -6464 890 -6430
rect 5214 -6260 5248 -6226
rect 13932 -5852 13966 -5818
rect 18290 -5784 18324 -5750
rect 13932 -5920 13966 -5886
rect 13932 -5988 13966 -5954
rect 13932 -6056 13966 -6022
rect 13932 -6124 13966 -6090
rect 9573 -6192 9607 -6158
rect 5214 -6328 5248 -6294
rect 5214 -6396 5248 -6362
rect 5214 -6464 5248 -6430
rect 9573 -6260 9607 -6226
rect 18290 -5852 18324 -5818
rect 18290 -5920 18324 -5886
rect 18290 -5988 18324 -5954
rect 18290 -6056 18324 -6022
rect 18290 -6124 18324 -6090
rect 13932 -6192 13966 -6158
rect 9573 -6328 9607 -6294
rect 9573 -6396 9607 -6362
rect 856 -6532 890 -6498
rect 856 -6600 890 -6566
rect 856 -6668 890 -6634
rect 856 -6804 890 -6702
rect 9573 -6464 9607 -6430
rect 13932 -6260 13966 -6226
rect 18290 -6192 18324 -6158
rect 13932 -6328 13966 -6294
rect 13932 -6396 13966 -6362
rect 5214 -6532 5248 -6498
rect 5214 -6600 5248 -6566
rect 5214 -6668 5248 -6634
rect 5214 -6804 5248 -6702
rect 13932 -6464 13966 -6430
rect 18290 -6260 18324 -6226
rect 18290 -6328 18324 -6294
rect 18290 -6396 18324 -6362
rect 9573 -6532 9607 -6498
rect 9573 -6600 9607 -6566
rect 9573 -6668 9607 -6634
rect 9573 -6804 9607 -6702
rect 18290 -6464 18324 -6430
rect 13932 -6532 13966 -6498
rect 13932 -6600 13966 -6566
rect 13932 -6668 13966 -6634
rect 13932 -6804 13966 -6702
rect 18290 -6532 18324 -6498
rect 18290 -6600 18324 -6566
rect 18290 -6668 18324 -6634
rect 18290 -6804 18324 -6702
rect 856 -6838 977 -6804
rect 1011 -6838 1045 -6804
rect 1079 -6838 1113 -6804
rect 1147 -6838 1181 -6804
rect 1215 -6838 1249 -6804
rect 1283 -6838 1317 -6804
rect 1351 -6838 1385 -6804
rect 1419 -6838 1453 -6804
rect 1487 -6838 1521 -6804
rect 1555 -6838 1589 -6804
rect 1623 -6838 1657 -6804
rect 1691 -6838 1725 -6804
rect 1759 -6838 1793 -6804
rect 1827 -6838 1861 -6804
rect 1895 -6838 1929 -6804
rect 1963 -6838 1997 -6804
rect 2031 -6838 2065 -6804
rect 2099 -6838 2133 -6804
rect 2167 -6838 2201 -6804
rect 2235 -6838 2269 -6804
rect 2303 -6838 2337 -6804
rect 2371 -6838 2405 -6804
rect 2439 -6838 2473 -6804
rect 2507 -6838 2541 -6804
rect 2575 -6838 2609 -6804
rect 2643 -6838 2677 -6804
rect 2711 -6838 2745 -6804
rect 2779 -6838 2813 -6804
rect 2847 -6838 2881 -6804
rect 2915 -6838 2949 -6804
rect 2983 -6838 3017 -6804
rect 3051 -6838 3085 -6804
rect 3119 -6838 3153 -6804
rect 3187 -6838 3221 -6804
rect 3255 -6838 3289 -6804
rect 3323 -6838 3357 -6804
rect 3391 -6838 3425 -6804
rect 3459 -6838 3493 -6804
rect 3527 -6838 3561 -6804
rect 3595 -6838 3629 -6804
rect 3663 -6838 3697 -6804
rect 3731 -6838 3765 -6804
rect 3799 -6838 3833 -6804
rect 3867 -6838 3901 -6804
rect 3935 -6838 3969 -6804
rect 4003 -6838 4037 -6804
rect 4071 -6838 4105 -6804
rect 4139 -6838 4173 -6804
rect 4207 -6838 4241 -6804
rect 4275 -6838 4309 -6804
rect 4343 -6838 4377 -6804
rect 4411 -6838 4445 -6804
rect 4479 -6838 4513 -6804
rect 4547 -6838 4581 -6804
rect 4615 -6838 4649 -6804
rect 4683 -6838 4717 -6804
rect 4751 -6838 4785 -6804
rect 4819 -6838 4853 -6804
rect 4887 -6838 4921 -6804
rect 4955 -6838 4989 -6804
rect 5023 -6838 5057 -6804
rect 5091 -6838 5372 -6804
rect 5406 -6838 5440 -6804
rect 5474 -6838 5508 -6804
rect 5542 -6838 5576 -6804
rect 5610 -6838 5644 -6804
rect 5678 -6838 5712 -6804
rect 5746 -6838 5780 -6804
rect 5814 -6838 5848 -6804
rect 5882 -6838 5916 -6804
rect 5950 -6838 5984 -6804
rect 6018 -6838 6052 -6804
rect 6086 -6838 6120 -6804
rect 6154 -6838 6188 -6804
rect 6222 -6838 6256 -6804
rect 6290 -6838 6324 -6804
rect 6358 -6838 6392 -6804
rect 6426 -6838 6460 -6804
rect 6494 -6838 6528 -6804
rect 6562 -6838 6596 -6804
rect 6630 -6838 6664 -6804
rect 6698 -6838 6732 -6804
rect 6766 -6838 6800 -6804
rect 6834 -6838 6868 -6804
rect 6902 -6838 6936 -6804
rect 6970 -6838 7004 -6804
rect 7038 -6838 7072 -6804
rect 7106 -6838 7140 -6804
rect 7174 -6838 7208 -6804
rect 7242 -6838 7276 -6804
rect 7310 -6838 7344 -6804
rect 7378 -6838 7412 -6804
rect 7446 -6838 7480 -6804
rect 7514 -6838 7548 -6804
rect 7582 -6838 7616 -6804
rect 7650 -6838 7684 -6804
rect 7718 -6838 7752 -6804
rect 7786 -6838 7820 -6804
rect 7854 -6838 7888 -6804
rect 7922 -6838 7956 -6804
rect 7990 -6838 8024 -6804
rect 8058 -6838 8092 -6804
rect 8126 -6838 8160 -6804
rect 8194 -6838 8228 -6804
rect 8262 -6838 8296 -6804
rect 8330 -6838 8364 -6804
rect 8398 -6838 8432 -6804
rect 8466 -6838 8500 -6804
rect 8534 -6838 8568 -6804
rect 8602 -6838 8636 -6804
rect 8670 -6838 8704 -6804
rect 8738 -6838 8772 -6804
rect 8806 -6838 8840 -6804
rect 8874 -6838 8908 -6804
rect 8942 -6838 8976 -6804
rect 9010 -6838 9044 -6804
rect 9078 -6838 9112 -6804
rect 9146 -6838 9180 -6804
rect 9214 -6838 9248 -6804
rect 9282 -6838 9316 -6804
rect 9350 -6838 9384 -6804
rect 9418 -6838 9452 -6804
rect 9486 -6838 9694 -6804
rect 9728 -6838 9762 -6804
rect 9796 -6838 9830 -6804
rect 9864 -6838 9898 -6804
rect 9932 -6838 9966 -6804
rect 10000 -6838 10034 -6804
rect 10068 -6838 10102 -6804
rect 10136 -6838 10170 -6804
rect 10204 -6838 10238 -6804
rect 10272 -6838 10306 -6804
rect 10340 -6838 10374 -6804
rect 10408 -6838 10442 -6804
rect 10476 -6838 10510 -6804
rect 10544 -6838 10578 -6804
rect 10612 -6838 10646 -6804
rect 10680 -6838 10714 -6804
rect 10748 -6838 10782 -6804
rect 10816 -6838 10850 -6804
rect 10884 -6838 10918 -6804
rect 10952 -6838 10986 -6804
rect 11020 -6838 11054 -6804
rect 11088 -6838 11122 -6804
rect 11156 -6838 11190 -6804
rect 11224 -6838 11258 -6804
rect 11292 -6838 11326 -6804
rect 11360 -6838 11394 -6804
rect 11428 -6838 11462 -6804
rect 11496 -6838 11530 -6804
rect 11564 -6838 11598 -6804
rect 11632 -6838 11666 -6804
rect 11700 -6838 11734 -6804
rect 11768 -6838 11802 -6804
rect 11836 -6838 11870 -6804
rect 11904 -6838 11938 -6804
rect 11972 -6838 12006 -6804
rect 12040 -6838 12074 -6804
rect 12108 -6838 12142 -6804
rect 12176 -6838 12210 -6804
rect 12244 -6838 12278 -6804
rect 12312 -6838 12346 -6804
rect 12380 -6838 12414 -6804
rect 12448 -6838 12482 -6804
rect 12516 -6838 12550 -6804
rect 12584 -6838 12618 -6804
rect 12652 -6838 12686 -6804
rect 12720 -6838 12754 -6804
rect 12788 -6838 12822 -6804
rect 12856 -6838 12890 -6804
rect 12924 -6838 12958 -6804
rect 12992 -6838 13026 -6804
rect 13060 -6838 13094 -6804
rect 13128 -6838 13162 -6804
rect 13196 -6838 13230 -6804
rect 13264 -6838 13298 -6804
rect 13332 -6838 13366 -6804
rect 13400 -6838 13434 -6804
rect 13468 -6838 13502 -6804
rect 13536 -6838 13570 -6804
rect 13604 -6838 13638 -6804
rect 13672 -6838 13706 -6804
rect 13740 -6838 13774 -6804
rect 13808 -6838 14089 -6804
rect 14123 -6838 14157 -6804
rect 14191 -6838 14225 -6804
rect 14259 -6838 14293 -6804
rect 14327 -6838 14361 -6804
rect 14395 -6838 14429 -6804
rect 14463 -6838 14497 -6804
rect 14531 -6838 14565 -6804
rect 14599 -6838 14633 -6804
rect 14667 -6838 14701 -6804
rect 14735 -6838 14769 -6804
rect 14803 -6838 14837 -6804
rect 14871 -6838 14905 -6804
rect 14939 -6838 14973 -6804
rect 15007 -6838 15041 -6804
rect 15075 -6838 15109 -6804
rect 15143 -6838 15177 -6804
rect 15211 -6838 15245 -6804
rect 15279 -6838 15313 -6804
rect 15347 -6838 15381 -6804
rect 15415 -6838 15449 -6804
rect 15483 -6838 15517 -6804
rect 15551 -6838 15585 -6804
rect 15619 -6838 15653 -6804
rect 15687 -6838 15721 -6804
rect 15755 -6838 15789 -6804
rect 15823 -6838 15857 -6804
rect 15891 -6838 15925 -6804
rect 15959 -6838 15993 -6804
rect 16027 -6838 16061 -6804
rect 16095 -6838 16129 -6804
rect 16163 -6838 16197 -6804
rect 16231 -6838 16265 -6804
rect 16299 -6838 16333 -6804
rect 16367 -6838 16401 -6804
rect 16435 -6838 16469 -6804
rect 16503 -6838 16537 -6804
rect 16571 -6838 16605 -6804
rect 16639 -6838 16673 -6804
rect 16707 -6838 16741 -6804
rect 16775 -6838 16809 -6804
rect 16843 -6838 16877 -6804
rect 16911 -6838 16945 -6804
rect 16979 -6838 17013 -6804
rect 17047 -6838 17081 -6804
rect 17115 -6838 17149 -6804
rect 17183 -6838 17217 -6804
rect 17251 -6838 17285 -6804
rect 17319 -6838 17353 -6804
rect 17387 -6838 17421 -6804
rect 17455 -6838 17489 -6804
rect 17523 -6838 17557 -6804
rect 17591 -6838 17625 -6804
rect 17659 -6838 17693 -6804
rect 17727 -6838 17761 -6804
rect 17795 -6838 17829 -6804
rect 17863 -6838 17897 -6804
rect 17931 -6838 17965 -6804
rect 17999 -6838 18033 -6804
rect 18067 -6838 18101 -6804
rect 18135 -6838 18169 -6804
rect 18203 -6838 18324 -6804
rect 856 -6940 890 -6838
rect 856 -7008 890 -6974
rect 856 -7076 890 -7042
rect 856 -7144 890 -7110
rect 5214 -6940 5248 -6838
rect 5214 -7008 5248 -6974
rect 5214 -7076 5248 -7042
rect 5214 -7144 5248 -7110
rect 856 -7212 890 -7178
rect 9573 -6940 9607 -6838
rect 9573 -7008 9607 -6974
rect 9573 -7076 9607 -7042
rect 9573 -7144 9607 -7110
rect 856 -7280 890 -7246
rect 856 -7348 890 -7314
rect 856 -7416 890 -7382
rect 5214 -7212 5248 -7178
rect 13932 -6940 13966 -6838
rect 13932 -7008 13966 -6974
rect 13932 -7076 13966 -7042
rect 13932 -7144 13966 -7110
rect 5214 -7280 5248 -7246
rect 5214 -7348 5248 -7314
rect 856 -7484 890 -7450
rect 5214 -7416 5248 -7382
rect 9573 -7212 9607 -7178
rect 18290 -6940 18324 -6838
rect 18290 -7008 18324 -6974
rect 18290 -7076 18324 -7042
rect 18290 -7144 18324 -7110
rect 9573 -7280 9607 -7246
rect 9573 -7348 9607 -7314
rect 5214 -7484 5248 -7450
rect 856 -7552 890 -7518
rect 856 -7620 890 -7586
rect 856 -7688 890 -7654
rect 856 -7756 890 -7722
rect 9573 -7416 9607 -7382
rect 13932 -7212 13966 -7178
rect 13932 -7280 13966 -7246
rect 13932 -7348 13966 -7314
rect 9573 -7484 9607 -7450
rect 5214 -7552 5248 -7518
rect 5214 -7620 5248 -7586
rect 5214 -7688 5248 -7654
rect 5214 -7756 5248 -7722
rect 13932 -7416 13966 -7382
rect 18290 -7212 18324 -7178
rect 18290 -7280 18324 -7246
rect 18290 -7348 18324 -7314
rect 13932 -7484 13966 -7450
rect 9573 -7552 9607 -7518
rect 9573 -7620 9607 -7586
rect 9573 -7688 9607 -7654
rect 9573 -7756 9607 -7722
rect 18290 -7416 18324 -7382
rect 18290 -7484 18324 -7450
rect 13932 -7552 13966 -7518
rect 13932 -7620 13966 -7586
rect 13932 -7688 13966 -7654
rect 13932 -7756 13966 -7722
rect 18290 -7552 18324 -7518
rect 18290 -7620 18324 -7586
rect 18290 -7688 18324 -7654
rect 18290 -7756 18324 -7722
rect 856 -7824 890 -7790
rect 856 -7892 890 -7858
rect 5214 -7824 5248 -7790
rect 856 -7960 890 -7926
rect 856 -8028 890 -7994
rect 856 -8096 890 -8062
rect 5214 -7892 5248 -7858
rect 9573 -7824 9607 -7790
rect 5214 -7960 5248 -7926
rect 5214 -8028 5248 -7994
rect 5214 -8096 5248 -8062
rect 9573 -7892 9607 -7858
rect 13932 -7824 13966 -7790
rect 9573 -7960 9607 -7926
rect 9573 -8028 9607 -7994
rect 856 -8164 890 -8130
rect 856 -8232 890 -8198
rect 856 -8300 890 -8266
rect 856 -8368 890 -8334
rect 9573 -8096 9607 -8062
rect 13932 -7892 13966 -7858
rect 18290 -7824 18324 -7790
rect 13932 -7960 13966 -7926
rect 13932 -8028 13966 -7994
rect 5214 -8164 5248 -8130
rect 5214 -8232 5248 -8198
rect 5214 -8300 5248 -8266
rect 5214 -8368 5248 -8334
rect 13932 -8096 13966 -8062
rect 18290 -7892 18324 -7858
rect 18290 -7960 18324 -7926
rect 18290 -8028 18324 -7994
rect 9573 -8164 9607 -8130
rect 9573 -8232 9607 -8198
rect 9573 -8300 9607 -8266
rect 9573 -8368 9607 -8334
rect 18290 -8096 18324 -8062
rect 13932 -8164 13966 -8130
rect 13932 -8232 13966 -8198
rect 13932 -8300 13966 -8266
rect 13932 -8368 13966 -8334
rect 18290 -8164 18324 -8130
rect 18290 -8232 18324 -8198
rect 18290 -8300 18324 -8266
rect 18290 -8368 18324 -8334
rect 856 -8436 977 -8402
rect 1011 -8436 1045 -8402
rect 1079 -8436 1113 -8402
rect 1147 -8436 1181 -8402
rect 1215 -8436 1249 -8402
rect 1283 -8436 1317 -8402
rect 1351 -8436 1385 -8402
rect 1419 -8436 1453 -8402
rect 1487 -8436 1521 -8402
rect 1555 -8436 1589 -8402
rect 1623 -8436 1657 -8402
rect 1691 -8436 1725 -8402
rect 1759 -8436 1793 -8402
rect 1827 -8436 1861 -8402
rect 1895 -8436 1929 -8402
rect 1963 -8436 1997 -8402
rect 2031 -8436 2065 -8402
rect 2099 -8436 2133 -8402
rect 2167 -8436 2201 -8402
rect 2235 -8436 2269 -8402
rect 2303 -8436 2337 -8402
rect 2371 -8436 2405 -8402
rect 2439 -8436 2473 -8402
rect 2507 -8436 2541 -8402
rect 2575 -8436 2609 -8402
rect 2643 -8436 2677 -8402
rect 2711 -8436 2745 -8402
rect 2779 -8436 2813 -8402
rect 2847 -8436 2881 -8402
rect 2915 -8436 2949 -8402
rect 2983 -8436 3017 -8402
rect 3051 -8436 3085 -8402
rect 3119 -8436 3153 -8402
rect 3187 -8436 3221 -8402
rect 3255 -8436 3289 -8402
rect 3323 -8436 3357 -8402
rect 3391 -8436 3425 -8402
rect 3459 -8436 3493 -8402
rect 3527 -8436 3561 -8402
rect 3595 -8436 3629 -8402
rect 3663 -8436 3697 -8402
rect 3731 -8436 3765 -8402
rect 3799 -8436 3833 -8402
rect 3867 -8436 3901 -8402
rect 3935 -8436 3969 -8402
rect 4003 -8436 4037 -8402
rect 4071 -8436 4105 -8402
rect 4139 -8436 4173 -8402
rect 4207 -8436 4241 -8402
rect 4275 -8436 4309 -8402
rect 4343 -8436 4377 -8402
rect 4411 -8436 4445 -8402
rect 4479 -8436 4513 -8402
rect 4547 -8436 4581 -8402
rect 4615 -8436 4649 -8402
rect 4683 -8436 4717 -8402
rect 4751 -8436 4785 -8402
rect 4819 -8436 4853 -8402
rect 4887 -8436 4921 -8402
rect 4955 -8436 4989 -8402
rect 5023 -8436 5057 -8402
rect 5091 -8436 5372 -8402
rect 5406 -8436 5440 -8402
rect 5474 -8436 5508 -8402
rect 5542 -8436 5576 -8402
rect 5610 -8436 5644 -8402
rect 5678 -8436 5712 -8402
rect 5746 -8436 5780 -8402
rect 5814 -8436 5848 -8402
rect 5882 -8436 5916 -8402
rect 5950 -8436 5984 -8402
rect 6018 -8436 6052 -8402
rect 6086 -8436 6120 -8402
rect 6154 -8436 6188 -8402
rect 6222 -8436 6256 -8402
rect 6290 -8436 6324 -8402
rect 6358 -8436 6392 -8402
rect 6426 -8436 6460 -8402
rect 6494 -8436 6528 -8402
rect 6562 -8436 6596 -8402
rect 6630 -8436 6664 -8402
rect 6698 -8436 6732 -8402
rect 6766 -8436 6800 -8402
rect 6834 -8436 6868 -8402
rect 6902 -8436 6936 -8402
rect 6970 -8436 7004 -8402
rect 7038 -8436 7072 -8402
rect 7106 -8436 7140 -8402
rect 7174 -8436 7208 -8402
rect 7242 -8436 7276 -8402
rect 7310 -8436 7344 -8402
rect 7378 -8436 7412 -8402
rect 7446 -8436 7480 -8402
rect 7514 -8436 7548 -8402
rect 7582 -8436 7616 -8402
rect 7650 -8436 7684 -8402
rect 7718 -8436 7752 -8402
rect 7786 -8436 7820 -8402
rect 7854 -8436 7888 -8402
rect 7922 -8436 7956 -8402
rect 7990 -8436 8024 -8402
rect 8058 -8436 8092 -8402
rect 8126 -8436 8160 -8402
rect 8194 -8436 8228 -8402
rect 8262 -8436 8296 -8402
rect 8330 -8436 8364 -8402
rect 8398 -8436 8432 -8402
rect 8466 -8436 8500 -8402
rect 8534 -8436 8568 -8402
rect 8602 -8436 8636 -8402
rect 8670 -8436 8704 -8402
rect 8738 -8436 8772 -8402
rect 8806 -8436 8840 -8402
rect 8874 -8436 8908 -8402
rect 8942 -8436 8976 -8402
rect 9010 -8436 9044 -8402
rect 9078 -8436 9112 -8402
rect 9146 -8436 9180 -8402
rect 9214 -8436 9248 -8402
rect 9282 -8436 9316 -8402
rect 9350 -8436 9384 -8402
rect 9418 -8436 9452 -8402
rect 9486 -8436 9694 -8402
rect 9728 -8436 9762 -8402
rect 9796 -8436 9830 -8402
rect 9864 -8436 9898 -8402
rect 9932 -8436 9966 -8402
rect 10000 -8436 10034 -8402
rect 10068 -8436 10102 -8402
rect 10136 -8436 10170 -8402
rect 10204 -8436 10238 -8402
rect 10272 -8436 10306 -8402
rect 10340 -8436 10374 -8402
rect 10408 -8436 10442 -8402
rect 10476 -8436 10510 -8402
rect 10544 -8436 10578 -8402
rect 10612 -8436 10646 -8402
rect 10680 -8436 10714 -8402
rect 10748 -8436 10782 -8402
rect 10816 -8436 10850 -8402
rect 10884 -8436 10918 -8402
rect 10952 -8436 10986 -8402
rect 11020 -8436 11054 -8402
rect 11088 -8436 11122 -8402
rect 11156 -8436 11190 -8402
rect 11224 -8436 11258 -8402
rect 11292 -8436 11326 -8402
rect 11360 -8436 11394 -8402
rect 11428 -8436 11462 -8402
rect 11496 -8436 11530 -8402
rect 11564 -8436 11598 -8402
rect 11632 -8436 11666 -8402
rect 11700 -8436 11734 -8402
rect 11768 -8436 11802 -8402
rect 11836 -8436 11870 -8402
rect 11904 -8436 11938 -8402
rect 11972 -8436 12006 -8402
rect 12040 -8436 12074 -8402
rect 12108 -8436 12142 -8402
rect 12176 -8436 12210 -8402
rect 12244 -8436 12278 -8402
rect 12312 -8436 12346 -8402
rect 12380 -8436 12414 -8402
rect 12448 -8436 12482 -8402
rect 12516 -8436 12550 -8402
rect 12584 -8436 12618 -8402
rect 12652 -8436 12686 -8402
rect 12720 -8436 12754 -8402
rect 12788 -8436 12822 -8402
rect 12856 -8436 12890 -8402
rect 12924 -8436 12958 -8402
rect 12992 -8436 13026 -8402
rect 13060 -8436 13094 -8402
rect 13128 -8436 13162 -8402
rect 13196 -8436 13230 -8402
rect 13264 -8436 13298 -8402
rect 13332 -8436 13366 -8402
rect 13400 -8436 13434 -8402
rect 13468 -8436 13502 -8402
rect 13536 -8436 13570 -8402
rect 13604 -8436 13638 -8402
rect 13672 -8436 13706 -8402
rect 13740 -8436 13774 -8402
rect 13808 -8436 14089 -8402
rect 14123 -8436 14157 -8402
rect 14191 -8436 14225 -8402
rect 14259 -8436 14293 -8402
rect 14327 -8436 14361 -8402
rect 14395 -8436 14429 -8402
rect 14463 -8436 14497 -8402
rect 14531 -8436 14565 -8402
rect 14599 -8436 14633 -8402
rect 14667 -8436 14701 -8402
rect 14735 -8436 14769 -8402
rect 14803 -8436 14837 -8402
rect 14871 -8436 14905 -8402
rect 14939 -8436 14973 -8402
rect 15007 -8436 15041 -8402
rect 15075 -8436 15109 -8402
rect 15143 -8436 15177 -8402
rect 15211 -8436 15245 -8402
rect 15279 -8436 15313 -8402
rect 15347 -8436 15381 -8402
rect 15415 -8436 15449 -8402
rect 15483 -8436 15517 -8402
rect 15551 -8436 15585 -8402
rect 15619 -8436 15653 -8402
rect 15687 -8436 15721 -8402
rect 15755 -8436 15789 -8402
rect 15823 -8436 15857 -8402
rect 15891 -8436 15925 -8402
rect 15959 -8436 15993 -8402
rect 16027 -8436 16061 -8402
rect 16095 -8436 16129 -8402
rect 16163 -8436 16197 -8402
rect 16231 -8436 16265 -8402
rect 16299 -8436 16333 -8402
rect 16367 -8436 16401 -8402
rect 16435 -8436 16469 -8402
rect 16503 -8436 16537 -8402
rect 16571 -8436 16605 -8402
rect 16639 -8436 16673 -8402
rect 16707 -8436 16741 -8402
rect 16775 -8436 16809 -8402
rect 16843 -8436 16877 -8402
rect 16911 -8436 16945 -8402
rect 16979 -8436 17013 -8402
rect 17047 -8436 17081 -8402
rect 17115 -8436 17149 -8402
rect 17183 -8436 17217 -8402
rect 17251 -8436 17285 -8402
rect 17319 -8436 17353 -8402
rect 17387 -8436 17421 -8402
rect 17455 -8436 17489 -8402
rect 17523 -8436 17557 -8402
rect 17591 -8436 17625 -8402
rect 17659 -8436 17693 -8402
rect 17727 -8436 17761 -8402
rect 17795 -8436 17829 -8402
rect 17863 -8436 17897 -8402
rect 17931 -8436 17965 -8402
rect 17999 -8436 18033 -8402
rect 18067 -8436 18101 -8402
rect 18135 -8436 18169 -8402
rect 18203 -8436 18324 -8402
rect 856 -8504 890 -8470
rect 856 -8572 890 -8538
rect 856 -8640 890 -8606
rect 856 -8708 890 -8674
rect 856 -8776 890 -8742
rect 5214 -8504 5248 -8470
rect 5214 -8572 5248 -8538
rect 5214 -8640 5248 -8606
rect 5214 -8708 5248 -8674
rect 5214 -8776 5248 -8742
rect 856 -8844 890 -8810
rect 9573 -8504 9607 -8470
rect 9573 -8572 9607 -8538
rect 9573 -8640 9607 -8606
rect 9573 -8708 9607 -8674
rect 9573 -8776 9607 -8742
rect 856 -8912 890 -8878
rect 856 -8980 890 -8946
rect 856 -9192 890 -9014
rect 5214 -8844 5248 -8810
rect 13932 -8504 13966 -8470
rect 13932 -8572 13966 -8538
rect 13932 -8640 13966 -8606
rect 13932 -8708 13966 -8674
rect 13932 -8776 13966 -8742
rect 5214 -8912 5248 -8878
rect 5214 -8980 5248 -8946
rect 5214 -9192 5248 -9014
rect 9573 -8844 9607 -8810
rect 18290 -8504 18324 -8470
rect 18290 -8572 18324 -8538
rect 18290 -8640 18324 -8606
rect 18290 -8708 18324 -8674
rect 18290 -8776 18324 -8742
rect 9573 -8912 9607 -8878
rect 9573 -8980 9607 -8946
rect 9573 -9192 9607 -9014
rect 13932 -8844 13966 -8810
rect 13932 -8912 13966 -8878
rect 13932 -8980 13966 -8946
rect 13932 -9192 13966 -9014
rect 18290 -8844 18324 -8810
rect 18290 -8912 18324 -8878
rect 18290 -8980 18324 -8946
rect 18290 -9192 18324 -9014
rect 856 -9226 977 -9192
rect 1011 -9226 1045 -9192
rect 1079 -9226 1113 -9192
rect 1147 -9226 1181 -9192
rect 1215 -9226 1249 -9192
rect 1283 -9226 1317 -9192
rect 1351 -9226 1385 -9192
rect 1419 -9226 1453 -9192
rect 1487 -9226 1521 -9192
rect 1555 -9226 1589 -9192
rect 1623 -9226 1657 -9192
rect 1691 -9226 1725 -9192
rect 1759 -9226 1793 -9192
rect 1827 -9226 1861 -9192
rect 1895 -9226 1929 -9192
rect 1963 -9226 1997 -9192
rect 2031 -9226 2065 -9192
rect 2099 -9226 2133 -9192
rect 2167 -9226 2201 -9192
rect 2235 -9226 2269 -9192
rect 2303 -9226 2337 -9192
rect 2371 -9226 2405 -9192
rect 2439 -9226 2473 -9192
rect 2507 -9226 2541 -9192
rect 2575 -9226 2609 -9192
rect 2643 -9226 2677 -9192
rect 2711 -9226 2745 -9192
rect 2779 -9226 2813 -9192
rect 2847 -9226 2881 -9192
rect 2915 -9226 2949 -9192
rect 2983 -9226 3017 -9192
rect 3051 -9226 3085 -9192
rect 3119 -9226 3153 -9192
rect 3187 -9226 3221 -9192
rect 3255 -9226 3289 -9192
rect 3323 -9226 3357 -9192
rect 3391 -9226 3425 -9192
rect 3459 -9226 3493 -9192
rect 3527 -9226 3561 -9192
rect 3595 -9226 3629 -9192
rect 3663 -9226 3697 -9192
rect 3731 -9226 3765 -9192
rect 3799 -9226 3833 -9192
rect 3867 -9226 3901 -9192
rect 3935 -9226 3969 -9192
rect 4003 -9226 4037 -9192
rect 4071 -9226 4105 -9192
rect 4139 -9226 4173 -9192
rect 4207 -9226 4241 -9192
rect 4275 -9226 4309 -9192
rect 4343 -9226 4377 -9192
rect 4411 -9226 4445 -9192
rect 4479 -9226 4513 -9192
rect 4547 -9226 4581 -9192
rect 4615 -9226 4649 -9192
rect 4683 -9226 4717 -9192
rect 4751 -9226 4785 -9192
rect 4819 -9226 4853 -9192
rect 4887 -9226 4921 -9192
rect 4955 -9226 4989 -9192
rect 5023 -9226 5057 -9192
rect 5091 -9226 5372 -9192
rect 5406 -9226 5440 -9192
rect 5474 -9226 5508 -9192
rect 5542 -9226 5576 -9192
rect 5610 -9226 5644 -9192
rect 5678 -9226 5712 -9192
rect 5746 -9226 5780 -9192
rect 5814 -9226 5848 -9192
rect 5882 -9226 5916 -9192
rect 5950 -9226 5984 -9192
rect 6018 -9226 6052 -9192
rect 6086 -9226 6120 -9192
rect 6154 -9226 6188 -9192
rect 6222 -9226 6256 -9192
rect 6290 -9226 6324 -9192
rect 6358 -9226 6392 -9192
rect 6426 -9226 6460 -9192
rect 6494 -9226 6528 -9192
rect 6562 -9226 6596 -9192
rect 6630 -9226 6664 -9192
rect 6698 -9226 6732 -9192
rect 6766 -9226 6800 -9192
rect 6834 -9226 6868 -9192
rect 6902 -9226 6936 -9192
rect 6970 -9226 7004 -9192
rect 7038 -9226 7072 -9192
rect 7106 -9226 7140 -9192
rect 7174 -9226 7208 -9192
rect 7242 -9226 7276 -9192
rect 7310 -9226 7344 -9192
rect 7378 -9226 7412 -9192
rect 7446 -9226 7480 -9192
rect 7514 -9226 7548 -9192
rect 7582 -9226 7616 -9192
rect 7650 -9226 7684 -9192
rect 7718 -9226 7752 -9192
rect 7786 -9226 7820 -9192
rect 7854 -9226 7888 -9192
rect 7922 -9226 7956 -9192
rect 7990 -9226 8024 -9192
rect 8058 -9226 8092 -9192
rect 8126 -9226 8160 -9192
rect 8194 -9226 8228 -9192
rect 8262 -9226 8296 -9192
rect 8330 -9226 8364 -9192
rect 8398 -9226 8432 -9192
rect 8466 -9226 8500 -9192
rect 8534 -9226 8568 -9192
rect 8602 -9226 8636 -9192
rect 8670 -9226 8704 -9192
rect 8738 -9226 8772 -9192
rect 8806 -9226 8840 -9192
rect 8874 -9226 8908 -9192
rect 8942 -9226 8976 -9192
rect 9010 -9226 9044 -9192
rect 9078 -9226 9112 -9192
rect 9146 -9226 9180 -9192
rect 9214 -9226 9248 -9192
rect 9282 -9226 9316 -9192
rect 9350 -9226 9384 -9192
rect 9418 -9226 9452 -9192
rect 9486 -9226 9694 -9192
rect 9728 -9226 9762 -9192
rect 9796 -9226 9830 -9192
rect 9864 -9226 9898 -9192
rect 9932 -9226 9966 -9192
rect 10000 -9226 10034 -9192
rect 10068 -9226 10102 -9192
rect 10136 -9226 10170 -9192
rect 10204 -9226 10238 -9192
rect 10272 -9226 10306 -9192
rect 10340 -9226 10374 -9192
rect 10408 -9226 10442 -9192
rect 10476 -9226 10510 -9192
rect 10544 -9226 10578 -9192
rect 10612 -9226 10646 -9192
rect 10680 -9226 10714 -9192
rect 10748 -9226 10782 -9192
rect 10816 -9226 10850 -9192
rect 10884 -9226 10918 -9192
rect 10952 -9226 10986 -9192
rect 11020 -9226 11054 -9192
rect 11088 -9226 11122 -9192
rect 11156 -9226 11190 -9192
rect 11224 -9226 11258 -9192
rect 11292 -9226 11326 -9192
rect 11360 -9226 11394 -9192
rect 11428 -9226 11462 -9192
rect 11496 -9226 11530 -9192
rect 11564 -9226 11598 -9192
rect 11632 -9226 11666 -9192
rect 11700 -9226 11734 -9192
rect 11768 -9226 11802 -9192
rect 11836 -9226 11870 -9192
rect 11904 -9226 11938 -9192
rect 11972 -9226 12006 -9192
rect 12040 -9226 12074 -9192
rect 12108 -9226 12142 -9192
rect 12176 -9226 12210 -9192
rect 12244 -9226 12278 -9192
rect 12312 -9226 12346 -9192
rect 12380 -9226 12414 -9192
rect 12448 -9226 12482 -9192
rect 12516 -9226 12550 -9192
rect 12584 -9226 12618 -9192
rect 12652 -9226 12686 -9192
rect 12720 -9226 12754 -9192
rect 12788 -9226 12822 -9192
rect 12856 -9226 12890 -9192
rect 12924 -9226 12958 -9192
rect 12992 -9226 13026 -9192
rect 13060 -9226 13094 -9192
rect 13128 -9226 13162 -9192
rect 13196 -9226 13230 -9192
rect 13264 -9226 13298 -9192
rect 13332 -9226 13366 -9192
rect 13400 -9226 13434 -9192
rect 13468 -9226 13502 -9192
rect 13536 -9226 13570 -9192
rect 13604 -9226 13638 -9192
rect 13672 -9226 13706 -9192
rect 13740 -9226 13774 -9192
rect 13808 -9226 14089 -9192
rect 14123 -9226 14157 -9192
rect 14191 -9226 14225 -9192
rect 14259 -9226 14293 -9192
rect 14327 -9226 14361 -9192
rect 14395 -9226 14429 -9192
rect 14463 -9226 14497 -9192
rect 14531 -9226 14565 -9192
rect 14599 -9226 14633 -9192
rect 14667 -9226 14701 -9192
rect 14735 -9226 14769 -9192
rect 14803 -9226 14837 -9192
rect 14871 -9226 14905 -9192
rect 14939 -9226 14973 -9192
rect 15007 -9226 15041 -9192
rect 15075 -9226 15109 -9192
rect 15143 -9226 15177 -9192
rect 15211 -9226 15245 -9192
rect 15279 -9226 15313 -9192
rect 15347 -9226 15381 -9192
rect 15415 -9226 15449 -9192
rect 15483 -9226 15517 -9192
rect 15551 -9226 15585 -9192
rect 15619 -9226 15653 -9192
rect 15687 -9226 15721 -9192
rect 15755 -9226 15789 -9192
rect 15823 -9226 15857 -9192
rect 15891 -9226 15925 -9192
rect 15959 -9226 15993 -9192
rect 16027 -9226 16061 -9192
rect 16095 -9226 16129 -9192
rect 16163 -9226 16197 -9192
rect 16231 -9226 16265 -9192
rect 16299 -9226 16333 -9192
rect 16367 -9226 16401 -9192
rect 16435 -9226 16469 -9192
rect 16503 -9226 16537 -9192
rect 16571 -9226 16605 -9192
rect 16639 -9226 16673 -9192
rect 16707 -9226 16741 -9192
rect 16775 -9226 16809 -9192
rect 16843 -9226 16877 -9192
rect 16911 -9226 16945 -9192
rect 16979 -9226 17013 -9192
rect 17047 -9226 17081 -9192
rect 17115 -9226 17149 -9192
rect 17183 -9226 17217 -9192
rect 17251 -9226 17285 -9192
rect 17319 -9226 17353 -9192
rect 17387 -9226 17421 -9192
rect 17455 -9226 17489 -9192
rect 17523 -9226 17557 -9192
rect 17591 -9226 17625 -9192
rect 17659 -9226 17693 -9192
rect 17727 -9226 17761 -9192
rect 17795 -9226 17829 -9192
rect 17863 -9226 17897 -9192
rect 17931 -9226 17965 -9192
rect 17999 -9226 18033 -9192
rect 18067 -9226 18101 -9192
rect 18135 -9226 18169 -9192
rect 18203 -9226 18324 -9192
<< nsubdiffcont >>
rect 977 429 1011 463
rect 1045 429 1079 463
rect 1113 429 1147 463
rect 1181 429 1215 463
rect 1249 429 1283 463
rect 1317 429 1351 463
rect 1385 429 1419 463
rect 1453 429 1487 463
rect 1521 429 1555 463
rect 1589 429 1623 463
rect 1657 429 1691 463
rect 1725 429 1759 463
rect 1793 429 1827 463
rect 1861 429 1895 463
rect 1929 429 1963 463
rect 1997 429 2031 463
rect 2065 429 2099 463
rect 2133 429 2167 463
rect 2201 429 2235 463
rect 2269 429 2303 463
rect 2337 429 2371 463
rect 2405 429 2439 463
rect 2473 429 2507 463
rect 2541 429 2575 463
rect 2609 429 2643 463
rect 2677 429 2711 463
rect 2745 429 2779 463
rect 2813 429 2847 463
rect 2881 429 2915 463
rect 2949 429 2983 463
rect 3017 429 3051 463
rect 3085 429 3119 463
rect 3153 429 3187 463
rect 3221 429 3255 463
rect 3289 429 3323 463
rect 3357 429 3391 463
rect 3425 429 3459 463
rect 3493 429 3527 463
rect 3561 429 3595 463
rect 3629 429 3663 463
rect 3697 429 3731 463
rect 3765 429 3799 463
rect 3833 429 3867 463
rect 3901 429 3935 463
rect 3969 429 4003 463
rect 4037 429 4071 463
rect 4105 429 4139 463
rect 4173 429 4207 463
rect 4241 429 4275 463
rect 4309 429 4343 463
rect 4377 429 4411 463
rect 4445 429 4479 463
rect 4513 429 4547 463
rect 4581 429 4615 463
rect 4649 429 4683 463
rect 4717 429 4751 463
rect 4785 429 4819 463
rect 4853 429 4887 463
rect 4921 429 4955 463
rect 4989 429 5023 463
rect 5057 429 5091 463
rect 5372 429 5406 463
rect 5440 429 5474 463
rect 5508 429 5542 463
rect 5576 429 5610 463
rect 5644 429 5678 463
rect 5712 429 5746 463
rect 5780 429 5814 463
rect 5848 429 5882 463
rect 5916 429 5950 463
rect 5984 429 6018 463
rect 6052 429 6086 463
rect 6120 429 6154 463
rect 6188 429 6222 463
rect 6256 429 6290 463
rect 6324 429 6358 463
rect 6392 429 6426 463
rect 6460 429 6494 463
rect 6528 429 6562 463
rect 6596 429 6630 463
rect 6664 429 6698 463
rect 6732 429 6766 463
rect 6800 429 6834 463
rect 6868 429 6902 463
rect 6936 429 6970 463
rect 7004 429 7038 463
rect 7072 429 7106 463
rect 7140 429 7174 463
rect 7208 429 7242 463
rect 7276 429 7310 463
rect 7344 429 7378 463
rect 7412 429 7446 463
rect 7480 429 7514 463
rect 7548 429 7582 463
rect 7616 429 7650 463
rect 7684 429 7718 463
rect 7752 429 7786 463
rect 7820 429 7854 463
rect 7888 429 7922 463
rect 7956 429 7990 463
rect 8024 429 8058 463
rect 8092 429 8126 463
rect 8160 429 8194 463
rect 8228 429 8262 463
rect 8296 429 8330 463
rect 8364 429 8398 463
rect 8432 429 8466 463
rect 8500 429 8534 463
rect 8568 429 8602 463
rect 8636 429 8670 463
rect 8704 429 8738 463
rect 8772 429 8806 463
rect 8840 429 8874 463
rect 8908 429 8942 463
rect 8976 429 9010 463
rect 9044 429 9078 463
rect 9112 429 9146 463
rect 9180 429 9214 463
rect 9248 429 9282 463
rect 9316 429 9350 463
rect 9384 429 9418 463
rect 9452 429 9486 463
rect 9694 429 9728 463
rect 9762 429 9796 463
rect 9830 429 9864 463
rect 9898 429 9932 463
rect 9966 429 10000 463
rect 10034 429 10068 463
rect 10102 429 10136 463
rect 10170 429 10204 463
rect 10238 429 10272 463
rect 10306 429 10340 463
rect 10374 429 10408 463
rect 10442 429 10476 463
rect 10510 429 10544 463
rect 10578 429 10612 463
rect 10646 429 10680 463
rect 10714 429 10748 463
rect 10782 429 10816 463
rect 10850 429 10884 463
rect 10918 429 10952 463
rect 10986 429 11020 463
rect 11054 429 11088 463
rect 11122 429 11156 463
rect 11190 429 11224 463
rect 11258 429 11292 463
rect 11326 429 11360 463
rect 11394 429 11428 463
rect 11462 429 11496 463
rect 11530 429 11564 463
rect 11598 429 11632 463
rect 11666 429 11700 463
rect 11734 429 11768 463
rect 11802 429 11836 463
rect 11870 429 11904 463
rect 11938 429 11972 463
rect 12006 429 12040 463
rect 12074 429 12108 463
rect 12142 429 12176 463
rect 12210 429 12244 463
rect 12278 429 12312 463
rect 12346 429 12380 463
rect 12414 429 12448 463
rect 12482 429 12516 463
rect 12550 429 12584 463
rect 12618 429 12652 463
rect 12686 429 12720 463
rect 12754 429 12788 463
rect 12822 429 12856 463
rect 12890 429 12924 463
rect 12958 429 12992 463
rect 13026 429 13060 463
rect 13094 429 13128 463
rect 13162 429 13196 463
rect 13230 429 13264 463
rect 13298 429 13332 463
rect 13366 429 13400 463
rect 13434 429 13468 463
rect 13502 429 13536 463
rect 13570 429 13604 463
rect 13638 429 13672 463
rect 13706 429 13740 463
rect 13774 429 13808 463
rect 14089 429 14123 463
rect 14157 429 14191 463
rect 14225 429 14259 463
rect 14293 429 14327 463
rect 14361 429 14395 463
rect 14429 429 14463 463
rect 14497 429 14531 463
rect 14565 429 14599 463
rect 14633 429 14667 463
rect 14701 429 14735 463
rect 14769 429 14803 463
rect 14837 429 14871 463
rect 14905 429 14939 463
rect 14973 429 15007 463
rect 15041 429 15075 463
rect 15109 429 15143 463
rect 15177 429 15211 463
rect 15245 429 15279 463
rect 15313 429 15347 463
rect 15381 429 15415 463
rect 15449 429 15483 463
rect 15517 429 15551 463
rect 15585 429 15619 463
rect 15653 429 15687 463
rect 15721 429 15755 463
rect 15789 429 15823 463
rect 15857 429 15891 463
rect 15925 429 15959 463
rect 15993 429 16027 463
rect 16061 429 16095 463
rect 16129 429 16163 463
rect 16197 429 16231 463
rect 16265 429 16299 463
rect 16333 429 16367 463
rect 16401 429 16435 463
rect 16469 429 16503 463
rect 16537 429 16571 463
rect 16605 429 16639 463
rect 16673 429 16707 463
rect 16741 429 16775 463
rect 16809 429 16843 463
rect 16877 429 16911 463
rect 16945 429 16979 463
rect 17013 429 17047 463
rect 17081 429 17115 463
rect 17149 429 17183 463
rect 17217 429 17251 463
rect 17285 429 17319 463
rect 17353 429 17387 463
rect 17421 429 17455 463
rect 17489 429 17523 463
rect 17557 429 17591 463
rect 17625 429 17659 463
rect 17693 429 17727 463
rect 17761 429 17795 463
rect 17829 429 17863 463
rect 17897 429 17931 463
rect 17965 429 17999 463
rect 18033 429 18067 463
rect 18101 429 18135 463
rect 18169 429 18203 463
rect 856 216 890 250
rect 856 148 890 182
rect 856 80 890 114
rect 5214 216 5248 250
rect 5214 148 5248 182
rect 5214 80 5248 114
rect 856 12 890 46
rect 9573 216 9607 250
rect 9573 148 9607 182
rect 9573 80 9607 114
rect 856 -56 890 -22
rect 856 -124 890 -90
rect 856 -192 890 -158
rect 856 -260 890 -226
rect 856 -328 890 -294
rect 5214 12 5248 46
rect 13932 216 13966 250
rect 13932 148 13966 182
rect 13932 80 13966 114
rect 5214 -56 5248 -22
rect 5214 -124 5248 -90
rect 5214 -192 5248 -158
rect 5214 -260 5248 -226
rect 5214 -328 5248 -294
rect 9573 12 9607 46
rect 18290 216 18324 250
rect 18290 148 18324 182
rect 18290 80 18324 114
rect 9573 -56 9607 -22
rect 9573 -124 9607 -90
rect 9573 -192 9607 -158
rect 9573 -260 9607 -226
rect 9573 -328 9607 -294
rect 13932 12 13966 46
rect 13932 -56 13966 -22
rect 13932 -124 13966 -90
rect 13932 -192 13966 -158
rect 13932 -260 13966 -226
rect 13932 -328 13966 -294
rect 18290 12 18324 46
rect 18290 -56 18324 -22
rect 18290 -124 18324 -90
rect 18290 -192 18324 -158
rect 18290 -260 18324 -226
rect 18290 -328 18324 -294
rect 977 -362 1011 -328
rect 1045 -362 1079 -328
rect 1113 -362 1147 -328
rect 1181 -362 1215 -328
rect 1249 -362 1283 -328
rect 1317 -362 1351 -328
rect 1385 -362 1419 -328
rect 1453 -362 1487 -328
rect 1521 -362 1555 -328
rect 1589 -362 1623 -328
rect 1657 -362 1691 -328
rect 1725 -362 1759 -328
rect 1793 -362 1827 -328
rect 1861 -362 1895 -328
rect 1929 -362 1963 -328
rect 1997 -362 2031 -328
rect 2065 -362 2099 -328
rect 2133 -362 2167 -328
rect 2201 -362 2235 -328
rect 2269 -362 2303 -328
rect 2337 -362 2371 -328
rect 2405 -362 2439 -328
rect 2473 -362 2507 -328
rect 2541 -362 2575 -328
rect 2609 -362 2643 -328
rect 2677 -362 2711 -328
rect 2745 -362 2779 -328
rect 2813 -362 2847 -328
rect 2881 -362 2915 -328
rect 2949 -362 2983 -328
rect 3017 -362 3051 -328
rect 3085 -362 3119 -328
rect 3153 -362 3187 -328
rect 3221 -362 3255 -328
rect 3289 -362 3323 -328
rect 3357 -362 3391 -328
rect 3425 -362 3459 -328
rect 3493 -362 3527 -328
rect 3561 -362 3595 -328
rect 3629 -362 3663 -328
rect 3697 -362 3731 -328
rect 3765 -362 3799 -328
rect 3833 -362 3867 -328
rect 3901 -362 3935 -328
rect 3969 -362 4003 -328
rect 4037 -362 4071 -328
rect 4105 -362 4139 -328
rect 4173 -362 4207 -328
rect 4241 -362 4275 -328
rect 4309 -362 4343 -328
rect 4377 -362 4411 -328
rect 4445 -362 4479 -328
rect 4513 -362 4547 -328
rect 4581 -362 4615 -328
rect 4649 -362 4683 -328
rect 4717 -362 4751 -328
rect 4785 -362 4819 -328
rect 4853 -362 4887 -328
rect 4921 -362 4955 -328
rect 4989 -362 5023 -328
rect 5057 -362 5091 -328
rect 5372 -362 5406 -328
rect 5440 -362 5474 -328
rect 5508 -362 5542 -328
rect 5576 -362 5610 -328
rect 5644 -362 5678 -328
rect 5712 -362 5746 -328
rect 5780 -362 5814 -328
rect 5848 -362 5882 -328
rect 5916 -362 5950 -328
rect 5984 -362 6018 -328
rect 6052 -362 6086 -328
rect 6120 -362 6154 -328
rect 6188 -362 6222 -328
rect 6256 -362 6290 -328
rect 6324 -362 6358 -328
rect 6392 -362 6426 -328
rect 6460 -362 6494 -328
rect 6528 -362 6562 -328
rect 6596 -362 6630 -328
rect 6664 -362 6698 -328
rect 6732 -362 6766 -328
rect 6800 -362 6834 -328
rect 6868 -362 6902 -328
rect 6936 -362 6970 -328
rect 7004 -362 7038 -328
rect 7072 -362 7106 -328
rect 7140 -362 7174 -328
rect 7208 -362 7242 -328
rect 7276 -362 7310 -328
rect 7344 -362 7378 -328
rect 7412 -362 7446 -328
rect 7480 -362 7514 -328
rect 7548 -362 7582 -328
rect 7616 -362 7650 -328
rect 7684 -362 7718 -328
rect 7752 -362 7786 -328
rect 7820 -362 7854 -328
rect 7888 -362 7922 -328
rect 7956 -362 7990 -328
rect 8024 -362 8058 -328
rect 8092 -362 8126 -328
rect 8160 -362 8194 -328
rect 8228 -362 8262 -328
rect 8296 -362 8330 -328
rect 8364 -362 8398 -328
rect 8432 -362 8466 -328
rect 8500 -362 8534 -328
rect 8568 -362 8602 -328
rect 8636 -362 8670 -328
rect 8704 -362 8738 -328
rect 8772 -362 8806 -328
rect 8840 -362 8874 -328
rect 8908 -362 8942 -328
rect 8976 -362 9010 -328
rect 9044 -362 9078 -328
rect 9112 -362 9146 -328
rect 9180 -362 9214 -328
rect 9248 -362 9282 -328
rect 9316 -362 9350 -328
rect 9384 -362 9418 -328
rect 9452 -362 9486 -328
rect 9694 -362 9728 -328
rect 9762 -362 9796 -328
rect 9830 -362 9864 -328
rect 9898 -362 9932 -328
rect 9966 -362 10000 -328
rect 10034 -362 10068 -328
rect 10102 -362 10136 -328
rect 10170 -362 10204 -328
rect 10238 -362 10272 -328
rect 10306 -362 10340 -328
rect 10374 -362 10408 -328
rect 10442 -362 10476 -328
rect 10510 -362 10544 -328
rect 10578 -362 10612 -328
rect 10646 -362 10680 -328
rect 10714 -362 10748 -328
rect 10782 -362 10816 -328
rect 10850 -362 10884 -328
rect 10918 -362 10952 -328
rect 10986 -362 11020 -328
rect 11054 -362 11088 -328
rect 11122 -362 11156 -328
rect 11190 -362 11224 -328
rect 11258 -362 11292 -328
rect 11326 -362 11360 -328
rect 11394 -362 11428 -328
rect 11462 -362 11496 -328
rect 11530 -362 11564 -328
rect 11598 -362 11632 -328
rect 11666 -362 11700 -328
rect 11734 -362 11768 -328
rect 11802 -362 11836 -328
rect 11870 -362 11904 -328
rect 11938 -362 11972 -328
rect 12006 -362 12040 -328
rect 12074 -362 12108 -328
rect 12142 -362 12176 -328
rect 12210 -362 12244 -328
rect 12278 -362 12312 -328
rect 12346 -362 12380 -328
rect 12414 -362 12448 -328
rect 12482 -362 12516 -328
rect 12550 -362 12584 -328
rect 12618 -362 12652 -328
rect 12686 -362 12720 -328
rect 12754 -362 12788 -328
rect 12822 -362 12856 -328
rect 12890 -362 12924 -328
rect 12958 -362 12992 -328
rect 13026 -362 13060 -328
rect 13094 -362 13128 -328
rect 13162 -362 13196 -328
rect 13230 -362 13264 -328
rect 13298 -362 13332 -328
rect 13366 -362 13400 -328
rect 13434 -362 13468 -328
rect 13502 -362 13536 -328
rect 13570 -362 13604 -328
rect 13638 -362 13672 -328
rect 13706 -362 13740 -328
rect 13774 -362 13808 -328
rect 14089 -362 14123 -328
rect 14157 -362 14191 -328
rect 14225 -362 14259 -328
rect 14293 -362 14327 -328
rect 14361 -362 14395 -328
rect 14429 -362 14463 -328
rect 14497 -362 14531 -328
rect 14565 -362 14599 -328
rect 14633 -362 14667 -328
rect 14701 -362 14735 -328
rect 14769 -362 14803 -328
rect 14837 -362 14871 -328
rect 14905 -362 14939 -328
rect 14973 -362 15007 -328
rect 15041 -362 15075 -328
rect 15109 -362 15143 -328
rect 15177 -362 15211 -328
rect 15245 -362 15279 -328
rect 15313 -362 15347 -328
rect 15381 -362 15415 -328
rect 15449 -362 15483 -328
rect 15517 -362 15551 -328
rect 15585 -362 15619 -328
rect 15653 -362 15687 -328
rect 15721 -362 15755 -328
rect 15789 -362 15823 -328
rect 15857 -362 15891 -328
rect 15925 -362 15959 -328
rect 15993 -362 16027 -328
rect 16061 -362 16095 -328
rect 16129 -362 16163 -328
rect 16197 -362 16231 -328
rect 16265 -362 16299 -328
rect 16333 -362 16367 -328
rect 16401 -362 16435 -328
rect 16469 -362 16503 -328
rect 16537 -362 16571 -328
rect 16605 -362 16639 -328
rect 16673 -362 16707 -328
rect 16741 -362 16775 -328
rect 16809 -362 16843 -328
rect 16877 -362 16911 -328
rect 16945 -362 16979 -328
rect 17013 -362 17047 -328
rect 17081 -362 17115 -328
rect 17149 -362 17183 -328
rect 17217 -362 17251 -328
rect 17285 -362 17319 -328
rect 17353 -362 17387 -328
rect 17421 -362 17455 -328
rect 17489 -362 17523 -328
rect 17557 -362 17591 -328
rect 17625 -362 17659 -328
rect 17693 -362 17727 -328
rect 17761 -362 17795 -328
rect 17829 -362 17863 -328
rect 17897 -362 17931 -328
rect 17965 -362 17999 -328
rect 18033 -362 18067 -328
rect 18101 -362 18135 -328
rect 18169 -362 18203 -328
rect 856 -396 890 -362
rect 856 -464 890 -430
rect 856 -532 890 -498
rect 856 -600 890 -566
rect 856 -668 890 -634
rect 5214 -396 5248 -362
rect 5214 -464 5248 -430
rect 5214 -532 5248 -498
rect 5214 -600 5248 -566
rect 5214 -668 5248 -634
rect 9573 -396 9607 -362
rect 9573 -464 9607 -430
rect 9573 -532 9607 -498
rect 9573 -600 9607 -566
rect 856 -736 890 -702
rect 856 -804 890 -770
rect 856 -872 890 -838
rect 9573 -668 9607 -634
rect 13932 -396 13966 -362
rect 13932 -464 13966 -430
rect 13932 -532 13966 -498
rect 13932 -600 13966 -566
rect 5214 -736 5248 -702
rect 5214 -804 5248 -770
rect 5214 -872 5248 -838
rect 856 -940 890 -906
rect 13932 -668 13966 -634
rect 18290 -396 18324 -362
rect 18290 -464 18324 -430
rect 18290 -532 18324 -498
rect 18290 -600 18324 -566
rect 9573 -736 9607 -702
rect 9573 -804 9607 -770
rect 9573 -872 9607 -838
rect 5214 -940 5248 -906
rect 856 -1008 890 -974
rect 856 -1076 890 -1042
rect 856 -1144 890 -1110
rect 856 -1212 890 -1178
rect 856 -1280 890 -1246
rect 18290 -668 18324 -634
rect 13932 -736 13966 -702
rect 13932 -804 13966 -770
rect 13932 -872 13966 -838
rect 9573 -940 9607 -906
rect 5214 -1008 5248 -974
rect 5214 -1076 5248 -1042
rect 5214 -1144 5248 -1110
rect 5214 -1212 5248 -1178
rect 856 -1348 890 -1314
rect 5214 -1280 5248 -1246
rect 18290 -736 18324 -702
rect 18290 -804 18324 -770
rect 18290 -872 18324 -838
rect 13932 -940 13966 -906
rect 9573 -1008 9607 -974
rect 9573 -1076 9607 -1042
rect 9573 -1144 9607 -1110
rect 9573 -1212 9607 -1178
rect 5214 -1348 5248 -1314
rect 856 -1416 890 -1382
rect 856 -1484 890 -1450
rect 856 -1552 890 -1518
rect 9573 -1280 9607 -1246
rect 18290 -940 18324 -906
rect 13932 -1008 13966 -974
rect 13932 -1076 13966 -1042
rect 13932 -1144 13966 -1110
rect 13932 -1212 13966 -1178
rect 9573 -1348 9607 -1314
rect 5214 -1416 5248 -1382
rect 5214 -1484 5248 -1450
rect 5214 -1552 5248 -1518
rect 856 -1620 890 -1586
rect 13932 -1280 13966 -1246
rect 18290 -1008 18324 -974
rect 18290 -1076 18324 -1042
rect 18290 -1144 18324 -1110
rect 18290 -1212 18324 -1178
rect 13932 -1348 13966 -1314
rect 9573 -1416 9607 -1382
rect 9573 -1484 9607 -1450
rect 9573 -1552 9607 -1518
rect 856 -1688 890 -1654
rect 856 -1756 890 -1722
rect 856 -1824 890 -1790
rect 5214 -1620 5248 -1586
rect 18290 -1280 18324 -1246
rect 18290 -1348 18324 -1314
rect 13932 -1416 13966 -1382
rect 13932 -1484 13966 -1450
rect 13932 -1552 13966 -1518
rect 5214 -1688 5248 -1654
rect 5214 -1756 5248 -1722
rect 5214 -1824 5248 -1790
rect 9573 -1620 9607 -1586
rect 18290 -1416 18324 -1382
rect 18290 -1484 18324 -1450
rect 18290 -1552 18324 -1518
rect 9573 -1688 9607 -1654
rect 9573 -1756 9607 -1722
rect 9573 -1824 9607 -1790
rect 13932 -1620 13966 -1586
rect 13932 -1688 13966 -1654
rect 13932 -1756 13966 -1722
rect 13932 -1824 13966 -1790
rect 18290 -1620 18324 -1586
rect 18290 -1688 18324 -1654
rect 18290 -1756 18324 -1722
rect 18290 -1824 18324 -1790
rect 977 -1960 1011 -1926
rect 1045 -1960 1079 -1926
rect 1113 -1960 1147 -1926
rect 1181 -1960 1215 -1926
rect 1249 -1960 1283 -1926
rect 1317 -1960 1351 -1926
rect 1385 -1960 1419 -1926
rect 1453 -1960 1487 -1926
rect 1521 -1960 1555 -1926
rect 1589 -1960 1623 -1926
rect 1657 -1960 1691 -1926
rect 1725 -1960 1759 -1926
rect 1793 -1960 1827 -1926
rect 1861 -1960 1895 -1926
rect 1929 -1960 1963 -1926
rect 1997 -1960 2031 -1926
rect 2065 -1960 2099 -1926
rect 2133 -1960 2167 -1926
rect 2201 -1960 2235 -1926
rect 2269 -1960 2303 -1926
rect 2337 -1960 2371 -1926
rect 2405 -1960 2439 -1926
rect 2473 -1960 2507 -1926
rect 2541 -1960 2575 -1926
rect 2609 -1960 2643 -1926
rect 2677 -1960 2711 -1926
rect 2745 -1960 2779 -1926
rect 2813 -1960 2847 -1926
rect 2881 -1960 2915 -1926
rect 2949 -1960 2983 -1926
rect 3017 -1960 3051 -1926
rect 3085 -1960 3119 -1926
rect 3153 -1960 3187 -1926
rect 3221 -1960 3255 -1926
rect 3289 -1960 3323 -1926
rect 3357 -1960 3391 -1926
rect 3425 -1960 3459 -1926
rect 3493 -1960 3527 -1926
rect 3561 -1960 3595 -1926
rect 3629 -1960 3663 -1926
rect 3697 -1960 3731 -1926
rect 3765 -1960 3799 -1926
rect 3833 -1960 3867 -1926
rect 3901 -1960 3935 -1926
rect 3969 -1960 4003 -1926
rect 4037 -1960 4071 -1926
rect 4105 -1960 4139 -1926
rect 4173 -1960 4207 -1926
rect 4241 -1960 4275 -1926
rect 4309 -1960 4343 -1926
rect 4377 -1960 4411 -1926
rect 4445 -1960 4479 -1926
rect 4513 -1960 4547 -1926
rect 4581 -1960 4615 -1926
rect 4649 -1960 4683 -1926
rect 4717 -1960 4751 -1926
rect 4785 -1960 4819 -1926
rect 4853 -1960 4887 -1926
rect 4921 -1960 4955 -1926
rect 4989 -1960 5023 -1926
rect 5057 -1960 5091 -1926
rect 5372 -1960 5406 -1926
rect 5440 -1960 5474 -1926
rect 5508 -1960 5542 -1926
rect 5576 -1960 5610 -1926
rect 5644 -1960 5678 -1926
rect 5712 -1960 5746 -1926
rect 5780 -1960 5814 -1926
rect 5848 -1960 5882 -1926
rect 5916 -1960 5950 -1926
rect 5984 -1960 6018 -1926
rect 6052 -1960 6086 -1926
rect 6120 -1960 6154 -1926
rect 6188 -1960 6222 -1926
rect 6256 -1960 6290 -1926
rect 6324 -1960 6358 -1926
rect 6392 -1960 6426 -1926
rect 6460 -1960 6494 -1926
rect 6528 -1960 6562 -1926
rect 6596 -1960 6630 -1926
rect 6664 -1960 6698 -1926
rect 6732 -1960 6766 -1926
rect 6800 -1960 6834 -1926
rect 6868 -1960 6902 -1926
rect 6936 -1960 6970 -1926
rect 7004 -1960 7038 -1926
rect 7072 -1960 7106 -1926
rect 7140 -1960 7174 -1926
rect 7208 -1960 7242 -1926
rect 7276 -1960 7310 -1926
rect 7344 -1960 7378 -1926
rect 7412 -1960 7446 -1926
rect 7480 -1960 7514 -1926
rect 7548 -1960 7582 -1926
rect 7616 -1960 7650 -1926
rect 7684 -1960 7718 -1926
rect 7752 -1960 7786 -1926
rect 7820 -1960 7854 -1926
rect 7888 -1960 7922 -1926
rect 7956 -1960 7990 -1926
rect 8024 -1960 8058 -1926
rect 8092 -1960 8126 -1926
rect 8160 -1960 8194 -1926
rect 8228 -1960 8262 -1926
rect 8296 -1960 8330 -1926
rect 8364 -1960 8398 -1926
rect 8432 -1960 8466 -1926
rect 8500 -1960 8534 -1926
rect 8568 -1960 8602 -1926
rect 8636 -1960 8670 -1926
rect 8704 -1960 8738 -1926
rect 8772 -1960 8806 -1926
rect 8840 -1960 8874 -1926
rect 8908 -1960 8942 -1926
rect 8976 -1960 9010 -1926
rect 9044 -1960 9078 -1926
rect 9112 -1960 9146 -1926
rect 9180 -1960 9214 -1926
rect 9248 -1960 9282 -1926
rect 9316 -1960 9350 -1926
rect 9384 -1960 9418 -1926
rect 9452 -1960 9486 -1926
rect 9694 -1960 9728 -1926
rect 9762 -1960 9796 -1926
rect 9830 -1960 9864 -1926
rect 9898 -1960 9932 -1926
rect 9966 -1960 10000 -1926
rect 10034 -1960 10068 -1926
rect 10102 -1960 10136 -1926
rect 10170 -1960 10204 -1926
rect 10238 -1960 10272 -1926
rect 10306 -1960 10340 -1926
rect 10374 -1960 10408 -1926
rect 10442 -1960 10476 -1926
rect 10510 -1960 10544 -1926
rect 10578 -1960 10612 -1926
rect 10646 -1960 10680 -1926
rect 10714 -1960 10748 -1926
rect 10782 -1960 10816 -1926
rect 10850 -1960 10884 -1926
rect 10918 -1960 10952 -1926
rect 10986 -1960 11020 -1926
rect 11054 -1960 11088 -1926
rect 11122 -1960 11156 -1926
rect 11190 -1960 11224 -1926
rect 11258 -1960 11292 -1926
rect 11326 -1960 11360 -1926
rect 11394 -1960 11428 -1926
rect 11462 -1960 11496 -1926
rect 11530 -1960 11564 -1926
rect 11598 -1960 11632 -1926
rect 11666 -1960 11700 -1926
rect 11734 -1960 11768 -1926
rect 11802 -1960 11836 -1926
rect 11870 -1960 11904 -1926
rect 11938 -1960 11972 -1926
rect 12006 -1960 12040 -1926
rect 12074 -1960 12108 -1926
rect 12142 -1960 12176 -1926
rect 12210 -1960 12244 -1926
rect 12278 -1960 12312 -1926
rect 12346 -1960 12380 -1926
rect 12414 -1960 12448 -1926
rect 12482 -1960 12516 -1926
rect 12550 -1960 12584 -1926
rect 12618 -1960 12652 -1926
rect 12686 -1960 12720 -1926
rect 12754 -1960 12788 -1926
rect 12822 -1960 12856 -1926
rect 12890 -1960 12924 -1926
rect 12958 -1960 12992 -1926
rect 13026 -1960 13060 -1926
rect 13094 -1960 13128 -1926
rect 13162 -1960 13196 -1926
rect 13230 -1960 13264 -1926
rect 13298 -1960 13332 -1926
rect 13366 -1960 13400 -1926
rect 13434 -1960 13468 -1926
rect 13502 -1960 13536 -1926
rect 13570 -1960 13604 -1926
rect 13638 -1960 13672 -1926
rect 13706 -1960 13740 -1926
rect 13774 -1960 13808 -1926
rect 14089 -1960 14123 -1926
rect 14157 -1960 14191 -1926
rect 14225 -1960 14259 -1926
rect 14293 -1960 14327 -1926
rect 14361 -1960 14395 -1926
rect 14429 -1960 14463 -1926
rect 14497 -1960 14531 -1926
rect 14565 -1960 14599 -1926
rect 14633 -1960 14667 -1926
rect 14701 -1960 14735 -1926
rect 14769 -1960 14803 -1926
rect 14837 -1960 14871 -1926
rect 14905 -1960 14939 -1926
rect 14973 -1960 15007 -1926
rect 15041 -1960 15075 -1926
rect 15109 -1960 15143 -1926
rect 15177 -1960 15211 -1926
rect 15245 -1960 15279 -1926
rect 15313 -1960 15347 -1926
rect 15381 -1960 15415 -1926
rect 15449 -1960 15483 -1926
rect 15517 -1960 15551 -1926
rect 15585 -1960 15619 -1926
rect 15653 -1960 15687 -1926
rect 15721 -1960 15755 -1926
rect 15789 -1960 15823 -1926
rect 15857 -1960 15891 -1926
rect 15925 -1960 15959 -1926
rect 15993 -1960 16027 -1926
rect 16061 -1960 16095 -1926
rect 16129 -1960 16163 -1926
rect 16197 -1960 16231 -1926
rect 16265 -1960 16299 -1926
rect 16333 -1960 16367 -1926
rect 16401 -1960 16435 -1926
rect 16469 -1960 16503 -1926
rect 16537 -1960 16571 -1926
rect 16605 -1960 16639 -1926
rect 16673 -1960 16707 -1926
rect 16741 -1960 16775 -1926
rect 16809 -1960 16843 -1926
rect 16877 -1960 16911 -1926
rect 16945 -1960 16979 -1926
rect 17013 -1960 17047 -1926
rect 17081 -1960 17115 -1926
rect 17149 -1960 17183 -1926
rect 17217 -1960 17251 -1926
rect 17285 -1960 17319 -1926
rect 17353 -1960 17387 -1926
rect 17421 -1960 17455 -1926
rect 17489 -1960 17523 -1926
rect 17557 -1960 17591 -1926
rect 17625 -1960 17659 -1926
rect 17693 -1960 17727 -1926
rect 17761 -1960 17795 -1926
rect 17829 -1960 17863 -1926
rect 17897 -1960 17931 -1926
rect 17965 -1960 17999 -1926
rect 18033 -1960 18067 -1926
rect 18101 -1960 18135 -1926
rect 18169 -1960 18203 -1926
rect 856 -2096 890 -2062
rect 856 -2164 890 -2130
rect 856 -2232 890 -2198
rect 856 -2300 890 -2266
rect 5214 -2096 5248 -2062
rect 5214 -2164 5248 -2130
rect 5214 -2232 5248 -2198
rect 5214 -2300 5248 -2266
rect 9573 -2096 9607 -2062
rect 9573 -2164 9607 -2130
rect 9573 -2232 9607 -2198
rect 856 -2368 890 -2334
rect 856 -2436 890 -2402
rect 856 -2504 890 -2470
rect 9573 -2300 9607 -2266
rect 13932 -2096 13966 -2062
rect 13932 -2164 13966 -2130
rect 13932 -2232 13966 -2198
rect 5214 -2368 5248 -2334
rect 5214 -2436 5248 -2402
rect 5214 -2504 5248 -2470
rect 856 -2572 890 -2538
rect 856 -2640 890 -2606
rect 13932 -2300 13966 -2266
rect 18290 -2096 18324 -2062
rect 18290 -2164 18324 -2130
rect 18290 -2232 18324 -2198
rect 9573 -2368 9607 -2334
rect 9573 -2436 9607 -2402
rect 9573 -2504 9607 -2470
rect 5214 -2572 5248 -2538
rect 856 -2708 890 -2674
rect 856 -2776 890 -2742
rect 856 -2844 890 -2810
rect 856 -2912 890 -2878
rect 5214 -2640 5248 -2606
rect 18290 -2300 18324 -2266
rect 13932 -2368 13966 -2334
rect 13932 -2436 13966 -2402
rect 13932 -2504 13966 -2470
rect 9573 -2572 9607 -2538
rect 5214 -2708 5248 -2674
rect 5214 -2776 5248 -2742
rect 5214 -2844 5248 -2810
rect 5214 -2912 5248 -2878
rect 856 -2980 890 -2946
rect 9573 -2640 9607 -2606
rect 18290 -2368 18324 -2334
rect 18290 -2436 18324 -2402
rect 18290 -2504 18324 -2470
rect 13932 -2572 13966 -2538
rect 9573 -2708 9607 -2674
rect 9573 -2776 9607 -2742
rect 9573 -2844 9607 -2810
rect 9573 -2912 9607 -2878
rect 5214 -2980 5248 -2946
rect 13932 -2640 13966 -2606
rect 18290 -2572 18324 -2538
rect 13932 -2708 13966 -2674
rect 13932 -2776 13966 -2742
rect 13932 -2844 13966 -2810
rect 13932 -2912 13966 -2878
rect 9573 -2980 9607 -2946
rect 18290 -2640 18324 -2606
rect 18290 -2708 18324 -2674
rect 18290 -2776 18324 -2742
rect 18290 -2844 18324 -2810
rect 18290 -2912 18324 -2878
rect 13932 -2980 13966 -2946
rect 18290 -2980 18324 -2946
rect 856 -3048 890 -3014
rect 856 -3116 890 -3082
rect 856 -3184 890 -3150
rect 5214 -3048 5248 -3014
rect 5214 -3116 5248 -3082
rect 5214 -3184 5248 -3150
rect 856 -3252 890 -3218
rect 9573 -3048 9607 -3014
rect 9573 -3116 9607 -3082
rect 9573 -3184 9607 -3150
rect 856 -3320 890 -3286
rect 856 -3388 890 -3354
rect 856 -3456 890 -3422
rect 856 -3524 890 -3490
rect 856 -3592 890 -3558
rect 5214 -3252 5248 -3218
rect 13932 -3048 13966 -3014
rect 13932 -3116 13966 -3082
rect 13932 -3184 13966 -3150
rect 5214 -3320 5248 -3286
rect 5214 -3388 5248 -3354
rect 5214 -3456 5248 -3422
rect 5214 -3524 5248 -3490
rect 5214 -3592 5248 -3558
rect 9573 -3252 9607 -3218
rect 18290 -3048 18324 -3014
rect 18290 -3116 18324 -3082
rect 18290 -3184 18324 -3150
rect 9573 -3320 9607 -3286
rect 9573 -3388 9607 -3354
rect 9573 -3456 9607 -3422
rect 9573 -3524 9607 -3490
rect 9573 -3592 9607 -3558
rect 13932 -3252 13966 -3218
rect 13932 -3320 13966 -3286
rect 13932 -3388 13966 -3354
rect 13932 -3456 13966 -3422
rect 13932 -3524 13966 -3490
rect 13932 -3592 13966 -3558
rect 18290 -3252 18324 -3218
rect 18290 -3320 18324 -3286
rect 18290 -3388 18324 -3354
rect 18290 -3456 18324 -3422
rect 18290 -3524 18324 -3490
rect 18290 -3592 18324 -3558
rect 977 -3626 1011 -3592
rect 1045 -3626 1079 -3592
rect 1113 -3626 1147 -3592
rect 1181 -3626 1215 -3592
rect 1249 -3626 1283 -3592
rect 1317 -3626 1351 -3592
rect 1385 -3626 1419 -3592
rect 1453 -3626 1487 -3592
rect 1521 -3626 1555 -3592
rect 1589 -3626 1623 -3592
rect 1657 -3626 1691 -3592
rect 1725 -3626 1759 -3592
rect 1793 -3626 1827 -3592
rect 1861 -3626 1895 -3592
rect 1929 -3626 1963 -3592
rect 1997 -3626 2031 -3592
rect 2065 -3626 2099 -3592
rect 2133 -3626 2167 -3592
rect 2201 -3626 2235 -3592
rect 2269 -3626 2303 -3592
rect 2337 -3626 2371 -3592
rect 2405 -3626 2439 -3592
rect 2473 -3626 2507 -3592
rect 2541 -3626 2575 -3592
rect 2609 -3626 2643 -3592
rect 2677 -3626 2711 -3592
rect 2745 -3626 2779 -3592
rect 2813 -3626 2847 -3592
rect 2881 -3626 2915 -3592
rect 2949 -3626 2983 -3592
rect 3017 -3626 3051 -3592
rect 3085 -3626 3119 -3592
rect 3153 -3626 3187 -3592
rect 3221 -3626 3255 -3592
rect 3289 -3626 3323 -3592
rect 3357 -3626 3391 -3592
rect 3425 -3626 3459 -3592
rect 3493 -3626 3527 -3592
rect 3561 -3626 3595 -3592
rect 3629 -3626 3663 -3592
rect 3697 -3626 3731 -3592
rect 3765 -3626 3799 -3592
rect 3833 -3626 3867 -3592
rect 3901 -3626 3935 -3592
rect 3969 -3626 4003 -3592
rect 4037 -3626 4071 -3592
rect 4105 -3626 4139 -3592
rect 4173 -3626 4207 -3592
rect 4241 -3626 4275 -3592
rect 4309 -3626 4343 -3592
rect 4377 -3626 4411 -3592
rect 4445 -3626 4479 -3592
rect 4513 -3626 4547 -3592
rect 4581 -3626 4615 -3592
rect 4649 -3626 4683 -3592
rect 4717 -3626 4751 -3592
rect 4785 -3626 4819 -3592
rect 4853 -3626 4887 -3592
rect 4921 -3626 4955 -3592
rect 4989 -3626 5023 -3592
rect 5057 -3626 5091 -3592
rect 5372 -3626 5406 -3592
rect 5440 -3626 5474 -3592
rect 5508 -3626 5542 -3592
rect 5576 -3626 5610 -3592
rect 5644 -3626 5678 -3592
rect 5712 -3626 5746 -3592
rect 5780 -3626 5814 -3592
rect 5848 -3626 5882 -3592
rect 5916 -3626 5950 -3592
rect 5984 -3626 6018 -3592
rect 6052 -3626 6086 -3592
rect 6120 -3626 6154 -3592
rect 6188 -3626 6222 -3592
rect 6256 -3626 6290 -3592
rect 6324 -3626 6358 -3592
rect 6392 -3626 6426 -3592
rect 6460 -3626 6494 -3592
rect 6528 -3626 6562 -3592
rect 6596 -3626 6630 -3592
rect 6664 -3626 6698 -3592
rect 6732 -3626 6766 -3592
rect 6800 -3626 6834 -3592
rect 6868 -3626 6902 -3592
rect 6936 -3626 6970 -3592
rect 7004 -3626 7038 -3592
rect 7072 -3626 7106 -3592
rect 7140 -3626 7174 -3592
rect 7208 -3626 7242 -3592
rect 7276 -3626 7310 -3592
rect 7344 -3626 7378 -3592
rect 7412 -3626 7446 -3592
rect 7480 -3626 7514 -3592
rect 7548 -3626 7582 -3592
rect 7616 -3626 7650 -3592
rect 7684 -3626 7718 -3592
rect 7752 -3626 7786 -3592
rect 7820 -3626 7854 -3592
rect 7888 -3626 7922 -3592
rect 7956 -3626 7990 -3592
rect 8024 -3626 8058 -3592
rect 8092 -3626 8126 -3592
rect 8160 -3626 8194 -3592
rect 8228 -3626 8262 -3592
rect 8296 -3626 8330 -3592
rect 8364 -3626 8398 -3592
rect 8432 -3626 8466 -3592
rect 8500 -3626 8534 -3592
rect 8568 -3626 8602 -3592
rect 8636 -3626 8670 -3592
rect 8704 -3626 8738 -3592
rect 8772 -3626 8806 -3592
rect 8840 -3626 8874 -3592
rect 8908 -3626 8942 -3592
rect 8976 -3626 9010 -3592
rect 9044 -3626 9078 -3592
rect 9112 -3626 9146 -3592
rect 9180 -3626 9214 -3592
rect 9248 -3626 9282 -3592
rect 9316 -3626 9350 -3592
rect 9384 -3626 9418 -3592
rect 9452 -3626 9486 -3592
rect 9694 -3626 9728 -3592
rect 9762 -3626 9796 -3592
rect 9830 -3626 9864 -3592
rect 9898 -3626 9932 -3592
rect 9966 -3626 10000 -3592
rect 10034 -3626 10068 -3592
rect 10102 -3626 10136 -3592
rect 10170 -3626 10204 -3592
rect 10238 -3626 10272 -3592
rect 10306 -3626 10340 -3592
rect 10374 -3626 10408 -3592
rect 10442 -3626 10476 -3592
rect 10510 -3626 10544 -3592
rect 10578 -3626 10612 -3592
rect 10646 -3626 10680 -3592
rect 10714 -3626 10748 -3592
rect 10782 -3626 10816 -3592
rect 10850 -3626 10884 -3592
rect 10918 -3626 10952 -3592
rect 10986 -3626 11020 -3592
rect 11054 -3626 11088 -3592
rect 11122 -3626 11156 -3592
rect 11190 -3626 11224 -3592
rect 11258 -3626 11292 -3592
rect 11326 -3626 11360 -3592
rect 11394 -3626 11428 -3592
rect 11462 -3626 11496 -3592
rect 11530 -3626 11564 -3592
rect 11598 -3626 11632 -3592
rect 11666 -3626 11700 -3592
rect 11734 -3626 11768 -3592
rect 11802 -3626 11836 -3592
rect 11870 -3626 11904 -3592
rect 11938 -3626 11972 -3592
rect 12006 -3626 12040 -3592
rect 12074 -3626 12108 -3592
rect 12142 -3626 12176 -3592
rect 12210 -3626 12244 -3592
rect 12278 -3626 12312 -3592
rect 12346 -3626 12380 -3592
rect 12414 -3626 12448 -3592
rect 12482 -3626 12516 -3592
rect 12550 -3626 12584 -3592
rect 12618 -3626 12652 -3592
rect 12686 -3626 12720 -3592
rect 12754 -3626 12788 -3592
rect 12822 -3626 12856 -3592
rect 12890 -3626 12924 -3592
rect 12958 -3626 12992 -3592
rect 13026 -3626 13060 -3592
rect 13094 -3626 13128 -3592
rect 13162 -3626 13196 -3592
rect 13230 -3626 13264 -3592
rect 13298 -3626 13332 -3592
rect 13366 -3626 13400 -3592
rect 13434 -3626 13468 -3592
rect 13502 -3626 13536 -3592
rect 13570 -3626 13604 -3592
rect 13638 -3626 13672 -3592
rect 13706 -3626 13740 -3592
rect 13774 -3626 13808 -3592
rect 14089 -3626 14123 -3592
rect 14157 -3626 14191 -3592
rect 14225 -3626 14259 -3592
rect 14293 -3626 14327 -3592
rect 14361 -3626 14395 -3592
rect 14429 -3626 14463 -3592
rect 14497 -3626 14531 -3592
rect 14565 -3626 14599 -3592
rect 14633 -3626 14667 -3592
rect 14701 -3626 14735 -3592
rect 14769 -3626 14803 -3592
rect 14837 -3626 14871 -3592
rect 14905 -3626 14939 -3592
rect 14973 -3626 15007 -3592
rect 15041 -3626 15075 -3592
rect 15109 -3626 15143 -3592
rect 15177 -3626 15211 -3592
rect 15245 -3626 15279 -3592
rect 15313 -3626 15347 -3592
rect 15381 -3626 15415 -3592
rect 15449 -3626 15483 -3592
rect 15517 -3626 15551 -3592
rect 15585 -3626 15619 -3592
rect 15653 -3626 15687 -3592
rect 15721 -3626 15755 -3592
rect 15789 -3626 15823 -3592
rect 15857 -3626 15891 -3592
rect 15925 -3626 15959 -3592
rect 15993 -3626 16027 -3592
rect 16061 -3626 16095 -3592
rect 16129 -3626 16163 -3592
rect 16197 -3626 16231 -3592
rect 16265 -3626 16299 -3592
rect 16333 -3626 16367 -3592
rect 16401 -3626 16435 -3592
rect 16469 -3626 16503 -3592
rect 16537 -3626 16571 -3592
rect 16605 -3626 16639 -3592
rect 16673 -3626 16707 -3592
rect 16741 -3626 16775 -3592
rect 16809 -3626 16843 -3592
rect 16877 -3626 16911 -3592
rect 16945 -3626 16979 -3592
rect 17013 -3626 17047 -3592
rect 17081 -3626 17115 -3592
rect 17149 -3626 17183 -3592
rect 17217 -3626 17251 -3592
rect 17285 -3626 17319 -3592
rect 17353 -3626 17387 -3592
rect 17421 -3626 17455 -3592
rect 17489 -3626 17523 -3592
rect 17557 -3626 17591 -3592
rect 17625 -3626 17659 -3592
rect 17693 -3626 17727 -3592
rect 17761 -3626 17795 -3592
rect 17829 -3626 17863 -3592
rect 17897 -3626 17931 -3592
rect 17965 -3626 17999 -3592
rect 18033 -3626 18067 -3592
rect 18101 -3626 18135 -3592
rect 18169 -3626 18203 -3592
rect 856 -3660 890 -3626
rect 856 -3728 890 -3694
rect 856 -3796 890 -3762
rect 856 -3864 890 -3830
rect 856 -3932 890 -3898
rect 856 -4000 890 -3966
rect 5214 -3660 5248 -3626
rect 5214 -3728 5248 -3694
rect 5214 -3796 5248 -3762
rect 5214 -3864 5248 -3830
rect 5214 -3932 5248 -3898
rect 5214 -4000 5248 -3966
rect 9573 -3660 9607 -3626
rect 9573 -3728 9607 -3694
rect 9573 -3796 9607 -3762
rect 9573 -3864 9607 -3830
rect 9573 -3932 9607 -3898
rect 856 -4068 890 -4034
rect 856 -4136 890 -4102
rect 9573 -4000 9607 -3966
rect 13932 -3660 13966 -3626
rect 13932 -3728 13966 -3694
rect 13932 -3796 13966 -3762
rect 13932 -3864 13966 -3830
rect 13932 -3932 13966 -3898
rect 5214 -4068 5248 -4034
rect 5214 -4136 5248 -4102
rect 13932 -4000 13966 -3966
rect 18290 -3660 18324 -3626
rect 18290 -3728 18324 -3694
rect 18290 -3796 18324 -3762
rect 18290 -3864 18324 -3830
rect 18290 -3932 18324 -3898
rect 9573 -4068 9607 -4034
rect 9573 -4136 9607 -4102
rect 18290 -4000 18324 -3966
rect 13932 -4068 13966 -4034
rect 13932 -4136 13966 -4102
rect 18290 -4068 18324 -4034
rect 18290 -4136 18324 -4102
rect 977 -4399 1011 -4365
rect 1045 -4399 1079 -4365
rect 1113 -4399 1147 -4365
rect 1181 -4399 1215 -4365
rect 1249 -4399 1283 -4365
rect 1317 -4399 1351 -4365
rect 1385 -4399 1419 -4365
rect 1453 -4399 1487 -4365
rect 1521 -4399 1555 -4365
rect 1589 -4399 1623 -4365
rect 1657 -4399 1691 -4365
rect 1725 -4399 1759 -4365
rect 1793 -4399 1827 -4365
rect 1861 -4399 1895 -4365
rect 1929 -4399 1963 -4365
rect 1997 -4399 2031 -4365
rect 2065 -4399 2099 -4365
rect 2133 -4399 2167 -4365
rect 2201 -4399 2235 -4365
rect 2269 -4399 2303 -4365
rect 2337 -4399 2371 -4365
rect 2405 -4399 2439 -4365
rect 2473 -4399 2507 -4365
rect 2541 -4399 2575 -4365
rect 2609 -4399 2643 -4365
rect 2677 -4399 2711 -4365
rect 2745 -4399 2779 -4365
rect 2813 -4399 2847 -4365
rect 2881 -4399 2915 -4365
rect 2949 -4399 2983 -4365
rect 3017 -4399 3051 -4365
rect 3085 -4399 3119 -4365
rect 3153 -4399 3187 -4365
rect 3221 -4399 3255 -4365
rect 3289 -4399 3323 -4365
rect 3357 -4399 3391 -4365
rect 3425 -4399 3459 -4365
rect 3493 -4399 3527 -4365
rect 3561 -4399 3595 -4365
rect 3629 -4399 3663 -4365
rect 3697 -4399 3731 -4365
rect 3765 -4399 3799 -4365
rect 3833 -4399 3867 -4365
rect 3901 -4399 3935 -4365
rect 3969 -4399 4003 -4365
rect 4037 -4399 4071 -4365
rect 4105 -4399 4139 -4365
rect 4173 -4399 4207 -4365
rect 4241 -4399 4275 -4365
rect 4309 -4399 4343 -4365
rect 4377 -4399 4411 -4365
rect 4445 -4399 4479 -4365
rect 4513 -4399 4547 -4365
rect 4581 -4399 4615 -4365
rect 4649 -4399 4683 -4365
rect 4717 -4399 4751 -4365
rect 4785 -4399 4819 -4365
rect 4853 -4399 4887 -4365
rect 4921 -4399 4955 -4365
rect 4989 -4399 5023 -4365
rect 5057 -4399 5091 -4365
rect 5372 -4399 5406 -4365
rect 5440 -4399 5474 -4365
rect 5508 -4399 5542 -4365
rect 5576 -4399 5610 -4365
rect 5644 -4399 5678 -4365
rect 5712 -4399 5746 -4365
rect 5780 -4399 5814 -4365
rect 5848 -4399 5882 -4365
rect 5916 -4399 5950 -4365
rect 5984 -4399 6018 -4365
rect 6052 -4399 6086 -4365
rect 6120 -4399 6154 -4365
rect 6188 -4399 6222 -4365
rect 6256 -4399 6290 -4365
rect 6324 -4399 6358 -4365
rect 6392 -4399 6426 -4365
rect 6460 -4399 6494 -4365
rect 6528 -4399 6562 -4365
rect 6596 -4399 6630 -4365
rect 6664 -4399 6698 -4365
rect 6732 -4399 6766 -4365
rect 6800 -4399 6834 -4365
rect 6868 -4399 6902 -4365
rect 6936 -4399 6970 -4365
rect 7004 -4399 7038 -4365
rect 7072 -4399 7106 -4365
rect 7140 -4399 7174 -4365
rect 7208 -4399 7242 -4365
rect 7276 -4399 7310 -4365
rect 7344 -4399 7378 -4365
rect 7412 -4399 7446 -4365
rect 7480 -4399 7514 -4365
rect 7548 -4399 7582 -4365
rect 7616 -4399 7650 -4365
rect 7684 -4399 7718 -4365
rect 7752 -4399 7786 -4365
rect 7820 -4399 7854 -4365
rect 7888 -4399 7922 -4365
rect 7956 -4399 7990 -4365
rect 8024 -4399 8058 -4365
rect 8092 -4399 8126 -4365
rect 8160 -4399 8194 -4365
rect 8228 -4399 8262 -4365
rect 8296 -4399 8330 -4365
rect 8364 -4399 8398 -4365
rect 8432 -4399 8466 -4365
rect 8500 -4399 8534 -4365
rect 8568 -4399 8602 -4365
rect 8636 -4399 8670 -4365
rect 8704 -4399 8738 -4365
rect 8772 -4399 8806 -4365
rect 8840 -4399 8874 -4365
rect 8908 -4399 8942 -4365
rect 8976 -4399 9010 -4365
rect 9044 -4399 9078 -4365
rect 9112 -4399 9146 -4365
rect 9180 -4399 9214 -4365
rect 9248 -4399 9282 -4365
rect 9316 -4399 9350 -4365
rect 9384 -4399 9418 -4365
rect 9452 -4399 9486 -4365
rect 9694 -4399 9728 -4365
rect 9762 -4399 9796 -4365
rect 9830 -4399 9864 -4365
rect 9898 -4399 9932 -4365
rect 9966 -4399 10000 -4365
rect 10034 -4399 10068 -4365
rect 10102 -4399 10136 -4365
rect 10170 -4399 10204 -4365
rect 10238 -4399 10272 -4365
rect 10306 -4399 10340 -4365
rect 10374 -4399 10408 -4365
rect 10442 -4399 10476 -4365
rect 10510 -4399 10544 -4365
rect 10578 -4399 10612 -4365
rect 10646 -4399 10680 -4365
rect 10714 -4399 10748 -4365
rect 10782 -4399 10816 -4365
rect 10850 -4399 10884 -4365
rect 10918 -4399 10952 -4365
rect 10986 -4399 11020 -4365
rect 11054 -4399 11088 -4365
rect 11122 -4399 11156 -4365
rect 11190 -4399 11224 -4365
rect 11258 -4399 11292 -4365
rect 11326 -4399 11360 -4365
rect 11394 -4399 11428 -4365
rect 11462 -4399 11496 -4365
rect 11530 -4399 11564 -4365
rect 11598 -4399 11632 -4365
rect 11666 -4399 11700 -4365
rect 11734 -4399 11768 -4365
rect 11802 -4399 11836 -4365
rect 11870 -4399 11904 -4365
rect 11938 -4399 11972 -4365
rect 12006 -4399 12040 -4365
rect 12074 -4399 12108 -4365
rect 12142 -4399 12176 -4365
rect 12210 -4399 12244 -4365
rect 12278 -4399 12312 -4365
rect 12346 -4399 12380 -4365
rect 12414 -4399 12448 -4365
rect 12482 -4399 12516 -4365
rect 12550 -4399 12584 -4365
rect 12618 -4399 12652 -4365
rect 12686 -4399 12720 -4365
rect 12754 -4399 12788 -4365
rect 12822 -4399 12856 -4365
rect 12890 -4399 12924 -4365
rect 12958 -4399 12992 -4365
rect 13026 -4399 13060 -4365
rect 13094 -4399 13128 -4365
rect 13162 -4399 13196 -4365
rect 13230 -4399 13264 -4365
rect 13298 -4399 13332 -4365
rect 13366 -4399 13400 -4365
rect 13434 -4399 13468 -4365
rect 13502 -4399 13536 -4365
rect 13570 -4399 13604 -4365
rect 13638 -4399 13672 -4365
rect 13706 -4399 13740 -4365
rect 13774 -4399 13808 -4365
rect 14089 -4399 14123 -4365
rect 14157 -4399 14191 -4365
rect 14225 -4399 14259 -4365
rect 14293 -4399 14327 -4365
rect 14361 -4399 14395 -4365
rect 14429 -4399 14463 -4365
rect 14497 -4399 14531 -4365
rect 14565 -4399 14599 -4365
rect 14633 -4399 14667 -4365
rect 14701 -4399 14735 -4365
rect 14769 -4399 14803 -4365
rect 14837 -4399 14871 -4365
rect 14905 -4399 14939 -4365
rect 14973 -4399 15007 -4365
rect 15041 -4399 15075 -4365
rect 15109 -4399 15143 -4365
rect 15177 -4399 15211 -4365
rect 15245 -4399 15279 -4365
rect 15313 -4399 15347 -4365
rect 15381 -4399 15415 -4365
rect 15449 -4399 15483 -4365
rect 15517 -4399 15551 -4365
rect 15585 -4399 15619 -4365
rect 15653 -4399 15687 -4365
rect 15721 -4399 15755 -4365
rect 15789 -4399 15823 -4365
rect 15857 -4399 15891 -4365
rect 15925 -4399 15959 -4365
rect 15993 -4399 16027 -4365
rect 16061 -4399 16095 -4365
rect 16129 -4399 16163 -4365
rect 16197 -4399 16231 -4365
rect 16265 -4399 16299 -4365
rect 16333 -4399 16367 -4365
rect 16401 -4399 16435 -4365
rect 16469 -4399 16503 -4365
rect 16537 -4399 16571 -4365
rect 16605 -4399 16639 -4365
rect 16673 -4399 16707 -4365
rect 16741 -4399 16775 -4365
rect 16809 -4399 16843 -4365
rect 16877 -4399 16911 -4365
rect 16945 -4399 16979 -4365
rect 17013 -4399 17047 -4365
rect 17081 -4399 17115 -4365
rect 17149 -4399 17183 -4365
rect 17217 -4399 17251 -4365
rect 17285 -4399 17319 -4365
rect 17353 -4399 17387 -4365
rect 17421 -4399 17455 -4365
rect 17489 -4399 17523 -4365
rect 17557 -4399 17591 -4365
rect 17625 -4399 17659 -4365
rect 17693 -4399 17727 -4365
rect 17761 -4399 17795 -4365
rect 17829 -4399 17863 -4365
rect 17897 -4399 17931 -4365
rect 17965 -4399 17999 -4365
rect 18033 -4399 18067 -4365
rect 18101 -4399 18135 -4365
rect 18169 -4399 18203 -4365
rect 856 -4662 890 -4628
rect 856 -4730 890 -4696
rect 5214 -4662 5248 -4628
rect 5214 -4730 5248 -4696
rect 856 -4798 890 -4764
rect 9573 -4662 9607 -4628
rect 9573 -4730 9607 -4696
rect 856 -4866 890 -4832
rect 856 -4934 890 -4900
rect 856 -5002 890 -4968
rect 856 -5070 890 -5036
rect 856 -5138 890 -5104
rect 5214 -4798 5248 -4764
rect 13932 -4662 13966 -4628
rect 13932 -4730 13966 -4696
rect 5214 -4866 5248 -4832
rect 5214 -4934 5248 -4900
rect 5214 -5002 5248 -4968
rect 5214 -5070 5248 -5036
rect 5214 -5138 5248 -5104
rect 9573 -4798 9607 -4764
rect 18290 -4662 18324 -4628
rect 18290 -4730 18324 -4696
rect 9573 -4866 9607 -4832
rect 9573 -4934 9607 -4900
rect 9573 -5002 9607 -4968
rect 9573 -5070 9607 -5036
rect 9573 -5138 9607 -5104
rect 13932 -4798 13966 -4764
rect 13932 -4866 13966 -4832
rect 13932 -4934 13966 -4900
rect 13932 -5002 13966 -4968
rect 13932 -5070 13966 -5036
rect 13932 -5138 13966 -5104
rect 18290 -4798 18324 -4764
rect 18290 -4866 18324 -4832
rect 18290 -4934 18324 -4900
rect 18290 -5002 18324 -4968
rect 18290 -5070 18324 -5036
rect 18290 -5138 18324 -5104
rect 977 -5172 1011 -5138
rect 1045 -5172 1079 -5138
rect 1113 -5172 1147 -5138
rect 1181 -5172 1215 -5138
rect 1249 -5172 1283 -5138
rect 1317 -5172 1351 -5138
rect 1385 -5172 1419 -5138
rect 1453 -5172 1487 -5138
rect 1521 -5172 1555 -5138
rect 1589 -5172 1623 -5138
rect 1657 -5172 1691 -5138
rect 1725 -5172 1759 -5138
rect 1793 -5172 1827 -5138
rect 1861 -5172 1895 -5138
rect 1929 -5172 1963 -5138
rect 1997 -5172 2031 -5138
rect 2065 -5172 2099 -5138
rect 2133 -5172 2167 -5138
rect 2201 -5172 2235 -5138
rect 2269 -5172 2303 -5138
rect 2337 -5172 2371 -5138
rect 2405 -5172 2439 -5138
rect 2473 -5172 2507 -5138
rect 2541 -5172 2575 -5138
rect 2609 -5172 2643 -5138
rect 2677 -5172 2711 -5138
rect 2745 -5172 2779 -5138
rect 2813 -5172 2847 -5138
rect 2881 -5172 2915 -5138
rect 2949 -5172 2983 -5138
rect 3017 -5172 3051 -5138
rect 3085 -5172 3119 -5138
rect 3153 -5172 3187 -5138
rect 3221 -5172 3255 -5138
rect 3289 -5172 3323 -5138
rect 3357 -5172 3391 -5138
rect 3425 -5172 3459 -5138
rect 3493 -5172 3527 -5138
rect 3561 -5172 3595 -5138
rect 3629 -5172 3663 -5138
rect 3697 -5172 3731 -5138
rect 3765 -5172 3799 -5138
rect 3833 -5172 3867 -5138
rect 3901 -5172 3935 -5138
rect 3969 -5172 4003 -5138
rect 4037 -5172 4071 -5138
rect 4105 -5172 4139 -5138
rect 4173 -5172 4207 -5138
rect 4241 -5172 4275 -5138
rect 4309 -5172 4343 -5138
rect 4377 -5172 4411 -5138
rect 4445 -5172 4479 -5138
rect 4513 -5172 4547 -5138
rect 4581 -5172 4615 -5138
rect 4649 -5172 4683 -5138
rect 4717 -5172 4751 -5138
rect 4785 -5172 4819 -5138
rect 4853 -5172 4887 -5138
rect 4921 -5172 4955 -5138
rect 4989 -5172 5023 -5138
rect 5057 -5172 5091 -5138
rect 5372 -5172 5406 -5138
rect 5440 -5172 5474 -5138
rect 5508 -5172 5542 -5138
rect 5576 -5172 5610 -5138
rect 5644 -5172 5678 -5138
rect 5712 -5172 5746 -5138
rect 5780 -5172 5814 -5138
rect 5848 -5172 5882 -5138
rect 5916 -5172 5950 -5138
rect 5984 -5172 6018 -5138
rect 6052 -5172 6086 -5138
rect 6120 -5172 6154 -5138
rect 6188 -5172 6222 -5138
rect 6256 -5172 6290 -5138
rect 6324 -5172 6358 -5138
rect 6392 -5172 6426 -5138
rect 6460 -5172 6494 -5138
rect 6528 -5172 6562 -5138
rect 6596 -5172 6630 -5138
rect 6664 -5172 6698 -5138
rect 6732 -5172 6766 -5138
rect 6800 -5172 6834 -5138
rect 6868 -5172 6902 -5138
rect 6936 -5172 6970 -5138
rect 7004 -5172 7038 -5138
rect 7072 -5172 7106 -5138
rect 7140 -5172 7174 -5138
rect 7208 -5172 7242 -5138
rect 7276 -5172 7310 -5138
rect 7344 -5172 7378 -5138
rect 7412 -5172 7446 -5138
rect 7480 -5172 7514 -5138
rect 7548 -5172 7582 -5138
rect 7616 -5172 7650 -5138
rect 7684 -5172 7718 -5138
rect 7752 -5172 7786 -5138
rect 7820 -5172 7854 -5138
rect 7888 -5172 7922 -5138
rect 7956 -5172 7990 -5138
rect 8024 -5172 8058 -5138
rect 8092 -5172 8126 -5138
rect 8160 -5172 8194 -5138
rect 8228 -5172 8262 -5138
rect 8296 -5172 8330 -5138
rect 8364 -5172 8398 -5138
rect 8432 -5172 8466 -5138
rect 8500 -5172 8534 -5138
rect 8568 -5172 8602 -5138
rect 8636 -5172 8670 -5138
rect 8704 -5172 8738 -5138
rect 8772 -5172 8806 -5138
rect 8840 -5172 8874 -5138
rect 8908 -5172 8942 -5138
rect 8976 -5172 9010 -5138
rect 9044 -5172 9078 -5138
rect 9112 -5172 9146 -5138
rect 9180 -5172 9214 -5138
rect 9248 -5172 9282 -5138
rect 9316 -5172 9350 -5138
rect 9384 -5172 9418 -5138
rect 9452 -5172 9486 -5138
rect 9694 -5172 9728 -5138
rect 9762 -5172 9796 -5138
rect 9830 -5172 9864 -5138
rect 9898 -5172 9932 -5138
rect 9966 -5172 10000 -5138
rect 10034 -5172 10068 -5138
rect 10102 -5172 10136 -5138
rect 10170 -5172 10204 -5138
rect 10238 -5172 10272 -5138
rect 10306 -5172 10340 -5138
rect 10374 -5172 10408 -5138
rect 10442 -5172 10476 -5138
rect 10510 -5172 10544 -5138
rect 10578 -5172 10612 -5138
rect 10646 -5172 10680 -5138
rect 10714 -5172 10748 -5138
rect 10782 -5172 10816 -5138
rect 10850 -5172 10884 -5138
rect 10918 -5172 10952 -5138
rect 10986 -5172 11020 -5138
rect 11054 -5172 11088 -5138
rect 11122 -5172 11156 -5138
rect 11190 -5172 11224 -5138
rect 11258 -5172 11292 -5138
rect 11326 -5172 11360 -5138
rect 11394 -5172 11428 -5138
rect 11462 -5172 11496 -5138
rect 11530 -5172 11564 -5138
rect 11598 -5172 11632 -5138
rect 11666 -5172 11700 -5138
rect 11734 -5172 11768 -5138
rect 11802 -5172 11836 -5138
rect 11870 -5172 11904 -5138
rect 11938 -5172 11972 -5138
rect 12006 -5172 12040 -5138
rect 12074 -5172 12108 -5138
rect 12142 -5172 12176 -5138
rect 12210 -5172 12244 -5138
rect 12278 -5172 12312 -5138
rect 12346 -5172 12380 -5138
rect 12414 -5172 12448 -5138
rect 12482 -5172 12516 -5138
rect 12550 -5172 12584 -5138
rect 12618 -5172 12652 -5138
rect 12686 -5172 12720 -5138
rect 12754 -5172 12788 -5138
rect 12822 -5172 12856 -5138
rect 12890 -5172 12924 -5138
rect 12958 -5172 12992 -5138
rect 13026 -5172 13060 -5138
rect 13094 -5172 13128 -5138
rect 13162 -5172 13196 -5138
rect 13230 -5172 13264 -5138
rect 13298 -5172 13332 -5138
rect 13366 -5172 13400 -5138
rect 13434 -5172 13468 -5138
rect 13502 -5172 13536 -5138
rect 13570 -5172 13604 -5138
rect 13638 -5172 13672 -5138
rect 13706 -5172 13740 -5138
rect 13774 -5172 13808 -5138
rect 14089 -5172 14123 -5138
rect 14157 -5172 14191 -5138
rect 14225 -5172 14259 -5138
rect 14293 -5172 14327 -5138
rect 14361 -5172 14395 -5138
rect 14429 -5172 14463 -5138
rect 14497 -5172 14531 -5138
rect 14565 -5172 14599 -5138
rect 14633 -5172 14667 -5138
rect 14701 -5172 14735 -5138
rect 14769 -5172 14803 -5138
rect 14837 -5172 14871 -5138
rect 14905 -5172 14939 -5138
rect 14973 -5172 15007 -5138
rect 15041 -5172 15075 -5138
rect 15109 -5172 15143 -5138
rect 15177 -5172 15211 -5138
rect 15245 -5172 15279 -5138
rect 15313 -5172 15347 -5138
rect 15381 -5172 15415 -5138
rect 15449 -5172 15483 -5138
rect 15517 -5172 15551 -5138
rect 15585 -5172 15619 -5138
rect 15653 -5172 15687 -5138
rect 15721 -5172 15755 -5138
rect 15789 -5172 15823 -5138
rect 15857 -5172 15891 -5138
rect 15925 -5172 15959 -5138
rect 15993 -5172 16027 -5138
rect 16061 -5172 16095 -5138
rect 16129 -5172 16163 -5138
rect 16197 -5172 16231 -5138
rect 16265 -5172 16299 -5138
rect 16333 -5172 16367 -5138
rect 16401 -5172 16435 -5138
rect 16469 -5172 16503 -5138
rect 16537 -5172 16571 -5138
rect 16605 -5172 16639 -5138
rect 16673 -5172 16707 -5138
rect 16741 -5172 16775 -5138
rect 16809 -5172 16843 -5138
rect 16877 -5172 16911 -5138
rect 16945 -5172 16979 -5138
rect 17013 -5172 17047 -5138
rect 17081 -5172 17115 -5138
rect 17149 -5172 17183 -5138
rect 17217 -5172 17251 -5138
rect 17285 -5172 17319 -5138
rect 17353 -5172 17387 -5138
rect 17421 -5172 17455 -5138
rect 17489 -5172 17523 -5138
rect 17557 -5172 17591 -5138
rect 17625 -5172 17659 -5138
rect 17693 -5172 17727 -5138
rect 17761 -5172 17795 -5138
rect 17829 -5172 17863 -5138
rect 17897 -5172 17931 -5138
rect 17965 -5172 17999 -5138
rect 18033 -5172 18067 -5138
rect 18101 -5172 18135 -5138
rect 18169 -5172 18203 -5138
rect 856 -5206 890 -5172
rect 856 -5274 890 -5240
rect 856 -5342 890 -5308
rect 856 -5410 890 -5376
rect 856 -5478 890 -5444
rect 856 -5546 890 -5512
rect 5214 -5206 5248 -5172
rect 5214 -5274 5248 -5240
rect 5214 -5342 5248 -5308
rect 5214 -5410 5248 -5376
rect 5214 -5478 5248 -5444
rect 5214 -5546 5248 -5512
rect 9573 -5206 9607 -5172
rect 9573 -5274 9607 -5240
rect 9573 -5342 9607 -5308
rect 9573 -5410 9607 -5376
rect 9573 -5478 9607 -5444
rect 856 -5614 890 -5580
rect 856 -5682 890 -5648
rect 856 -5750 890 -5716
rect 9573 -5546 9607 -5512
rect 13932 -5206 13966 -5172
rect 13932 -5274 13966 -5240
rect 13932 -5342 13966 -5308
rect 13932 -5410 13966 -5376
rect 13932 -5478 13966 -5444
rect 5214 -5614 5248 -5580
rect 5214 -5682 5248 -5648
rect 5214 -5750 5248 -5716
rect 13932 -5546 13966 -5512
rect 18290 -5206 18324 -5172
rect 18290 -5274 18324 -5240
rect 18290 -5342 18324 -5308
rect 18290 -5410 18324 -5376
rect 18290 -5478 18324 -5444
rect 9573 -5614 9607 -5580
rect 9573 -5682 9607 -5648
rect 9573 -5750 9607 -5716
rect 18290 -5546 18324 -5512
rect 13932 -5614 13966 -5580
rect 13932 -5682 13966 -5648
rect 13932 -5750 13966 -5716
rect 18290 -5614 18324 -5580
rect 18290 -5682 18324 -5648
rect 18290 -5750 18324 -5716
rect 856 -5818 890 -5784
rect 5214 -5818 5248 -5784
rect 856 -5886 890 -5852
rect 856 -5954 890 -5920
rect 856 -6022 890 -5988
rect 856 -6090 890 -6056
rect 856 -6158 890 -6124
rect 9573 -5818 9607 -5784
rect 5214 -5886 5248 -5852
rect 5214 -5954 5248 -5920
rect 5214 -6022 5248 -5988
rect 5214 -6090 5248 -6056
rect 856 -6226 890 -6192
rect 5214 -6158 5248 -6124
rect 13932 -5818 13966 -5784
rect 9573 -5886 9607 -5852
rect 9573 -5954 9607 -5920
rect 9573 -6022 9607 -5988
rect 9573 -6090 9607 -6056
rect 5214 -6226 5248 -6192
rect 856 -6294 890 -6260
rect 856 -6362 890 -6328
rect 856 -6430 890 -6396
rect 9573 -6158 9607 -6124
rect 18290 -5818 18324 -5784
rect 13932 -5886 13966 -5852
rect 13932 -5954 13966 -5920
rect 13932 -6022 13966 -5988
rect 13932 -6090 13966 -6056
rect 9573 -6226 9607 -6192
rect 5214 -6294 5248 -6260
rect 5214 -6362 5248 -6328
rect 5214 -6430 5248 -6396
rect 856 -6498 890 -6464
rect 13932 -6158 13966 -6124
rect 18290 -5886 18324 -5852
rect 18290 -5954 18324 -5920
rect 18290 -6022 18324 -5988
rect 18290 -6090 18324 -6056
rect 13932 -6226 13966 -6192
rect 9573 -6294 9607 -6260
rect 9573 -6362 9607 -6328
rect 9573 -6430 9607 -6396
rect 856 -6566 890 -6532
rect 856 -6634 890 -6600
rect 856 -6702 890 -6668
rect 5214 -6498 5248 -6464
rect 18290 -6158 18324 -6124
rect 18290 -6226 18324 -6192
rect 13932 -6294 13966 -6260
rect 13932 -6362 13966 -6328
rect 13932 -6430 13966 -6396
rect 5214 -6566 5248 -6532
rect 5214 -6634 5248 -6600
rect 5214 -6702 5248 -6668
rect 9573 -6498 9607 -6464
rect 18290 -6294 18324 -6260
rect 18290 -6362 18324 -6328
rect 18290 -6430 18324 -6396
rect 9573 -6566 9607 -6532
rect 9573 -6634 9607 -6600
rect 9573 -6702 9607 -6668
rect 13932 -6498 13966 -6464
rect 13932 -6566 13966 -6532
rect 13932 -6634 13966 -6600
rect 13932 -6702 13966 -6668
rect 18290 -6498 18324 -6464
rect 18290 -6566 18324 -6532
rect 18290 -6634 18324 -6600
rect 18290 -6702 18324 -6668
rect 977 -6838 1011 -6804
rect 1045 -6838 1079 -6804
rect 1113 -6838 1147 -6804
rect 1181 -6838 1215 -6804
rect 1249 -6838 1283 -6804
rect 1317 -6838 1351 -6804
rect 1385 -6838 1419 -6804
rect 1453 -6838 1487 -6804
rect 1521 -6838 1555 -6804
rect 1589 -6838 1623 -6804
rect 1657 -6838 1691 -6804
rect 1725 -6838 1759 -6804
rect 1793 -6838 1827 -6804
rect 1861 -6838 1895 -6804
rect 1929 -6838 1963 -6804
rect 1997 -6838 2031 -6804
rect 2065 -6838 2099 -6804
rect 2133 -6838 2167 -6804
rect 2201 -6838 2235 -6804
rect 2269 -6838 2303 -6804
rect 2337 -6838 2371 -6804
rect 2405 -6838 2439 -6804
rect 2473 -6838 2507 -6804
rect 2541 -6838 2575 -6804
rect 2609 -6838 2643 -6804
rect 2677 -6838 2711 -6804
rect 2745 -6838 2779 -6804
rect 2813 -6838 2847 -6804
rect 2881 -6838 2915 -6804
rect 2949 -6838 2983 -6804
rect 3017 -6838 3051 -6804
rect 3085 -6838 3119 -6804
rect 3153 -6838 3187 -6804
rect 3221 -6838 3255 -6804
rect 3289 -6838 3323 -6804
rect 3357 -6838 3391 -6804
rect 3425 -6838 3459 -6804
rect 3493 -6838 3527 -6804
rect 3561 -6838 3595 -6804
rect 3629 -6838 3663 -6804
rect 3697 -6838 3731 -6804
rect 3765 -6838 3799 -6804
rect 3833 -6838 3867 -6804
rect 3901 -6838 3935 -6804
rect 3969 -6838 4003 -6804
rect 4037 -6838 4071 -6804
rect 4105 -6838 4139 -6804
rect 4173 -6838 4207 -6804
rect 4241 -6838 4275 -6804
rect 4309 -6838 4343 -6804
rect 4377 -6838 4411 -6804
rect 4445 -6838 4479 -6804
rect 4513 -6838 4547 -6804
rect 4581 -6838 4615 -6804
rect 4649 -6838 4683 -6804
rect 4717 -6838 4751 -6804
rect 4785 -6838 4819 -6804
rect 4853 -6838 4887 -6804
rect 4921 -6838 4955 -6804
rect 4989 -6838 5023 -6804
rect 5057 -6838 5091 -6804
rect 5372 -6838 5406 -6804
rect 5440 -6838 5474 -6804
rect 5508 -6838 5542 -6804
rect 5576 -6838 5610 -6804
rect 5644 -6838 5678 -6804
rect 5712 -6838 5746 -6804
rect 5780 -6838 5814 -6804
rect 5848 -6838 5882 -6804
rect 5916 -6838 5950 -6804
rect 5984 -6838 6018 -6804
rect 6052 -6838 6086 -6804
rect 6120 -6838 6154 -6804
rect 6188 -6838 6222 -6804
rect 6256 -6838 6290 -6804
rect 6324 -6838 6358 -6804
rect 6392 -6838 6426 -6804
rect 6460 -6838 6494 -6804
rect 6528 -6838 6562 -6804
rect 6596 -6838 6630 -6804
rect 6664 -6838 6698 -6804
rect 6732 -6838 6766 -6804
rect 6800 -6838 6834 -6804
rect 6868 -6838 6902 -6804
rect 6936 -6838 6970 -6804
rect 7004 -6838 7038 -6804
rect 7072 -6838 7106 -6804
rect 7140 -6838 7174 -6804
rect 7208 -6838 7242 -6804
rect 7276 -6838 7310 -6804
rect 7344 -6838 7378 -6804
rect 7412 -6838 7446 -6804
rect 7480 -6838 7514 -6804
rect 7548 -6838 7582 -6804
rect 7616 -6838 7650 -6804
rect 7684 -6838 7718 -6804
rect 7752 -6838 7786 -6804
rect 7820 -6838 7854 -6804
rect 7888 -6838 7922 -6804
rect 7956 -6838 7990 -6804
rect 8024 -6838 8058 -6804
rect 8092 -6838 8126 -6804
rect 8160 -6838 8194 -6804
rect 8228 -6838 8262 -6804
rect 8296 -6838 8330 -6804
rect 8364 -6838 8398 -6804
rect 8432 -6838 8466 -6804
rect 8500 -6838 8534 -6804
rect 8568 -6838 8602 -6804
rect 8636 -6838 8670 -6804
rect 8704 -6838 8738 -6804
rect 8772 -6838 8806 -6804
rect 8840 -6838 8874 -6804
rect 8908 -6838 8942 -6804
rect 8976 -6838 9010 -6804
rect 9044 -6838 9078 -6804
rect 9112 -6838 9146 -6804
rect 9180 -6838 9214 -6804
rect 9248 -6838 9282 -6804
rect 9316 -6838 9350 -6804
rect 9384 -6838 9418 -6804
rect 9452 -6838 9486 -6804
rect 9694 -6838 9728 -6804
rect 9762 -6838 9796 -6804
rect 9830 -6838 9864 -6804
rect 9898 -6838 9932 -6804
rect 9966 -6838 10000 -6804
rect 10034 -6838 10068 -6804
rect 10102 -6838 10136 -6804
rect 10170 -6838 10204 -6804
rect 10238 -6838 10272 -6804
rect 10306 -6838 10340 -6804
rect 10374 -6838 10408 -6804
rect 10442 -6838 10476 -6804
rect 10510 -6838 10544 -6804
rect 10578 -6838 10612 -6804
rect 10646 -6838 10680 -6804
rect 10714 -6838 10748 -6804
rect 10782 -6838 10816 -6804
rect 10850 -6838 10884 -6804
rect 10918 -6838 10952 -6804
rect 10986 -6838 11020 -6804
rect 11054 -6838 11088 -6804
rect 11122 -6838 11156 -6804
rect 11190 -6838 11224 -6804
rect 11258 -6838 11292 -6804
rect 11326 -6838 11360 -6804
rect 11394 -6838 11428 -6804
rect 11462 -6838 11496 -6804
rect 11530 -6838 11564 -6804
rect 11598 -6838 11632 -6804
rect 11666 -6838 11700 -6804
rect 11734 -6838 11768 -6804
rect 11802 -6838 11836 -6804
rect 11870 -6838 11904 -6804
rect 11938 -6838 11972 -6804
rect 12006 -6838 12040 -6804
rect 12074 -6838 12108 -6804
rect 12142 -6838 12176 -6804
rect 12210 -6838 12244 -6804
rect 12278 -6838 12312 -6804
rect 12346 -6838 12380 -6804
rect 12414 -6838 12448 -6804
rect 12482 -6838 12516 -6804
rect 12550 -6838 12584 -6804
rect 12618 -6838 12652 -6804
rect 12686 -6838 12720 -6804
rect 12754 -6838 12788 -6804
rect 12822 -6838 12856 -6804
rect 12890 -6838 12924 -6804
rect 12958 -6838 12992 -6804
rect 13026 -6838 13060 -6804
rect 13094 -6838 13128 -6804
rect 13162 -6838 13196 -6804
rect 13230 -6838 13264 -6804
rect 13298 -6838 13332 -6804
rect 13366 -6838 13400 -6804
rect 13434 -6838 13468 -6804
rect 13502 -6838 13536 -6804
rect 13570 -6838 13604 -6804
rect 13638 -6838 13672 -6804
rect 13706 -6838 13740 -6804
rect 13774 -6838 13808 -6804
rect 14089 -6838 14123 -6804
rect 14157 -6838 14191 -6804
rect 14225 -6838 14259 -6804
rect 14293 -6838 14327 -6804
rect 14361 -6838 14395 -6804
rect 14429 -6838 14463 -6804
rect 14497 -6838 14531 -6804
rect 14565 -6838 14599 -6804
rect 14633 -6838 14667 -6804
rect 14701 -6838 14735 -6804
rect 14769 -6838 14803 -6804
rect 14837 -6838 14871 -6804
rect 14905 -6838 14939 -6804
rect 14973 -6838 15007 -6804
rect 15041 -6838 15075 -6804
rect 15109 -6838 15143 -6804
rect 15177 -6838 15211 -6804
rect 15245 -6838 15279 -6804
rect 15313 -6838 15347 -6804
rect 15381 -6838 15415 -6804
rect 15449 -6838 15483 -6804
rect 15517 -6838 15551 -6804
rect 15585 -6838 15619 -6804
rect 15653 -6838 15687 -6804
rect 15721 -6838 15755 -6804
rect 15789 -6838 15823 -6804
rect 15857 -6838 15891 -6804
rect 15925 -6838 15959 -6804
rect 15993 -6838 16027 -6804
rect 16061 -6838 16095 -6804
rect 16129 -6838 16163 -6804
rect 16197 -6838 16231 -6804
rect 16265 -6838 16299 -6804
rect 16333 -6838 16367 -6804
rect 16401 -6838 16435 -6804
rect 16469 -6838 16503 -6804
rect 16537 -6838 16571 -6804
rect 16605 -6838 16639 -6804
rect 16673 -6838 16707 -6804
rect 16741 -6838 16775 -6804
rect 16809 -6838 16843 -6804
rect 16877 -6838 16911 -6804
rect 16945 -6838 16979 -6804
rect 17013 -6838 17047 -6804
rect 17081 -6838 17115 -6804
rect 17149 -6838 17183 -6804
rect 17217 -6838 17251 -6804
rect 17285 -6838 17319 -6804
rect 17353 -6838 17387 -6804
rect 17421 -6838 17455 -6804
rect 17489 -6838 17523 -6804
rect 17557 -6838 17591 -6804
rect 17625 -6838 17659 -6804
rect 17693 -6838 17727 -6804
rect 17761 -6838 17795 -6804
rect 17829 -6838 17863 -6804
rect 17897 -6838 17931 -6804
rect 17965 -6838 17999 -6804
rect 18033 -6838 18067 -6804
rect 18101 -6838 18135 -6804
rect 18169 -6838 18203 -6804
rect 856 -6974 890 -6940
rect 856 -7042 890 -7008
rect 856 -7110 890 -7076
rect 856 -7178 890 -7144
rect 5214 -6974 5248 -6940
rect 5214 -7042 5248 -7008
rect 5214 -7110 5248 -7076
rect 5214 -7178 5248 -7144
rect 9573 -6974 9607 -6940
rect 9573 -7042 9607 -7008
rect 9573 -7110 9607 -7076
rect 856 -7246 890 -7212
rect 856 -7314 890 -7280
rect 856 -7382 890 -7348
rect 9573 -7178 9607 -7144
rect 13932 -6974 13966 -6940
rect 13932 -7042 13966 -7008
rect 13932 -7110 13966 -7076
rect 5214 -7246 5248 -7212
rect 5214 -7314 5248 -7280
rect 5214 -7382 5248 -7348
rect 856 -7450 890 -7416
rect 856 -7518 890 -7484
rect 13932 -7178 13966 -7144
rect 18290 -6974 18324 -6940
rect 18290 -7042 18324 -7008
rect 18290 -7110 18324 -7076
rect 9573 -7246 9607 -7212
rect 9573 -7314 9607 -7280
rect 9573 -7382 9607 -7348
rect 5214 -7450 5248 -7416
rect 856 -7586 890 -7552
rect 856 -7654 890 -7620
rect 856 -7722 890 -7688
rect 856 -7790 890 -7756
rect 5214 -7518 5248 -7484
rect 18290 -7178 18324 -7144
rect 13932 -7246 13966 -7212
rect 13932 -7314 13966 -7280
rect 13932 -7382 13966 -7348
rect 9573 -7450 9607 -7416
rect 5214 -7586 5248 -7552
rect 5214 -7654 5248 -7620
rect 5214 -7722 5248 -7688
rect 5214 -7790 5248 -7756
rect 9573 -7518 9607 -7484
rect 18290 -7246 18324 -7212
rect 18290 -7314 18324 -7280
rect 18290 -7382 18324 -7348
rect 13932 -7450 13966 -7416
rect 9573 -7586 9607 -7552
rect 9573 -7654 9607 -7620
rect 9573 -7722 9607 -7688
rect 9573 -7790 9607 -7756
rect 13932 -7518 13966 -7484
rect 18290 -7450 18324 -7416
rect 13932 -7586 13966 -7552
rect 13932 -7654 13966 -7620
rect 13932 -7722 13966 -7688
rect 13932 -7790 13966 -7756
rect 18290 -7518 18324 -7484
rect 18290 -7586 18324 -7552
rect 18290 -7654 18324 -7620
rect 18290 -7722 18324 -7688
rect 18290 -7790 18324 -7756
rect 856 -7858 890 -7824
rect 5214 -7858 5248 -7824
rect 856 -7926 890 -7892
rect 856 -7994 890 -7960
rect 856 -8062 890 -8028
rect 9573 -7858 9607 -7824
rect 5214 -7926 5248 -7892
rect 5214 -7994 5248 -7960
rect 5214 -8062 5248 -8028
rect 856 -8130 890 -8096
rect 13932 -7858 13966 -7824
rect 9573 -7926 9607 -7892
rect 9573 -7994 9607 -7960
rect 9573 -8062 9607 -8028
rect 856 -8198 890 -8164
rect 856 -8266 890 -8232
rect 856 -8334 890 -8300
rect 856 -8402 890 -8368
rect 5214 -8130 5248 -8096
rect 18290 -7858 18324 -7824
rect 13932 -7926 13966 -7892
rect 13932 -7994 13966 -7960
rect 13932 -8062 13966 -8028
rect 5214 -8198 5248 -8164
rect 5214 -8266 5248 -8232
rect 5214 -8334 5248 -8300
rect 5214 -8402 5248 -8368
rect 9573 -8130 9607 -8096
rect 18290 -7926 18324 -7892
rect 18290 -7994 18324 -7960
rect 18290 -8062 18324 -8028
rect 9573 -8198 9607 -8164
rect 9573 -8266 9607 -8232
rect 9573 -8334 9607 -8300
rect 9573 -8402 9607 -8368
rect 13932 -8130 13966 -8096
rect 13932 -8198 13966 -8164
rect 13932 -8266 13966 -8232
rect 13932 -8334 13966 -8300
rect 13932 -8402 13966 -8368
rect 18290 -8130 18324 -8096
rect 18290 -8198 18324 -8164
rect 18290 -8266 18324 -8232
rect 18290 -8334 18324 -8300
rect 18290 -8402 18324 -8368
rect 977 -8436 1011 -8402
rect 1045 -8436 1079 -8402
rect 1113 -8436 1147 -8402
rect 1181 -8436 1215 -8402
rect 1249 -8436 1283 -8402
rect 1317 -8436 1351 -8402
rect 1385 -8436 1419 -8402
rect 1453 -8436 1487 -8402
rect 1521 -8436 1555 -8402
rect 1589 -8436 1623 -8402
rect 1657 -8436 1691 -8402
rect 1725 -8436 1759 -8402
rect 1793 -8436 1827 -8402
rect 1861 -8436 1895 -8402
rect 1929 -8436 1963 -8402
rect 1997 -8436 2031 -8402
rect 2065 -8436 2099 -8402
rect 2133 -8436 2167 -8402
rect 2201 -8436 2235 -8402
rect 2269 -8436 2303 -8402
rect 2337 -8436 2371 -8402
rect 2405 -8436 2439 -8402
rect 2473 -8436 2507 -8402
rect 2541 -8436 2575 -8402
rect 2609 -8436 2643 -8402
rect 2677 -8436 2711 -8402
rect 2745 -8436 2779 -8402
rect 2813 -8436 2847 -8402
rect 2881 -8436 2915 -8402
rect 2949 -8436 2983 -8402
rect 3017 -8436 3051 -8402
rect 3085 -8436 3119 -8402
rect 3153 -8436 3187 -8402
rect 3221 -8436 3255 -8402
rect 3289 -8436 3323 -8402
rect 3357 -8436 3391 -8402
rect 3425 -8436 3459 -8402
rect 3493 -8436 3527 -8402
rect 3561 -8436 3595 -8402
rect 3629 -8436 3663 -8402
rect 3697 -8436 3731 -8402
rect 3765 -8436 3799 -8402
rect 3833 -8436 3867 -8402
rect 3901 -8436 3935 -8402
rect 3969 -8436 4003 -8402
rect 4037 -8436 4071 -8402
rect 4105 -8436 4139 -8402
rect 4173 -8436 4207 -8402
rect 4241 -8436 4275 -8402
rect 4309 -8436 4343 -8402
rect 4377 -8436 4411 -8402
rect 4445 -8436 4479 -8402
rect 4513 -8436 4547 -8402
rect 4581 -8436 4615 -8402
rect 4649 -8436 4683 -8402
rect 4717 -8436 4751 -8402
rect 4785 -8436 4819 -8402
rect 4853 -8436 4887 -8402
rect 4921 -8436 4955 -8402
rect 4989 -8436 5023 -8402
rect 5057 -8436 5091 -8402
rect 5372 -8436 5406 -8402
rect 5440 -8436 5474 -8402
rect 5508 -8436 5542 -8402
rect 5576 -8436 5610 -8402
rect 5644 -8436 5678 -8402
rect 5712 -8436 5746 -8402
rect 5780 -8436 5814 -8402
rect 5848 -8436 5882 -8402
rect 5916 -8436 5950 -8402
rect 5984 -8436 6018 -8402
rect 6052 -8436 6086 -8402
rect 6120 -8436 6154 -8402
rect 6188 -8436 6222 -8402
rect 6256 -8436 6290 -8402
rect 6324 -8436 6358 -8402
rect 6392 -8436 6426 -8402
rect 6460 -8436 6494 -8402
rect 6528 -8436 6562 -8402
rect 6596 -8436 6630 -8402
rect 6664 -8436 6698 -8402
rect 6732 -8436 6766 -8402
rect 6800 -8436 6834 -8402
rect 6868 -8436 6902 -8402
rect 6936 -8436 6970 -8402
rect 7004 -8436 7038 -8402
rect 7072 -8436 7106 -8402
rect 7140 -8436 7174 -8402
rect 7208 -8436 7242 -8402
rect 7276 -8436 7310 -8402
rect 7344 -8436 7378 -8402
rect 7412 -8436 7446 -8402
rect 7480 -8436 7514 -8402
rect 7548 -8436 7582 -8402
rect 7616 -8436 7650 -8402
rect 7684 -8436 7718 -8402
rect 7752 -8436 7786 -8402
rect 7820 -8436 7854 -8402
rect 7888 -8436 7922 -8402
rect 7956 -8436 7990 -8402
rect 8024 -8436 8058 -8402
rect 8092 -8436 8126 -8402
rect 8160 -8436 8194 -8402
rect 8228 -8436 8262 -8402
rect 8296 -8436 8330 -8402
rect 8364 -8436 8398 -8402
rect 8432 -8436 8466 -8402
rect 8500 -8436 8534 -8402
rect 8568 -8436 8602 -8402
rect 8636 -8436 8670 -8402
rect 8704 -8436 8738 -8402
rect 8772 -8436 8806 -8402
rect 8840 -8436 8874 -8402
rect 8908 -8436 8942 -8402
rect 8976 -8436 9010 -8402
rect 9044 -8436 9078 -8402
rect 9112 -8436 9146 -8402
rect 9180 -8436 9214 -8402
rect 9248 -8436 9282 -8402
rect 9316 -8436 9350 -8402
rect 9384 -8436 9418 -8402
rect 9452 -8436 9486 -8402
rect 9694 -8436 9728 -8402
rect 9762 -8436 9796 -8402
rect 9830 -8436 9864 -8402
rect 9898 -8436 9932 -8402
rect 9966 -8436 10000 -8402
rect 10034 -8436 10068 -8402
rect 10102 -8436 10136 -8402
rect 10170 -8436 10204 -8402
rect 10238 -8436 10272 -8402
rect 10306 -8436 10340 -8402
rect 10374 -8436 10408 -8402
rect 10442 -8436 10476 -8402
rect 10510 -8436 10544 -8402
rect 10578 -8436 10612 -8402
rect 10646 -8436 10680 -8402
rect 10714 -8436 10748 -8402
rect 10782 -8436 10816 -8402
rect 10850 -8436 10884 -8402
rect 10918 -8436 10952 -8402
rect 10986 -8436 11020 -8402
rect 11054 -8436 11088 -8402
rect 11122 -8436 11156 -8402
rect 11190 -8436 11224 -8402
rect 11258 -8436 11292 -8402
rect 11326 -8436 11360 -8402
rect 11394 -8436 11428 -8402
rect 11462 -8436 11496 -8402
rect 11530 -8436 11564 -8402
rect 11598 -8436 11632 -8402
rect 11666 -8436 11700 -8402
rect 11734 -8436 11768 -8402
rect 11802 -8436 11836 -8402
rect 11870 -8436 11904 -8402
rect 11938 -8436 11972 -8402
rect 12006 -8436 12040 -8402
rect 12074 -8436 12108 -8402
rect 12142 -8436 12176 -8402
rect 12210 -8436 12244 -8402
rect 12278 -8436 12312 -8402
rect 12346 -8436 12380 -8402
rect 12414 -8436 12448 -8402
rect 12482 -8436 12516 -8402
rect 12550 -8436 12584 -8402
rect 12618 -8436 12652 -8402
rect 12686 -8436 12720 -8402
rect 12754 -8436 12788 -8402
rect 12822 -8436 12856 -8402
rect 12890 -8436 12924 -8402
rect 12958 -8436 12992 -8402
rect 13026 -8436 13060 -8402
rect 13094 -8436 13128 -8402
rect 13162 -8436 13196 -8402
rect 13230 -8436 13264 -8402
rect 13298 -8436 13332 -8402
rect 13366 -8436 13400 -8402
rect 13434 -8436 13468 -8402
rect 13502 -8436 13536 -8402
rect 13570 -8436 13604 -8402
rect 13638 -8436 13672 -8402
rect 13706 -8436 13740 -8402
rect 13774 -8436 13808 -8402
rect 14089 -8436 14123 -8402
rect 14157 -8436 14191 -8402
rect 14225 -8436 14259 -8402
rect 14293 -8436 14327 -8402
rect 14361 -8436 14395 -8402
rect 14429 -8436 14463 -8402
rect 14497 -8436 14531 -8402
rect 14565 -8436 14599 -8402
rect 14633 -8436 14667 -8402
rect 14701 -8436 14735 -8402
rect 14769 -8436 14803 -8402
rect 14837 -8436 14871 -8402
rect 14905 -8436 14939 -8402
rect 14973 -8436 15007 -8402
rect 15041 -8436 15075 -8402
rect 15109 -8436 15143 -8402
rect 15177 -8436 15211 -8402
rect 15245 -8436 15279 -8402
rect 15313 -8436 15347 -8402
rect 15381 -8436 15415 -8402
rect 15449 -8436 15483 -8402
rect 15517 -8436 15551 -8402
rect 15585 -8436 15619 -8402
rect 15653 -8436 15687 -8402
rect 15721 -8436 15755 -8402
rect 15789 -8436 15823 -8402
rect 15857 -8436 15891 -8402
rect 15925 -8436 15959 -8402
rect 15993 -8436 16027 -8402
rect 16061 -8436 16095 -8402
rect 16129 -8436 16163 -8402
rect 16197 -8436 16231 -8402
rect 16265 -8436 16299 -8402
rect 16333 -8436 16367 -8402
rect 16401 -8436 16435 -8402
rect 16469 -8436 16503 -8402
rect 16537 -8436 16571 -8402
rect 16605 -8436 16639 -8402
rect 16673 -8436 16707 -8402
rect 16741 -8436 16775 -8402
rect 16809 -8436 16843 -8402
rect 16877 -8436 16911 -8402
rect 16945 -8436 16979 -8402
rect 17013 -8436 17047 -8402
rect 17081 -8436 17115 -8402
rect 17149 -8436 17183 -8402
rect 17217 -8436 17251 -8402
rect 17285 -8436 17319 -8402
rect 17353 -8436 17387 -8402
rect 17421 -8436 17455 -8402
rect 17489 -8436 17523 -8402
rect 17557 -8436 17591 -8402
rect 17625 -8436 17659 -8402
rect 17693 -8436 17727 -8402
rect 17761 -8436 17795 -8402
rect 17829 -8436 17863 -8402
rect 17897 -8436 17931 -8402
rect 17965 -8436 17999 -8402
rect 18033 -8436 18067 -8402
rect 18101 -8436 18135 -8402
rect 18169 -8436 18203 -8402
rect 856 -8470 890 -8436
rect 856 -8538 890 -8504
rect 856 -8606 890 -8572
rect 856 -8674 890 -8640
rect 856 -8742 890 -8708
rect 856 -8810 890 -8776
rect 5214 -8470 5248 -8436
rect 5214 -8538 5248 -8504
rect 5214 -8606 5248 -8572
rect 5214 -8674 5248 -8640
rect 5214 -8742 5248 -8708
rect 5214 -8810 5248 -8776
rect 9573 -8470 9607 -8436
rect 9573 -8538 9607 -8504
rect 9573 -8606 9607 -8572
rect 9573 -8674 9607 -8640
rect 9573 -8742 9607 -8708
rect 856 -8878 890 -8844
rect 856 -8946 890 -8912
rect 856 -9014 890 -8980
rect 9573 -8810 9607 -8776
rect 13932 -8470 13966 -8436
rect 13932 -8538 13966 -8504
rect 13932 -8606 13966 -8572
rect 13932 -8674 13966 -8640
rect 13932 -8742 13966 -8708
rect 5214 -8878 5248 -8844
rect 5214 -8946 5248 -8912
rect 5214 -9014 5248 -8980
rect 13932 -8810 13966 -8776
rect 18290 -8470 18324 -8436
rect 18290 -8538 18324 -8504
rect 18290 -8606 18324 -8572
rect 18290 -8674 18324 -8640
rect 18290 -8742 18324 -8708
rect 9573 -8878 9607 -8844
rect 9573 -8946 9607 -8912
rect 9573 -9014 9607 -8980
rect 18290 -8810 18324 -8776
rect 13932 -8878 13966 -8844
rect 13932 -8946 13966 -8912
rect 13932 -9014 13966 -8980
rect 18290 -8878 18324 -8844
rect 18290 -8946 18324 -8912
rect 18290 -9014 18324 -8980
rect 977 -9226 1011 -9192
rect 1045 -9226 1079 -9192
rect 1113 -9226 1147 -9192
rect 1181 -9226 1215 -9192
rect 1249 -9226 1283 -9192
rect 1317 -9226 1351 -9192
rect 1385 -9226 1419 -9192
rect 1453 -9226 1487 -9192
rect 1521 -9226 1555 -9192
rect 1589 -9226 1623 -9192
rect 1657 -9226 1691 -9192
rect 1725 -9226 1759 -9192
rect 1793 -9226 1827 -9192
rect 1861 -9226 1895 -9192
rect 1929 -9226 1963 -9192
rect 1997 -9226 2031 -9192
rect 2065 -9226 2099 -9192
rect 2133 -9226 2167 -9192
rect 2201 -9226 2235 -9192
rect 2269 -9226 2303 -9192
rect 2337 -9226 2371 -9192
rect 2405 -9226 2439 -9192
rect 2473 -9226 2507 -9192
rect 2541 -9226 2575 -9192
rect 2609 -9226 2643 -9192
rect 2677 -9226 2711 -9192
rect 2745 -9226 2779 -9192
rect 2813 -9226 2847 -9192
rect 2881 -9226 2915 -9192
rect 2949 -9226 2983 -9192
rect 3017 -9226 3051 -9192
rect 3085 -9226 3119 -9192
rect 3153 -9226 3187 -9192
rect 3221 -9226 3255 -9192
rect 3289 -9226 3323 -9192
rect 3357 -9226 3391 -9192
rect 3425 -9226 3459 -9192
rect 3493 -9226 3527 -9192
rect 3561 -9226 3595 -9192
rect 3629 -9226 3663 -9192
rect 3697 -9226 3731 -9192
rect 3765 -9226 3799 -9192
rect 3833 -9226 3867 -9192
rect 3901 -9226 3935 -9192
rect 3969 -9226 4003 -9192
rect 4037 -9226 4071 -9192
rect 4105 -9226 4139 -9192
rect 4173 -9226 4207 -9192
rect 4241 -9226 4275 -9192
rect 4309 -9226 4343 -9192
rect 4377 -9226 4411 -9192
rect 4445 -9226 4479 -9192
rect 4513 -9226 4547 -9192
rect 4581 -9226 4615 -9192
rect 4649 -9226 4683 -9192
rect 4717 -9226 4751 -9192
rect 4785 -9226 4819 -9192
rect 4853 -9226 4887 -9192
rect 4921 -9226 4955 -9192
rect 4989 -9226 5023 -9192
rect 5057 -9226 5091 -9192
rect 5372 -9226 5406 -9192
rect 5440 -9226 5474 -9192
rect 5508 -9226 5542 -9192
rect 5576 -9226 5610 -9192
rect 5644 -9226 5678 -9192
rect 5712 -9226 5746 -9192
rect 5780 -9226 5814 -9192
rect 5848 -9226 5882 -9192
rect 5916 -9226 5950 -9192
rect 5984 -9226 6018 -9192
rect 6052 -9226 6086 -9192
rect 6120 -9226 6154 -9192
rect 6188 -9226 6222 -9192
rect 6256 -9226 6290 -9192
rect 6324 -9226 6358 -9192
rect 6392 -9226 6426 -9192
rect 6460 -9226 6494 -9192
rect 6528 -9226 6562 -9192
rect 6596 -9226 6630 -9192
rect 6664 -9226 6698 -9192
rect 6732 -9226 6766 -9192
rect 6800 -9226 6834 -9192
rect 6868 -9226 6902 -9192
rect 6936 -9226 6970 -9192
rect 7004 -9226 7038 -9192
rect 7072 -9226 7106 -9192
rect 7140 -9226 7174 -9192
rect 7208 -9226 7242 -9192
rect 7276 -9226 7310 -9192
rect 7344 -9226 7378 -9192
rect 7412 -9226 7446 -9192
rect 7480 -9226 7514 -9192
rect 7548 -9226 7582 -9192
rect 7616 -9226 7650 -9192
rect 7684 -9226 7718 -9192
rect 7752 -9226 7786 -9192
rect 7820 -9226 7854 -9192
rect 7888 -9226 7922 -9192
rect 7956 -9226 7990 -9192
rect 8024 -9226 8058 -9192
rect 8092 -9226 8126 -9192
rect 8160 -9226 8194 -9192
rect 8228 -9226 8262 -9192
rect 8296 -9226 8330 -9192
rect 8364 -9226 8398 -9192
rect 8432 -9226 8466 -9192
rect 8500 -9226 8534 -9192
rect 8568 -9226 8602 -9192
rect 8636 -9226 8670 -9192
rect 8704 -9226 8738 -9192
rect 8772 -9226 8806 -9192
rect 8840 -9226 8874 -9192
rect 8908 -9226 8942 -9192
rect 8976 -9226 9010 -9192
rect 9044 -9226 9078 -9192
rect 9112 -9226 9146 -9192
rect 9180 -9226 9214 -9192
rect 9248 -9226 9282 -9192
rect 9316 -9226 9350 -9192
rect 9384 -9226 9418 -9192
rect 9452 -9226 9486 -9192
rect 9694 -9226 9728 -9192
rect 9762 -9226 9796 -9192
rect 9830 -9226 9864 -9192
rect 9898 -9226 9932 -9192
rect 9966 -9226 10000 -9192
rect 10034 -9226 10068 -9192
rect 10102 -9226 10136 -9192
rect 10170 -9226 10204 -9192
rect 10238 -9226 10272 -9192
rect 10306 -9226 10340 -9192
rect 10374 -9226 10408 -9192
rect 10442 -9226 10476 -9192
rect 10510 -9226 10544 -9192
rect 10578 -9226 10612 -9192
rect 10646 -9226 10680 -9192
rect 10714 -9226 10748 -9192
rect 10782 -9226 10816 -9192
rect 10850 -9226 10884 -9192
rect 10918 -9226 10952 -9192
rect 10986 -9226 11020 -9192
rect 11054 -9226 11088 -9192
rect 11122 -9226 11156 -9192
rect 11190 -9226 11224 -9192
rect 11258 -9226 11292 -9192
rect 11326 -9226 11360 -9192
rect 11394 -9226 11428 -9192
rect 11462 -9226 11496 -9192
rect 11530 -9226 11564 -9192
rect 11598 -9226 11632 -9192
rect 11666 -9226 11700 -9192
rect 11734 -9226 11768 -9192
rect 11802 -9226 11836 -9192
rect 11870 -9226 11904 -9192
rect 11938 -9226 11972 -9192
rect 12006 -9226 12040 -9192
rect 12074 -9226 12108 -9192
rect 12142 -9226 12176 -9192
rect 12210 -9226 12244 -9192
rect 12278 -9226 12312 -9192
rect 12346 -9226 12380 -9192
rect 12414 -9226 12448 -9192
rect 12482 -9226 12516 -9192
rect 12550 -9226 12584 -9192
rect 12618 -9226 12652 -9192
rect 12686 -9226 12720 -9192
rect 12754 -9226 12788 -9192
rect 12822 -9226 12856 -9192
rect 12890 -9226 12924 -9192
rect 12958 -9226 12992 -9192
rect 13026 -9226 13060 -9192
rect 13094 -9226 13128 -9192
rect 13162 -9226 13196 -9192
rect 13230 -9226 13264 -9192
rect 13298 -9226 13332 -9192
rect 13366 -9226 13400 -9192
rect 13434 -9226 13468 -9192
rect 13502 -9226 13536 -9192
rect 13570 -9226 13604 -9192
rect 13638 -9226 13672 -9192
rect 13706 -9226 13740 -9192
rect 13774 -9226 13808 -9192
rect 14089 -9226 14123 -9192
rect 14157 -9226 14191 -9192
rect 14225 -9226 14259 -9192
rect 14293 -9226 14327 -9192
rect 14361 -9226 14395 -9192
rect 14429 -9226 14463 -9192
rect 14497 -9226 14531 -9192
rect 14565 -9226 14599 -9192
rect 14633 -9226 14667 -9192
rect 14701 -9226 14735 -9192
rect 14769 -9226 14803 -9192
rect 14837 -9226 14871 -9192
rect 14905 -9226 14939 -9192
rect 14973 -9226 15007 -9192
rect 15041 -9226 15075 -9192
rect 15109 -9226 15143 -9192
rect 15177 -9226 15211 -9192
rect 15245 -9226 15279 -9192
rect 15313 -9226 15347 -9192
rect 15381 -9226 15415 -9192
rect 15449 -9226 15483 -9192
rect 15517 -9226 15551 -9192
rect 15585 -9226 15619 -9192
rect 15653 -9226 15687 -9192
rect 15721 -9226 15755 -9192
rect 15789 -9226 15823 -9192
rect 15857 -9226 15891 -9192
rect 15925 -9226 15959 -9192
rect 15993 -9226 16027 -9192
rect 16061 -9226 16095 -9192
rect 16129 -9226 16163 -9192
rect 16197 -9226 16231 -9192
rect 16265 -9226 16299 -9192
rect 16333 -9226 16367 -9192
rect 16401 -9226 16435 -9192
rect 16469 -9226 16503 -9192
rect 16537 -9226 16571 -9192
rect 16605 -9226 16639 -9192
rect 16673 -9226 16707 -9192
rect 16741 -9226 16775 -9192
rect 16809 -9226 16843 -9192
rect 16877 -9226 16911 -9192
rect 16945 -9226 16979 -9192
rect 17013 -9226 17047 -9192
rect 17081 -9226 17115 -9192
rect 17149 -9226 17183 -9192
rect 17217 -9226 17251 -9192
rect 17285 -9226 17319 -9192
rect 17353 -9226 17387 -9192
rect 17421 -9226 17455 -9192
rect 17489 -9226 17523 -9192
rect 17557 -9226 17591 -9192
rect 17625 -9226 17659 -9192
rect 17693 -9226 17727 -9192
rect 17761 -9226 17795 -9192
rect 17829 -9226 17863 -9192
rect 17897 -9226 17931 -9192
rect 17965 -9226 17999 -9192
rect 18033 -9226 18067 -9192
rect 18101 -9226 18135 -9192
rect 18169 -9226 18203 -9192
<< poly >>
rect 1017 349 1217 365
rect 1017 315 1066 349
rect 1100 315 1134 349
rect 1168 315 1217 349
rect 1017 268 1217 315
rect 1469 349 1669 365
rect 1469 315 1518 349
rect 1552 315 1586 349
rect 1620 315 1669 349
rect 1469 268 1669 315
rect 1727 349 1927 365
rect 1727 315 1776 349
rect 1810 315 1844 349
rect 1878 315 1927 349
rect 1727 268 1927 315
rect 1985 349 2185 365
rect 1985 315 2034 349
rect 2068 315 2102 349
rect 2136 315 2185 349
rect 1985 268 2185 315
rect 2243 349 2443 365
rect 2243 315 2292 349
rect 2326 315 2360 349
rect 2394 315 2443 349
rect 2243 268 2443 315
rect 2695 349 2895 365
rect 2695 315 2744 349
rect 2778 315 2812 349
rect 2846 315 2895 349
rect 2695 268 2895 315
rect 2953 349 3153 365
rect 2953 315 3002 349
rect 3036 315 3070 349
rect 3104 315 3153 349
rect 2953 268 3153 315
rect 3211 349 3411 365
rect 3211 315 3260 349
rect 3294 315 3328 349
rect 3362 315 3411 349
rect 3211 268 3411 315
rect 3663 349 3863 365
rect 3663 315 3712 349
rect 3746 315 3780 349
rect 3814 315 3863 349
rect 3663 268 3863 315
rect 3921 349 4121 365
rect 3921 315 3970 349
rect 4004 315 4038 349
rect 4072 315 4121 349
rect 3921 268 4121 315
rect 4179 349 4379 365
rect 4179 315 4228 349
rect 4262 315 4296 349
rect 4330 315 4379 349
rect 4179 268 4379 315
rect 4437 349 4637 365
rect 4437 315 4486 349
rect 4520 315 4554 349
rect 4588 315 4637 349
rect 4437 268 4637 315
rect 4888 349 5088 365
rect 4888 315 4937 349
rect 4971 315 5005 349
rect 5039 315 5088 349
rect 4888 268 5088 315
rect 5374 349 5574 365
rect 5374 315 5423 349
rect 5457 315 5491 349
rect 5525 315 5574 349
rect 5374 268 5574 315
rect 5826 349 6026 365
rect 5826 315 5875 349
rect 5909 315 5943 349
rect 5977 315 6026 349
rect 5826 268 6026 315
rect 6084 349 6284 365
rect 6084 315 6133 349
rect 6167 315 6201 349
rect 6235 315 6284 349
rect 6084 268 6284 315
rect 6342 349 6542 365
rect 6342 315 6391 349
rect 6425 315 6459 349
rect 6493 315 6542 349
rect 6342 268 6542 315
rect 6600 349 6800 365
rect 6600 315 6649 349
rect 6683 315 6717 349
rect 6751 315 6800 349
rect 6600 268 6800 315
rect 7052 349 7252 365
rect 7052 315 7101 349
rect 7135 315 7169 349
rect 7203 315 7252 349
rect 7052 268 7252 315
rect 7310 349 7510 365
rect 7310 315 7359 349
rect 7393 315 7427 349
rect 7461 315 7510 349
rect 7310 268 7510 315
rect 7568 349 7768 365
rect 7568 315 7617 349
rect 7651 315 7685 349
rect 7719 315 7768 349
rect 7568 268 7768 315
rect 8020 349 8220 365
rect 8020 315 8069 349
rect 8103 315 8137 349
rect 8171 315 8220 349
rect 8020 268 8220 315
rect 8278 349 8478 365
rect 8278 315 8327 349
rect 8361 315 8395 349
rect 8429 315 8478 349
rect 8278 268 8478 315
rect 8536 349 8736 365
rect 8536 315 8585 349
rect 8619 315 8653 349
rect 8687 315 8736 349
rect 8536 268 8736 315
rect 8794 349 8994 365
rect 8794 315 8843 349
rect 8877 315 8911 349
rect 8945 315 8994 349
rect 8794 268 8994 315
rect 9246 349 9446 365
rect 9246 315 9295 349
rect 9329 315 9363 349
rect 9397 315 9446 349
rect 9246 268 9446 315
rect 1017 42 1217 68
rect 1469 42 1669 68
rect 1727 42 1927 68
rect 1985 42 2185 68
rect 2243 42 2443 68
rect 2695 42 2895 68
rect 2953 42 3153 68
rect 3211 42 3411 68
rect 3663 42 3863 68
rect 3921 42 4121 68
rect 4179 42 4379 68
rect 4437 42 4637 68
rect 4888 42 5088 68
rect 9734 349 9934 365
rect 9734 315 9783 349
rect 9817 315 9851 349
rect 9885 315 9934 349
rect 9734 268 9934 315
rect 10186 349 10386 365
rect 10186 315 10235 349
rect 10269 315 10303 349
rect 10337 315 10386 349
rect 10186 268 10386 315
rect 10444 349 10644 365
rect 10444 315 10493 349
rect 10527 315 10561 349
rect 10595 315 10644 349
rect 10444 268 10644 315
rect 10702 349 10902 365
rect 10702 315 10751 349
rect 10785 315 10819 349
rect 10853 315 10902 349
rect 10702 268 10902 315
rect 10960 349 11160 365
rect 10960 315 11009 349
rect 11043 315 11077 349
rect 11111 315 11160 349
rect 10960 268 11160 315
rect 11412 349 11612 365
rect 11412 315 11461 349
rect 11495 315 11529 349
rect 11563 315 11612 349
rect 11412 268 11612 315
rect 11670 349 11870 365
rect 11670 315 11719 349
rect 11753 315 11787 349
rect 11821 315 11870 349
rect 11670 268 11870 315
rect 11928 349 12128 365
rect 11928 315 11977 349
rect 12011 315 12045 349
rect 12079 315 12128 349
rect 11928 268 12128 315
rect 12380 349 12580 365
rect 12380 315 12429 349
rect 12463 315 12497 349
rect 12531 315 12580 349
rect 12380 268 12580 315
rect 12638 349 12838 365
rect 12638 315 12687 349
rect 12721 315 12755 349
rect 12789 315 12838 349
rect 12638 268 12838 315
rect 12896 349 13096 365
rect 12896 315 12945 349
rect 12979 315 13013 349
rect 13047 315 13096 349
rect 12896 268 13096 315
rect 13154 349 13354 365
rect 13154 315 13203 349
rect 13237 315 13271 349
rect 13305 315 13354 349
rect 13154 268 13354 315
rect 13606 349 13806 365
rect 13606 315 13655 349
rect 13689 315 13723 349
rect 13757 315 13806 349
rect 13606 268 13806 315
rect 5374 42 5574 68
rect 5826 42 6026 68
rect 6084 42 6284 68
rect 6342 42 6542 68
rect 6600 42 6800 68
rect 7052 42 7252 68
rect 7310 42 7510 68
rect 7568 42 7768 68
rect 8020 42 8220 68
rect 8278 42 8478 68
rect 8536 42 8736 68
rect 8794 42 8994 68
rect 9246 42 9446 68
rect 14092 349 14292 365
rect 14092 315 14141 349
rect 14175 315 14209 349
rect 14243 315 14292 349
rect 14092 268 14292 315
rect 14543 349 14743 365
rect 14543 315 14592 349
rect 14626 315 14660 349
rect 14694 315 14743 349
rect 14543 268 14743 315
rect 14801 349 15001 365
rect 14801 315 14850 349
rect 14884 315 14918 349
rect 14952 315 15001 349
rect 14801 268 15001 315
rect 15059 349 15259 365
rect 15059 315 15108 349
rect 15142 315 15176 349
rect 15210 315 15259 349
rect 15059 268 15259 315
rect 15317 349 15517 365
rect 15317 315 15366 349
rect 15400 315 15434 349
rect 15468 315 15517 349
rect 15317 268 15517 315
rect 15769 349 15969 365
rect 15769 315 15818 349
rect 15852 315 15886 349
rect 15920 315 15969 349
rect 15769 268 15969 315
rect 16027 349 16227 365
rect 16027 315 16076 349
rect 16110 315 16144 349
rect 16178 315 16227 349
rect 16027 268 16227 315
rect 16285 349 16485 365
rect 16285 315 16334 349
rect 16368 315 16402 349
rect 16436 315 16485 349
rect 16285 268 16485 315
rect 16737 349 16937 365
rect 16737 315 16786 349
rect 16820 315 16854 349
rect 16888 315 16937 349
rect 16737 268 16937 315
rect 16995 349 17195 365
rect 16995 315 17044 349
rect 17078 315 17112 349
rect 17146 315 17195 349
rect 16995 268 17195 315
rect 17253 349 17453 365
rect 17253 315 17302 349
rect 17336 315 17370 349
rect 17404 315 17453 349
rect 17253 268 17453 315
rect 17511 349 17711 365
rect 17511 315 17560 349
rect 17594 315 17628 349
rect 17662 315 17711 349
rect 17511 268 17711 315
rect 17963 349 18163 365
rect 17963 315 18012 349
rect 18046 315 18080 349
rect 18114 315 18163 349
rect 17963 268 18163 315
rect 9734 42 9934 68
rect 10186 42 10386 68
rect 10444 42 10644 68
rect 10702 42 10902 68
rect 10960 42 11160 68
rect 11412 42 11612 68
rect 11670 42 11870 68
rect 11928 42 12128 68
rect 12380 42 12580 68
rect 12638 42 12838 68
rect 12896 42 13096 68
rect 13154 42 13354 68
rect 13606 42 13806 68
rect 14092 42 14292 68
rect 14543 42 14743 68
rect 14801 42 15001 68
rect 15059 42 15259 68
rect 15317 42 15517 68
rect 15769 42 15969 68
rect 16027 42 16227 68
rect 16285 42 16485 68
rect 16737 42 16937 68
rect 16995 42 17195 68
rect 17253 42 17453 68
rect 17511 42 17711 68
rect 17963 42 18163 68
rect 1017 -676 1217 -650
rect 1469 -676 1669 -650
rect 1727 -676 1927 -650
rect 1985 -676 2185 -650
rect 2243 -676 2443 -650
rect 2695 -676 2895 -650
rect 2953 -676 3153 -650
rect 3211 -676 3411 -650
rect 3663 -676 3863 -650
rect 3921 -676 4121 -650
rect 4179 -676 4379 -650
rect 4437 -676 4637 -650
rect 4888 -676 5088 -650
rect 5374 -676 5574 -650
rect 5826 -676 6026 -650
rect 6084 -676 6284 -650
rect 6342 -676 6542 -650
rect 6600 -676 6800 -650
rect 7052 -676 7252 -650
rect 7310 -676 7510 -650
rect 7568 -676 7768 -650
rect 8020 -676 8220 -650
rect 8278 -676 8478 -650
rect 8536 -676 8736 -650
rect 8794 -676 8994 -650
rect 9246 -676 9446 -650
rect 1017 -923 1217 -876
rect 1017 -957 1066 -923
rect 1100 -957 1134 -923
rect 1168 -957 1217 -923
rect 1017 -973 1217 -957
rect 1469 -923 1669 -876
rect 1469 -957 1518 -923
rect 1552 -957 1586 -923
rect 1620 -957 1669 -923
rect 1469 -973 1669 -957
rect 1727 -923 1927 -876
rect 1727 -957 1776 -923
rect 1810 -957 1844 -923
rect 1878 -957 1927 -923
rect 1727 -973 1927 -957
rect 1985 -923 2185 -876
rect 1985 -957 2034 -923
rect 2068 -957 2102 -923
rect 2136 -957 2185 -923
rect 1985 -973 2185 -957
rect 2243 -923 2443 -876
rect 2243 -957 2292 -923
rect 2326 -957 2360 -923
rect 2394 -957 2443 -923
rect 2243 -973 2443 -957
rect 2695 -923 2895 -876
rect 2695 -957 2744 -923
rect 2778 -957 2812 -923
rect 2846 -957 2895 -923
rect 2695 -973 2895 -957
rect 2953 -923 3153 -876
rect 2953 -957 3002 -923
rect 3036 -957 3070 -923
rect 3104 -957 3153 -923
rect 2953 -973 3153 -957
rect 3211 -923 3411 -876
rect 3211 -957 3260 -923
rect 3294 -957 3328 -923
rect 3362 -957 3411 -923
rect 3211 -973 3411 -957
rect 3663 -923 3863 -876
rect 3663 -957 3712 -923
rect 3746 -957 3780 -923
rect 3814 -957 3863 -923
rect 3663 -973 3863 -957
rect 3921 -923 4121 -876
rect 3921 -957 3970 -923
rect 4004 -957 4038 -923
rect 4072 -957 4121 -923
rect 3921 -973 4121 -957
rect 4179 -923 4379 -876
rect 4179 -957 4228 -923
rect 4262 -957 4296 -923
rect 4330 -957 4379 -923
rect 4179 -973 4379 -957
rect 4437 -923 4637 -876
rect 4437 -957 4486 -923
rect 4520 -957 4554 -923
rect 4588 -957 4637 -923
rect 4437 -973 4637 -957
rect 4888 -923 5088 -876
rect 4888 -957 4937 -923
rect 4971 -957 5005 -923
rect 5039 -957 5088 -923
rect 4888 -973 5088 -957
rect 9734 -676 9934 -650
rect 10186 -676 10386 -650
rect 10444 -676 10644 -650
rect 10702 -676 10902 -650
rect 10960 -676 11160 -650
rect 11412 -676 11612 -650
rect 11670 -676 11870 -650
rect 11928 -676 12128 -650
rect 12380 -676 12580 -650
rect 12638 -676 12838 -650
rect 12896 -676 13096 -650
rect 13154 -676 13354 -650
rect 13606 -676 13806 -650
rect 5374 -923 5574 -876
rect 5374 -957 5423 -923
rect 5457 -957 5491 -923
rect 5525 -957 5574 -923
rect 5374 -973 5574 -957
rect 5826 -923 6026 -876
rect 5826 -957 5875 -923
rect 5909 -957 5943 -923
rect 5977 -957 6026 -923
rect 5826 -973 6026 -957
rect 6084 -923 6284 -876
rect 6084 -957 6133 -923
rect 6167 -957 6201 -923
rect 6235 -957 6284 -923
rect 6084 -973 6284 -957
rect 6342 -923 6542 -876
rect 6342 -957 6391 -923
rect 6425 -957 6459 -923
rect 6493 -957 6542 -923
rect 6342 -973 6542 -957
rect 6600 -923 6800 -876
rect 6600 -957 6649 -923
rect 6683 -957 6717 -923
rect 6751 -957 6800 -923
rect 6600 -973 6800 -957
rect 7052 -923 7252 -876
rect 7052 -957 7101 -923
rect 7135 -957 7169 -923
rect 7203 -957 7252 -923
rect 7052 -973 7252 -957
rect 7310 -923 7510 -876
rect 7310 -957 7359 -923
rect 7393 -957 7427 -923
rect 7461 -957 7510 -923
rect 7310 -973 7510 -957
rect 7568 -923 7768 -876
rect 7568 -957 7617 -923
rect 7651 -957 7685 -923
rect 7719 -957 7768 -923
rect 7568 -973 7768 -957
rect 8020 -923 8220 -876
rect 8020 -957 8069 -923
rect 8103 -957 8137 -923
rect 8171 -957 8220 -923
rect 8020 -973 8220 -957
rect 8278 -923 8478 -876
rect 8278 -957 8327 -923
rect 8361 -957 8395 -923
rect 8429 -957 8478 -923
rect 8278 -973 8478 -957
rect 8536 -923 8736 -876
rect 8536 -957 8585 -923
rect 8619 -957 8653 -923
rect 8687 -957 8736 -923
rect 8536 -973 8736 -957
rect 8794 -923 8994 -876
rect 8794 -957 8843 -923
rect 8877 -957 8911 -923
rect 8945 -957 8994 -923
rect 8794 -973 8994 -957
rect 9246 -923 9446 -876
rect 9246 -957 9295 -923
rect 9329 -957 9363 -923
rect 9397 -957 9446 -923
rect 9246 -973 9446 -957
rect 14092 -676 14292 -650
rect 14543 -676 14743 -650
rect 14801 -676 15001 -650
rect 15059 -676 15259 -650
rect 15317 -676 15517 -650
rect 15769 -676 15969 -650
rect 16027 -676 16227 -650
rect 16285 -676 16485 -650
rect 16737 -676 16937 -650
rect 16995 -676 17195 -650
rect 17253 -676 17453 -650
rect 17511 -676 17711 -650
rect 17963 -676 18163 -650
rect 1017 -1286 1217 -1270
rect 1017 -1320 1066 -1286
rect 1100 -1320 1134 -1286
rect 1168 -1320 1217 -1286
rect 1017 -1367 1217 -1320
rect 1469 -1286 1669 -1270
rect 1469 -1320 1518 -1286
rect 1552 -1320 1586 -1286
rect 1620 -1320 1669 -1286
rect 1469 -1367 1669 -1320
rect 1727 -1286 1927 -1270
rect 1727 -1320 1776 -1286
rect 1810 -1320 1844 -1286
rect 1878 -1320 1927 -1286
rect 1727 -1367 1927 -1320
rect 1985 -1286 2185 -1270
rect 1985 -1320 2034 -1286
rect 2068 -1320 2102 -1286
rect 2136 -1320 2185 -1286
rect 1985 -1367 2185 -1320
rect 2243 -1286 2443 -1270
rect 2243 -1320 2292 -1286
rect 2326 -1320 2360 -1286
rect 2394 -1320 2443 -1286
rect 2243 -1367 2443 -1320
rect 2695 -1286 2895 -1270
rect 2695 -1320 2744 -1286
rect 2778 -1320 2812 -1286
rect 2846 -1320 2895 -1286
rect 2695 -1367 2895 -1320
rect 2953 -1286 3153 -1270
rect 2953 -1320 3002 -1286
rect 3036 -1320 3070 -1286
rect 3104 -1320 3153 -1286
rect 2953 -1367 3153 -1320
rect 3211 -1286 3411 -1270
rect 3211 -1320 3260 -1286
rect 3294 -1320 3328 -1286
rect 3362 -1320 3411 -1286
rect 3211 -1367 3411 -1320
rect 3663 -1286 3863 -1270
rect 3663 -1320 3712 -1286
rect 3746 -1320 3780 -1286
rect 3814 -1320 3863 -1286
rect 3663 -1367 3863 -1320
rect 3921 -1286 4121 -1270
rect 3921 -1320 3970 -1286
rect 4004 -1320 4038 -1286
rect 4072 -1320 4121 -1286
rect 3921 -1367 4121 -1320
rect 4179 -1286 4379 -1270
rect 4179 -1320 4228 -1286
rect 4262 -1320 4296 -1286
rect 4330 -1320 4379 -1286
rect 4179 -1367 4379 -1320
rect 4437 -1286 4637 -1270
rect 4437 -1320 4486 -1286
rect 4520 -1320 4554 -1286
rect 4588 -1320 4637 -1286
rect 4437 -1367 4637 -1320
rect 4888 -1286 5088 -1270
rect 4888 -1320 4937 -1286
rect 4971 -1320 5005 -1286
rect 5039 -1320 5088 -1286
rect 4888 -1367 5088 -1320
rect 9734 -923 9934 -876
rect 9734 -957 9783 -923
rect 9817 -957 9851 -923
rect 9885 -957 9934 -923
rect 9734 -973 9934 -957
rect 10186 -923 10386 -876
rect 10186 -957 10235 -923
rect 10269 -957 10303 -923
rect 10337 -957 10386 -923
rect 10186 -973 10386 -957
rect 10444 -923 10644 -876
rect 10444 -957 10493 -923
rect 10527 -957 10561 -923
rect 10595 -957 10644 -923
rect 10444 -973 10644 -957
rect 10702 -923 10902 -876
rect 10702 -957 10751 -923
rect 10785 -957 10819 -923
rect 10853 -957 10902 -923
rect 10702 -973 10902 -957
rect 10960 -923 11160 -876
rect 10960 -957 11009 -923
rect 11043 -957 11077 -923
rect 11111 -957 11160 -923
rect 10960 -973 11160 -957
rect 11412 -923 11612 -876
rect 11412 -957 11461 -923
rect 11495 -957 11529 -923
rect 11563 -957 11612 -923
rect 11412 -973 11612 -957
rect 11670 -923 11870 -876
rect 11670 -957 11719 -923
rect 11753 -957 11787 -923
rect 11821 -957 11870 -923
rect 11670 -973 11870 -957
rect 11928 -923 12128 -876
rect 11928 -957 11977 -923
rect 12011 -957 12045 -923
rect 12079 -957 12128 -923
rect 11928 -973 12128 -957
rect 12380 -923 12580 -876
rect 12380 -957 12429 -923
rect 12463 -957 12497 -923
rect 12531 -957 12580 -923
rect 12380 -973 12580 -957
rect 12638 -923 12838 -876
rect 12638 -957 12687 -923
rect 12721 -957 12755 -923
rect 12789 -957 12838 -923
rect 12638 -973 12838 -957
rect 12896 -923 13096 -876
rect 12896 -957 12945 -923
rect 12979 -957 13013 -923
rect 13047 -957 13096 -923
rect 12896 -973 13096 -957
rect 13154 -923 13354 -876
rect 13154 -957 13203 -923
rect 13237 -957 13271 -923
rect 13305 -957 13354 -923
rect 13154 -973 13354 -957
rect 13606 -923 13806 -876
rect 13606 -957 13655 -923
rect 13689 -957 13723 -923
rect 13757 -957 13806 -923
rect 13606 -973 13806 -957
rect 5374 -1286 5574 -1270
rect 5374 -1320 5423 -1286
rect 5457 -1320 5491 -1286
rect 5525 -1320 5574 -1286
rect 5374 -1367 5574 -1320
rect 5826 -1286 6026 -1270
rect 5826 -1320 5875 -1286
rect 5909 -1320 5943 -1286
rect 5977 -1320 6026 -1286
rect 5826 -1367 6026 -1320
rect 6084 -1286 6284 -1270
rect 6084 -1320 6133 -1286
rect 6167 -1320 6201 -1286
rect 6235 -1320 6284 -1286
rect 6084 -1367 6284 -1320
rect 6342 -1286 6542 -1270
rect 6342 -1320 6391 -1286
rect 6425 -1320 6459 -1286
rect 6493 -1320 6542 -1286
rect 6342 -1367 6542 -1320
rect 6600 -1286 6800 -1270
rect 6600 -1320 6649 -1286
rect 6683 -1320 6717 -1286
rect 6751 -1320 6800 -1286
rect 6600 -1367 6800 -1320
rect 7052 -1286 7252 -1270
rect 7052 -1320 7101 -1286
rect 7135 -1320 7169 -1286
rect 7203 -1320 7252 -1286
rect 7052 -1367 7252 -1320
rect 7310 -1286 7510 -1270
rect 7310 -1320 7359 -1286
rect 7393 -1320 7427 -1286
rect 7461 -1320 7510 -1286
rect 7310 -1367 7510 -1320
rect 7568 -1286 7768 -1270
rect 7568 -1320 7617 -1286
rect 7651 -1320 7685 -1286
rect 7719 -1320 7768 -1286
rect 7568 -1367 7768 -1320
rect 8020 -1286 8220 -1270
rect 8020 -1320 8069 -1286
rect 8103 -1320 8137 -1286
rect 8171 -1320 8220 -1286
rect 8020 -1367 8220 -1320
rect 8278 -1286 8478 -1270
rect 8278 -1320 8327 -1286
rect 8361 -1320 8395 -1286
rect 8429 -1320 8478 -1286
rect 8278 -1367 8478 -1320
rect 8536 -1286 8736 -1270
rect 8536 -1320 8585 -1286
rect 8619 -1320 8653 -1286
rect 8687 -1320 8736 -1286
rect 8536 -1367 8736 -1320
rect 8794 -1286 8994 -1270
rect 8794 -1320 8843 -1286
rect 8877 -1320 8911 -1286
rect 8945 -1320 8994 -1286
rect 8794 -1367 8994 -1320
rect 9246 -1286 9446 -1270
rect 9246 -1320 9295 -1286
rect 9329 -1320 9363 -1286
rect 9397 -1320 9446 -1286
rect 9246 -1367 9446 -1320
rect 14092 -923 14292 -876
rect 14092 -957 14141 -923
rect 14175 -957 14209 -923
rect 14243 -957 14292 -923
rect 14092 -973 14292 -957
rect 14543 -923 14743 -876
rect 14543 -957 14592 -923
rect 14626 -957 14660 -923
rect 14694 -957 14743 -923
rect 14543 -973 14743 -957
rect 14801 -923 15001 -876
rect 14801 -957 14850 -923
rect 14884 -957 14918 -923
rect 14952 -957 15001 -923
rect 14801 -973 15001 -957
rect 15059 -923 15259 -876
rect 15059 -957 15108 -923
rect 15142 -957 15176 -923
rect 15210 -957 15259 -923
rect 15059 -973 15259 -957
rect 15317 -923 15517 -876
rect 15317 -957 15366 -923
rect 15400 -957 15434 -923
rect 15468 -957 15517 -923
rect 15317 -973 15517 -957
rect 15769 -923 15969 -876
rect 15769 -957 15818 -923
rect 15852 -957 15886 -923
rect 15920 -957 15969 -923
rect 15769 -973 15969 -957
rect 16027 -923 16227 -876
rect 16027 -957 16076 -923
rect 16110 -957 16144 -923
rect 16178 -957 16227 -923
rect 16027 -973 16227 -957
rect 16285 -923 16485 -876
rect 16285 -957 16334 -923
rect 16368 -957 16402 -923
rect 16436 -957 16485 -923
rect 16285 -973 16485 -957
rect 16737 -923 16937 -876
rect 16737 -957 16786 -923
rect 16820 -957 16854 -923
rect 16888 -957 16937 -923
rect 16737 -973 16937 -957
rect 16995 -923 17195 -876
rect 16995 -957 17044 -923
rect 17078 -957 17112 -923
rect 17146 -957 17195 -923
rect 16995 -973 17195 -957
rect 17253 -923 17453 -876
rect 17253 -957 17302 -923
rect 17336 -957 17370 -923
rect 17404 -957 17453 -923
rect 17253 -973 17453 -957
rect 17511 -923 17711 -876
rect 17511 -957 17560 -923
rect 17594 -957 17628 -923
rect 17662 -957 17711 -923
rect 17511 -973 17711 -957
rect 17963 -923 18163 -876
rect 17963 -957 18012 -923
rect 18046 -957 18080 -923
rect 18114 -957 18163 -923
rect 17963 -973 18163 -957
rect 1017 -1593 1217 -1567
rect 1469 -1593 1669 -1567
rect 1727 -1593 1927 -1567
rect 1985 -1593 2185 -1567
rect 2243 -1593 2443 -1567
rect 2695 -1593 2895 -1567
rect 2953 -1593 3153 -1567
rect 3211 -1593 3411 -1567
rect 3663 -1593 3863 -1567
rect 3921 -1593 4121 -1567
rect 4179 -1593 4379 -1567
rect 4437 -1593 4637 -1567
rect 4888 -1593 5088 -1567
rect 9734 -1286 9934 -1270
rect 9734 -1320 9783 -1286
rect 9817 -1320 9851 -1286
rect 9885 -1320 9934 -1286
rect 9734 -1367 9934 -1320
rect 10186 -1286 10386 -1270
rect 10186 -1320 10235 -1286
rect 10269 -1320 10303 -1286
rect 10337 -1320 10386 -1286
rect 10186 -1367 10386 -1320
rect 10444 -1286 10644 -1270
rect 10444 -1320 10493 -1286
rect 10527 -1320 10561 -1286
rect 10595 -1320 10644 -1286
rect 10444 -1367 10644 -1320
rect 10702 -1286 10902 -1270
rect 10702 -1320 10751 -1286
rect 10785 -1320 10819 -1286
rect 10853 -1320 10902 -1286
rect 10702 -1367 10902 -1320
rect 10960 -1286 11160 -1270
rect 10960 -1320 11009 -1286
rect 11043 -1320 11077 -1286
rect 11111 -1320 11160 -1286
rect 10960 -1367 11160 -1320
rect 11412 -1286 11612 -1270
rect 11412 -1320 11461 -1286
rect 11495 -1320 11529 -1286
rect 11563 -1320 11612 -1286
rect 11412 -1367 11612 -1320
rect 11670 -1286 11870 -1270
rect 11670 -1320 11719 -1286
rect 11753 -1320 11787 -1286
rect 11821 -1320 11870 -1286
rect 11670 -1367 11870 -1320
rect 11928 -1286 12128 -1270
rect 11928 -1320 11977 -1286
rect 12011 -1320 12045 -1286
rect 12079 -1320 12128 -1286
rect 11928 -1367 12128 -1320
rect 12380 -1286 12580 -1270
rect 12380 -1320 12429 -1286
rect 12463 -1320 12497 -1286
rect 12531 -1320 12580 -1286
rect 12380 -1367 12580 -1320
rect 12638 -1286 12838 -1270
rect 12638 -1320 12687 -1286
rect 12721 -1320 12755 -1286
rect 12789 -1320 12838 -1286
rect 12638 -1367 12838 -1320
rect 12896 -1286 13096 -1270
rect 12896 -1320 12945 -1286
rect 12979 -1320 13013 -1286
rect 13047 -1320 13096 -1286
rect 12896 -1367 13096 -1320
rect 13154 -1286 13354 -1270
rect 13154 -1320 13203 -1286
rect 13237 -1320 13271 -1286
rect 13305 -1320 13354 -1286
rect 13154 -1367 13354 -1320
rect 13606 -1286 13806 -1270
rect 13606 -1320 13655 -1286
rect 13689 -1320 13723 -1286
rect 13757 -1320 13806 -1286
rect 13606 -1367 13806 -1320
rect 5374 -1593 5574 -1567
rect 5826 -1593 6026 -1567
rect 6084 -1593 6284 -1567
rect 6342 -1593 6542 -1567
rect 6600 -1593 6800 -1567
rect 7052 -1593 7252 -1567
rect 7310 -1593 7510 -1567
rect 7568 -1593 7768 -1567
rect 8020 -1593 8220 -1567
rect 8278 -1593 8478 -1567
rect 8536 -1593 8736 -1567
rect 8794 -1593 8994 -1567
rect 9246 -1593 9446 -1567
rect 14092 -1286 14292 -1270
rect 14092 -1320 14141 -1286
rect 14175 -1320 14209 -1286
rect 14243 -1320 14292 -1286
rect 14092 -1367 14292 -1320
rect 14543 -1286 14743 -1270
rect 14543 -1320 14592 -1286
rect 14626 -1320 14660 -1286
rect 14694 -1320 14743 -1286
rect 14543 -1367 14743 -1320
rect 14801 -1286 15001 -1270
rect 14801 -1320 14850 -1286
rect 14884 -1320 14918 -1286
rect 14952 -1320 15001 -1286
rect 14801 -1367 15001 -1320
rect 15059 -1286 15259 -1270
rect 15059 -1320 15108 -1286
rect 15142 -1320 15176 -1286
rect 15210 -1320 15259 -1286
rect 15059 -1367 15259 -1320
rect 15317 -1286 15517 -1270
rect 15317 -1320 15366 -1286
rect 15400 -1320 15434 -1286
rect 15468 -1320 15517 -1286
rect 15317 -1367 15517 -1320
rect 15769 -1286 15969 -1270
rect 15769 -1320 15818 -1286
rect 15852 -1320 15886 -1286
rect 15920 -1320 15969 -1286
rect 15769 -1367 15969 -1320
rect 16027 -1286 16227 -1270
rect 16027 -1320 16076 -1286
rect 16110 -1320 16144 -1286
rect 16178 -1320 16227 -1286
rect 16027 -1367 16227 -1320
rect 16285 -1286 16485 -1270
rect 16285 -1320 16334 -1286
rect 16368 -1320 16402 -1286
rect 16436 -1320 16485 -1286
rect 16285 -1367 16485 -1320
rect 16737 -1286 16937 -1270
rect 16737 -1320 16786 -1286
rect 16820 -1320 16854 -1286
rect 16888 -1320 16937 -1286
rect 16737 -1367 16937 -1320
rect 16995 -1286 17195 -1270
rect 16995 -1320 17044 -1286
rect 17078 -1320 17112 -1286
rect 17146 -1320 17195 -1286
rect 16995 -1367 17195 -1320
rect 17253 -1286 17453 -1270
rect 17253 -1320 17302 -1286
rect 17336 -1320 17370 -1286
rect 17404 -1320 17453 -1286
rect 17253 -1367 17453 -1320
rect 17511 -1286 17711 -1270
rect 17511 -1320 17560 -1286
rect 17594 -1320 17628 -1286
rect 17662 -1320 17711 -1286
rect 17511 -1367 17711 -1320
rect 17963 -1286 18163 -1270
rect 17963 -1320 18012 -1286
rect 18046 -1320 18080 -1286
rect 18114 -1320 18163 -1286
rect 17963 -1367 18163 -1320
rect 9734 -1593 9934 -1567
rect 10186 -1593 10386 -1567
rect 10444 -1593 10644 -1567
rect 10702 -1593 10902 -1567
rect 10960 -1593 11160 -1567
rect 11412 -1593 11612 -1567
rect 11670 -1593 11870 -1567
rect 11928 -1593 12128 -1567
rect 12380 -1593 12580 -1567
rect 12638 -1593 12838 -1567
rect 12896 -1593 13096 -1567
rect 13154 -1593 13354 -1567
rect 13606 -1593 13806 -1567
rect 14092 -1593 14292 -1567
rect 14543 -1593 14743 -1567
rect 14801 -1593 15001 -1567
rect 15059 -1593 15259 -1567
rect 15317 -1593 15517 -1567
rect 15769 -1593 15969 -1567
rect 16027 -1593 16227 -1567
rect 16285 -1593 16485 -1567
rect 16737 -1593 16937 -1567
rect 16995 -1593 17195 -1567
rect 17253 -1593 17453 -1567
rect 17511 -1593 17711 -1567
rect 17963 -1593 18163 -1567
rect 1017 -2323 1217 -2297
rect 1469 -2323 1669 -2297
rect 1727 -2323 1927 -2297
rect 1985 -2323 2185 -2297
rect 2243 -2323 2443 -2297
rect 2695 -2323 2895 -2297
rect 2953 -2323 3153 -2297
rect 3211 -2323 3411 -2297
rect 3663 -2323 3863 -2297
rect 3921 -2323 4121 -2297
rect 4179 -2323 4379 -2297
rect 4437 -2323 4637 -2297
rect 4888 -2323 5088 -2297
rect 5374 -2323 5574 -2297
rect 5826 -2323 6026 -2297
rect 6084 -2323 6284 -2297
rect 6342 -2323 6542 -2297
rect 6600 -2323 6800 -2297
rect 7052 -2323 7252 -2297
rect 7310 -2323 7510 -2297
rect 7568 -2323 7768 -2297
rect 8020 -2323 8220 -2297
rect 8278 -2323 8478 -2297
rect 8536 -2323 8736 -2297
rect 8794 -2323 8994 -2297
rect 9246 -2323 9446 -2297
rect 1017 -2570 1217 -2523
rect 1017 -2604 1066 -2570
rect 1100 -2604 1134 -2570
rect 1168 -2604 1217 -2570
rect 1017 -2620 1217 -2604
rect 1469 -2570 1669 -2523
rect 1469 -2604 1518 -2570
rect 1552 -2604 1586 -2570
rect 1620 -2604 1669 -2570
rect 1469 -2620 1669 -2604
rect 1727 -2570 1927 -2523
rect 1727 -2604 1776 -2570
rect 1810 -2604 1844 -2570
rect 1878 -2604 1927 -2570
rect 1727 -2620 1927 -2604
rect 1985 -2570 2185 -2523
rect 1985 -2604 2034 -2570
rect 2068 -2604 2102 -2570
rect 2136 -2604 2185 -2570
rect 1985 -2620 2185 -2604
rect 2243 -2570 2443 -2523
rect 2243 -2604 2292 -2570
rect 2326 -2604 2360 -2570
rect 2394 -2604 2443 -2570
rect 2243 -2620 2443 -2604
rect 2695 -2570 2895 -2523
rect 2695 -2604 2744 -2570
rect 2778 -2604 2812 -2570
rect 2846 -2604 2895 -2570
rect 2695 -2620 2895 -2604
rect 2953 -2570 3153 -2523
rect 2953 -2604 3002 -2570
rect 3036 -2604 3070 -2570
rect 3104 -2604 3153 -2570
rect 2953 -2620 3153 -2604
rect 3211 -2570 3411 -2523
rect 3211 -2604 3260 -2570
rect 3294 -2604 3328 -2570
rect 3362 -2604 3411 -2570
rect 3211 -2620 3411 -2604
rect 3663 -2570 3863 -2523
rect 3663 -2604 3712 -2570
rect 3746 -2604 3780 -2570
rect 3814 -2604 3863 -2570
rect 3663 -2620 3863 -2604
rect 3921 -2570 4121 -2523
rect 3921 -2604 3970 -2570
rect 4004 -2604 4038 -2570
rect 4072 -2604 4121 -2570
rect 3921 -2620 4121 -2604
rect 4179 -2570 4379 -2523
rect 4179 -2604 4228 -2570
rect 4262 -2604 4296 -2570
rect 4330 -2604 4379 -2570
rect 4179 -2620 4379 -2604
rect 4437 -2570 4637 -2523
rect 4437 -2604 4486 -2570
rect 4520 -2604 4554 -2570
rect 4588 -2604 4637 -2570
rect 4437 -2620 4637 -2604
rect 4888 -2570 5088 -2523
rect 4888 -2604 4937 -2570
rect 4971 -2604 5005 -2570
rect 5039 -2604 5088 -2570
rect 4888 -2620 5088 -2604
rect 9734 -2323 9934 -2297
rect 10186 -2323 10386 -2297
rect 10444 -2323 10644 -2297
rect 10702 -2323 10902 -2297
rect 10960 -2323 11160 -2297
rect 11412 -2323 11612 -2297
rect 11670 -2323 11870 -2297
rect 11928 -2323 12128 -2297
rect 12380 -2323 12580 -2297
rect 12638 -2323 12838 -2297
rect 12896 -2323 13096 -2297
rect 13154 -2323 13354 -2297
rect 13606 -2323 13806 -2297
rect 5374 -2570 5574 -2523
rect 5374 -2604 5423 -2570
rect 5457 -2604 5491 -2570
rect 5525 -2604 5574 -2570
rect 5374 -2620 5574 -2604
rect 5826 -2570 6026 -2523
rect 5826 -2604 5875 -2570
rect 5909 -2604 5943 -2570
rect 5977 -2604 6026 -2570
rect 5826 -2620 6026 -2604
rect 6084 -2570 6284 -2523
rect 6084 -2604 6133 -2570
rect 6167 -2604 6201 -2570
rect 6235 -2604 6284 -2570
rect 6084 -2620 6284 -2604
rect 6342 -2570 6542 -2523
rect 6342 -2604 6391 -2570
rect 6425 -2604 6459 -2570
rect 6493 -2604 6542 -2570
rect 6342 -2620 6542 -2604
rect 6600 -2570 6800 -2523
rect 6600 -2604 6649 -2570
rect 6683 -2604 6717 -2570
rect 6751 -2604 6800 -2570
rect 6600 -2620 6800 -2604
rect 7052 -2570 7252 -2523
rect 7052 -2604 7101 -2570
rect 7135 -2604 7169 -2570
rect 7203 -2604 7252 -2570
rect 7052 -2620 7252 -2604
rect 7310 -2570 7510 -2523
rect 7310 -2604 7359 -2570
rect 7393 -2604 7427 -2570
rect 7461 -2604 7510 -2570
rect 7310 -2620 7510 -2604
rect 7568 -2570 7768 -2523
rect 7568 -2604 7617 -2570
rect 7651 -2604 7685 -2570
rect 7719 -2604 7768 -2570
rect 7568 -2620 7768 -2604
rect 8020 -2570 8220 -2523
rect 8020 -2604 8069 -2570
rect 8103 -2604 8137 -2570
rect 8171 -2604 8220 -2570
rect 8020 -2620 8220 -2604
rect 8278 -2570 8478 -2523
rect 8278 -2604 8327 -2570
rect 8361 -2604 8395 -2570
rect 8429 -2604 8478 -2570
rect 8278 -2620 8478 -2604
rect 8536 -2570 8736 -2523
rect 8536 -2604 8585 -2570
rect 8619 -2604 8653 -2570
rect 8687 -2604 8736 -2570
rect 8536 -2620 8736 -2604
rect 8794 -2570 8994 -2523
rect 8794 -2604 8843 -2570
rect 8877 -2604 8911 -2570
rect 8945 -2604 8994 -2570
rect 8794 -2620 8994 -2604
rect 9246 -2570 9446 -2523
rect 9246 -2604 9295 -2570
rect 9329 -2604 9363 -2570
rect 9397 -2604 9446 -2570
rect 9246 -2620 9446 -2604
rect 14092 -2323 14292 -2297
rect 14543 -2323 14743 -2297
rect 14801 -2323 15001 -2297
rect 15059 -2323 15259 -2297
rect 15317 -2323 15517 -2297
rect 15769 -2323 15969 -2297
rect 16027 -2323 16227 -2297
rect 16285 -2323 16485 -2297
rect 16737 -2323 16937 -2297
rect 16995 -2323 17195 -2297
rect 17253 -2323 17453 -2297
rect 17511 -2323 17711 -2297
rect 17963 -2323 18163 -2297
rect 1017 -2933 1217 -2917
rect 1017 -2967 1066 -2933
rect 1100 -2967 1134 -2933
rect 1168 -2967 1217 -2933
rect 1017 -3014 1217 -2967
rect 1469 -2933 1669 -2917
rect 1469 -2967 1518 -2933
rect 1552 -2967 1586 -2933
rect 1620 -2967 1669 -2933
rect 1469 -3014 1669 -2967
rect 1727 -2933 1927 -2917
rect 1727 -2967 1776 -2933
rect 1810 -2967 1844 -2933
rect 1878 -2967 1927 -2933
rect 1727 -3014 1927 -2967
rect 1985 -2933 2185 -2917
rect 1985 -2967 2034 -2933
rect 2068 -2967 2102 -2933
rect 2136 -2967 2185 -2933
rect 1985 -3014 2185 -2967
rect 2243 -2933 2443 -2917
rect 2243 -2967 2292 -2933
rect 2326 -2967 2360 -2933
rect 2394 -2967 2443 -2933
rect 2243 -3014 2443 -2967
rect 2695 -2933 2895 -2917
rect 2695 -2967 2744 -2933
rect 2778 -2967 2812 -2933
rect 2846 -2967 2895 -2933
rect 2695 -3014 2895 -2967
rect 2953 -2933 3153 -2917
rect 2953 -2967 3002 -2933
rect 3036 -2967 3070 -2933
rect 3104 -2967 3153 -2933
rect 2953 -3014 3153 -2967
rect 3211 -2933 3411 -2917
rect 3211 -2967 3260 -2933
rect 3294 -2967 3328 -2933
rect 3362 -2967 3411 -2933
rect 3211 -3014 3411 -2967
rect 3663 -2933 3863 -2917
rect 3663 -2967 3712 -2933
rect 3746 -2967 3780 -2933
rect 3814 -2967 3863 -2933
rect 3663 -3014 3863 -2967
rect 3921 -2933 4121 -2917
rect 3921 -2967 3970 -2933
rect 4004 -2967 4038 -2933
rect 4072 -2967 4121 -2933
rect 3921 -3014 4121 -2967
rect 4179 -2933 4379 -2917
rect 4179 -2967 4228 -2933
rect 4262 -2967 4296 -2933
rect 4330 -2967 4379 -2933
rect 4179 -3014 4379 -2967
rect 4437 -2933 4637 -2917
rect 4437 -2967 4486 -2933
rect 4520 -2967 4554 -2933
rect 4588 -2967 4637 -2933
rect 4437 -3014 4637 -2967
rect 4888 -2933 5088 -2917
rect 4888 -2967 4937 -2933
rect 4971 -2967 5005 -2933
rect 5039 -2967 5088 -2933
rect 4888 -3014 5088 -2967
rect 9734 -2570 9934 -2523
rect 9734 -2604 9783 -2570
rect 9817 -2604 9851 -2570
rect 9885 -2604 9934 -2570
rect 9734 -2620 9934 -2604
rect 10186 -2570 10386 -2523
rect 10186 -2604 10235 -2570
rect 10269 -2604 10303 -2570
rect 10337 -2604 10386 -2570
rect 10186 -2620 10386 -2604
rect 10444 -2570 10644 -2523
rect 10444 -2604 10493 -2570
rect 10527 -2604 10561 -2570
rect 10595 -2604 10644 -2570
rect 10444 -2620 10644 -2604
rect 10702 -2570 10902 -2523
rect 10702 -2604 10751 -2570
rect 10785 -2604 10819 -2570
rect 10853 -2604 10902 -2570
rect 10702 -2620 10902 -2604
rect 10960 -2570 11160 -2523
rect 10960 -2604 11009 -2570
rect 11043 -2604 11077 -2570
rect 11111 -2604 11160 -2570
rect 10960 -2620 11160 -2604
rect 11412 -2570 11612 -2523
rect 11412 -2604 11461 -2570
rect 11495 -2604 11529 -2570
rect 11563 -2604 11612 -2570
rect 11412 -2620 11612 -2604
rect 11670 -2570 11870 -2523
rect 11670 -2604 11719 -2570
rect 11753 -2604 11787 -2570
rect 11821 -2604 11870 -2570
rect 11670 -2620 11870 -2604
rect 11928 -2570 12128 -2523
rect 11928 -2604 11977 -2570
rect 12011 -2604 12045 -2570
rect 12079 -2604 12128 -2570
rect 11928 -2620 12128 -2604
rect 12380 -2570 12580 -2523
rect 12380 -2604 12429 -2570
rect 12463 -2604 12497 -2570
rect 12531 -2604 12580 -2570
rect 12380 -2620 12580 -2604
rect 12638 -2570 12838 -2523
rect 12638 -2604 12687 -2570
rect 12721 -2604 12755 -2570
rect 12789 -2604 12838 -2570
rect 12638 -2620 12838 -2604
rect 12896 -2570 13096 -2523
rect 12896 -2604 12945 -2570
rect 12979 -2604 13013 -2570
rect 13047 -2604 13096 -2570
rect 12896 -2620 13096 -2604
rect 13154 -2570 13354 -2523
rect 13154 -2604 13203 -2570
rect 13237 -2604 13271 -2570
rect 13305 -2604 13354 -2570
rect 13154 -2620 13354 -2604
rect 13606 -2570 13806 -2523
rect 13606 -2604 13655 -2570
rect 13689 -2604 13723 -2570
rect 13757 -2604 13806 -2570
rect 13606 -2620 13806 -2604
rect 5374 -2933 5574 -2917
rect 5374 -2967 5423 -2933
rect 5457 -2967 5491 -2933
rect 5525 -2967 5574 -2933
rect 5374 -3014 5574 -2967
rect 5826 -2933 6026 -2917
rect 5826 -2967 5875 -2933
rect 5909 -2967 5943 -2933
rect 5977 -2967 6026 -2933
rect 5826 -3014 6026 -2967
rect 6084 -2933 6284 -2917
rect 6084 -2967 6133 -2933
rect 6167 -2967 6201 -2933
rect 6235 -2967 6284 -2933
rect 6084 -3014 6284 -2967
rect 6342 -2933 6542 -2917
rect 6342 -2967 6391 -2933
rect 6425 -2967 6459 -2933
rect 6493 -2967 6542 -2933
rect 6342 -3014 6542 -2967
rect 6600 -2933 6800 -2917
rect 6600 -2967 6649 -2933
rect 6683 -2967 6717 -2933
rect 6751 -2967 6800 -2933
rect 6600 -3014 6800 -2967
rect 7052 -2933 7252 -2917
rect 7052 -2967 7101 -2933
rect 7135 -2967 7169 -2933
rect 7203 -2967 7252 -2933
rect 7052 -3014 7252 -2967
rect 7310 -2933 7510 -2917
rect 7310 -2967 7359 -2933
rect 7393 -2967 7427 -2933
rect 7461 -2967 7510 -2933
rect 7310 -3014 7510 -2967
rect 7568 -2933 7768 -2917
rect 7568 -2967 7617 -2933
rect 7651 -2967 7685 -2933
rect 7719 -2967 7768 -2933
rect 7568 -3014 7768 -2967
rect 8020 -2933 8220 -2917
rect 8020 -2967 8069 -2933
rect 8103 -2967 8137 -2933
rect 8171 -2967 8220 -2933
rect 8020 -3014 8220 -2967
rect 8278 -2933 8478 -2917
rect 8278 -2967 8327 -2933
rect 8361 -2967 8395 -2933
rect 8429 -2967 8478 -2933
rect 8278 -3014 8478 -2967
rect 8536 -2933 8736 -2917
rect 8536 -2967 8585 -2933
rect 8619 -2967 8653 -2933
rect 8687 -2967 8736 -2933
rect 8536 -3014 8736 -2967
rect 8794 -2933 8994 -2917
rect 8794 -2967 8843 -2933
rect 8877 -2967 8911 -2933
rect 8945 -2967 8994 -2933
rect 8794 -3014 8994 -2967
rect 9246 -2933 9446 -2917
rect 9246 -2967 9295 -2933
rect 9329 -2967 9363 -2933
rect 9397 -2967 9446 -2933
rect 9246 -3014 9446 -2967
rect 14092 -2570 14292 -2523
rect 14092 -2604 14141 -2570
rect 14175 -2604 14209 -2570
rect 14243 -2604 14292 -2570
rect 14092 -2620 14292 -2604
rect 14543 -2570 14743 -2523
rect 14543 -2604 14592 -2570
rect 14626 -2604 14660 -2570
rect 14694 -2604 14743 -2570
rect 14543 -2620 14743 -2604
rect 14801 -2570 15001 -2523
rect 14801 -2604 14850 -2570
rect 14884 -2604 14918 -2570
rect 14952 -2604 15001 -2570
rect 14801 -2620 15001 -2604
rect 15059 -2570 15259 -2523
rect 15059 -2604 15108 -2570
rect 15142 -2604 15176 -2570
rect 15210 -2604 15259 -2570
rect 15059 -2620 15259 -2604
rect 15317 -2570 15517 -2523
rect 15317 -2604 15366 -2570
rect 15400 -2604 15434 -2570
rect 15468 -2604 15517 -2570
rect 15317 -2620 15517 -2604
rect 15769 -2570 15969 -2523
rect 15769 -2604 15818 -2570
rect 15852 -2604 15886 -2570
rect 15920 -2604 15969 -2570
rect 15769 -2620 15969 -2604
rect 16027 -2570 16227 -2523
rect 16027 -2604 16076 -2570
rect 16110 -2604 16144 -2570
rect 16178 -2604 16227 -2570
rect 16027 -2620 16227 -2604
rect 16285 -2570 16485 -2523
rect 16285 -2604 16334 -2570
rect 16368 -2604 16402 -2570
rect 16436 -2604 16485 -2570
rect 16285 -2620 16485 -2604
rect 16737 -2570 16937 -2523
rect 16737 -2604 16786 -2570
rect 16820 -2604 16854 -2570
rect 16888 -2604 16937 -2570
rect 16737 -2620 16937 -2604
rect 16995 -2570 17195 -2523
rect 16995 -2604 17044 -2570
rect 17078 -2604 17112 -2570
rect 17146 -2604 17195 -2570
rect 16995 -2620 17195 -2604
rect 17253 -2570 17453 -2523
rect 17253 -2604 17302 -2570
rect 17336 -2604 17370 -2570
rect 17404 -2604 17453 -2570
rect 17253 -2620 17453 -2604
rect 17511 -2570 17711 -2523
rect 17511 -2604 17560 -2570
rect 17594 -2604 17628 -2570
rect 17662 -2604 17711 -2570
rect 17511 -2620 17711 -2604
rect 17963 -2570 18163 -2523
rect 17963 -2604 18012 -2570
rect 18046 -2604 18080 -2570
rect 18114 -2604 18163 -2570
rect 17963 -2620 18163 -2604
rect 9734 -2933 9934 -2917
rect 9734 -2967 9783 -2933
rect 9817 -2967 9851 -2933
rect 9885 -2967 9934 -2933
rect 9734 -3014 9934 -2967
rect 10186 -2933 10386 -2917
rect 10186 -2967 10235 -2933
rect 10269 -2967 10303 -2933
rect 10337 -2967 10386 -2933
rect 10186 -3014 10386 -2967
rect 10444 -2933 10644 -2917
rect 10444 -2967 10493 -2933
rect 10527 -2967 10561 -2933
rect 10595 -2967 10644 -2933
rect 10444 -3014 10644 -2967
rect 10702 -2933 10902 -2917
rect 10702 -2967 10751 -2933
rect 10785 -2967 10819 -2933
rect 10853 -2967 10902 -2933
rect 10702 -3014 10902 -2967
rect 10960 -2933 11160 -2917
rect 10960 -2967 11009 -2933
rect 11043 -2967 11077 -2933
rect 11111 -2967 11160 -2933
rect 10960 -3014 11160 -2967
rect 11412 -2933 11612 -2917
rect 11412 -2967 11461 -2933
rect 11495 -2967 11529 -2933
rect 11563 -2967 11612 -2933
rect 11412 -3014 11612 -2967
rect 11670 -2933 11870 -2917
rect 11670 -2967 11719 -2933
rect 11753 -2967 11787 -2933
rect 11821 -2967 11870 -2933
rect 11670 -3014 11870 -2967
rect 11928 -2933 12128 -2917
rect 11928 -2967 11977 -2933
rect 12011 -2967 12045 -2933
rect 12079 -2967 12128 -2933
rect 11928 -3014 12128 -2967
rect 12380 -2933 12580 -2917
rect 12380 -2967 12429 -2933
rect 12463 -2967 12497 -2933
rect 12531 -2967 12580 -2933
rect 12380 -3014 12580 -2967
rect 12638 -2933 12838 -2917
rect 12638 -2967 12687 -2933
rect 12721 -2967 12755 -2933
rect 12789 -2967 12838 -2933
rect 12638 -3014 12838 -2967
rect 12896 -2933 13096 -2917
rect 12896 -2967 12945 -2933
rect 12979 -2967 13013 -2933
rect 13047 -2967 13096 -2933
rect 12896 -3014 13096 -2967
rect 13154 -2933 13354 -2917
rect 13154 -2967 13203 -2933
rect 13237 -2967 13271 -2933
rect 13305 -2967 13354 -2933
rect 13154 -3014 13354 -2967
rect 13606 -2933 13806 -2917
rect 13606 -2967 13655 -2933
rect 13689 -2967 13723 -2933
rect 13757 -2967 13806 -2933
rect 13606 -3014 13806 -2967
rect 14092 -2933 14292 -2917
rect 14092 -2967 14141 -2933
rect 14175 -2967 14209 -2933
rect 14243 -2967 14292 -2933
rect 14092 -3014 14292 -2967
rect 14543 -2933 14743 -2917
rect 14543 -2967 14592 -2933
rect 14626 -2967 14660 -2933
rect 14694 -2967 14743 -2933
rect 14543 -3014 14743 -2967
rect 14801 -2933 15001 -2917
rect 14801 -2967 14850 -2933
rect 14884 -2967 14918 -2933
rect 14952 -2967 15001 -2933
rect 14801 -3014 15001 -2967
rect 15059 -2933 15259 -2917
rect 15059 -2967 15108 -2933
rect 15142 -2967 15176 -2933
rect 15210 -2967 15259 -2933
rect 15059 -3014 15259 -2967
rect 15317 -2933 15517 -2917
rect 15317 -2967 15366 -2933
rect 15400 -2967 15434 -2933
rect 15468 -2967 15517 -2933
rect 15317 -3014 15517 -2967
rect 15769 -2933 15969 -2917
rect 15769 -2967 15818 -2933
rect 15852 -2967 15886 -2933
rect 15920 -2967 15969 -2933
rect 15769 -3014 15969 -2967
rect 16027 -2933 16227 -2917
rect 16027 -2967 16076 -2933
rect 16110 -2967 16144 -2933
rect 16178 -2967 16227 -2933
rect 16027 -3014 16227 -2967
rect 16285 -2933 16485 -2917
rect 16285 -2967 16334 -2933
rect 16368 -2967 16402 -2933
rect 16436 -2967 16485 -2933
rect 16285 -3014 16485 -2967
rect 16737 -2933 16937 -2917
rect 16737 -2967 16786 -2933
rect 16820 -2967 16854 -2933
rect 16888 -2967 16937 -2933
rect 16737 -3014 16937 -2967
rect 16995 -2933 17195 -2917
rect 16995 -2967 17044 -2933
rect 17078 -2967 17112 -2933
rect 17146 -2967 17195 -2933
rect 16995 -3014 17195 -2967
rect 17253 -2933 17453 -2917
rect 17253 -2967 17302 -2933
rect 17336 -2967 17370 -2933
rect 17404 -2967 17453 -2933
rect 17253 -3014 17453 -2967
rect 17511 -2933 17711 -2917
rect 17511 -2967 17560 -2933
rect 17594 -2967 17628 -2933
rect 17662 -2967 17711 -2933
rect 17511 -3014 17711 -2967
rect 17963 -2933 18163 -2917
rect 17963 -2967 18012 -2933
rect 18046 -2967 18080 -2933
rect 18114 -2967 18163 -2933
rect 17963 -3014 18163 -2967
rect 1017 -3240 1217 -3214
rect 1469 -3240 1669 -3214
rect 1727 -3240 1927 -3214
rect 1985 -3240 2185 -3214
rect 2243 -3240 2443 -3214
rect 2695 -3240 2895 -3214
rect 2953 -3240 3153 -3214
rect 3211 -3240 3411 -3214
rect 3663 -3240 3863 -3214
rect 3921 -3240 4121 -3214
rect 4179 -3240 4379 -3214
rect 4437 -3240 4637 -3214
rect 4888 -3240 5088 -3214
rect 5374 -3240 5574 -3214
rect 5826 -3240 6026 -3214
rect 6084 -3240 6284 -3214
rect 6342 -3240 6542 -3214
rect 6600 -3240 6800 -3214
rect 7052 -3240 7252 -3214
rect 7310 -3240 7510 -3214
rect 7568 -3240 7768 -3214
rect 8020 -3240 8220 -3214
rect 8278 -3240 8478 -3214
rect 8536 -3240 8736 -3214
rect 8794 -3240 8994 -3214
rect 9246 -3240 9446 -3214
rect 9734 -3240 9934 -3214
rect 10186 -3240 10386 -3214
rect 10444 -3240 10644 -3214
rect 10702 -3240 10902 -3214
rect 10960 -3240 11160 -3214
rect 11412 -3240 11612 -3214
rect 11670 -3240 11870 -3214
rect 11928 -3240 12128 -3214
rect 12380 -3240 12580 -3214
rect 12638 -3240 12838 -3214
rect 12896 -3240 13096 -3214
rect 13154 -3240 13354 -3214
rect 13606 -3240 13806 -3214
rect 14092 -3240 14292 -3214
rect 14543 -3240 14743 -3214
rect 14801 -3240 15001 -3214
rect 15059 -3240 15259 -3214
rect 15317 -3240 15517 -3214
rect 15769 -3240 15969 -3214
rect 16027 -3240 16227 -3214
rect 16285 -3240 16485 -3214
rect 16737 -3240 16937 -3214
rect 16995 -3240 17195 -3214
rect 17253 -3240 17453 -3214
rect 17511 -3240 17711 -3214
rect 17963 -3240 18163 -3214
rect 1017 -4004 1217 -3978
rect 1469 -4004 1669 -3978
rect 1727 -4004 1927 -3978
rect 1985 -4004 2185 -3978
rect 2243 -4004 2443 -3978
rect 2695 -4004 2895 -3978
rect 2953 -4004 3153 -3978
rect 3211 -4004 3411 -3978
rect 3663 -4004 3863 -3978
rect 3921 -4004 4121 -3978
rect 4179 -4004 4379 -3978
rect 4437 -4004 4637 -3978
rect 4888 -4004 5088 -3978
rect 5374 -4004 5574 -3978
rect 5826 -4004 6026 -3978
rect 6084 -4004 6284 -3978
rect 6342 -4004 6542 -3978
rect 6600 -4004 6800 -3978
rect 7052 -4004 7252 -3978
rect 7310 -4004 7510 -3978
rect 7568 -4004 7768 -3978
rect 8020 -4004 8220 -3978
rect 8278 -4004 8478 -3978
rect 8536 -4004 8736 -3978
rect 8794 -4004 8994 -3978
rect 9246 -4004 9446 -3978
rect 1017 -4251 1217 -4204
rect 1017 -4285 1066 -4251
rect 1100 -4285 1134 -4251
rect 1168 -4285 1217 -4251
rect 1017 -4301 1217 -4285
rect 1469 -4251 1669 -4204
rect 1469 -4285 1518 -4251
rect 1552 -4285 1586 -4251
rect 1620 -4285 1669 -4251
rect 1469 -4301 1669 -4285
rect 1727 -4251 1927 -4204
rect 1727 -4285 1776 -4251
rect 1810 -4285 1844 -4251
rect 1878 -4285 1927 -4251
rect 1727 -4301 1927 -4285
rect 1985 -4251 2185 -4204
rect 1985 -4285 2034 -4251
rect 2068 -4285 2102 -4251
rect 2136 -4285 2185 -4251
rect 1985 -4301 2185 -4285
rect 2243 -4251 2443 -4204
rect 2243 -4285 2292 -4251
rect 2326 -4285 2360 -4251
rect 2394 -4285 2443 -4251
rect 2243 -4301 2443 -4285
rect 2695 -4251 2895 -4204
rect 2695 -4285 2744 -4251
rect 2778 -4285 2812 -4251
rect 2846 -4285 2895 -4251
rect 2695 -4301 2895 -4285
rect 2953 -4251 3153 -4204
rect 2953 -4285 3002 -4251
rect 3036 -4285 3070 -4251
rect 3104 -4285 3153 -4251
rect 2953 -4301 3153 -4285
rect 3211 -4251 3411 -4204
rect 3211 -4285 3260 -4251
rect 3294 -4285 3328 -4251
rect 3362 -4285 3411 -4251
rect 3211 -4301 3411 -4285
rect 3663 -4251 3863 -4204
rect 3663 -4285 3712 -4251
rect 3746 -4285 3780 -4251
rect 3814 -4285 3863 -4251
rect 3663 -4301 3863 -4285
rect 3921 -4251 4121 -4204
rect 3921 -4285 3970 -4251
rect 4004 -4285 4038 -4251
rect 4072 -4285 4121 -4251
rect 3921 -4301 4121 -4285
rect 4179 -4251 4379 -4204
rect 4179 -4285 4228 -4251
rect 4262 -4285 4296 -4251
rect 4330 -4285 4379 -4251
rect 4179 -4301 4379 -4285
rect 4437 -4251 4637 -4204
rect 4437 -4285 4486 -4251
rect 4520 -4285 4554 -4251
rect 4588 -4285 4637 -4251
rect 4437 -4301 4637 -4285
rect 4888 -4251 5088 -4204
rect 4888 -4285 4937 -4251
rect 4971 -4285 5005 -4251
rect 5039 -4285 5088 -4251
rect 4888 -4301 5088 -4285
rect 9734 -4004 9934 -3978
rect 10186 -4004 10386 -3978
rect 10444 -4004 10644 -3978
rect 10702 -4004 10902 -3978
rect 10960 -4004 11160 -3978
rect 11412 -4004 11612 -3978
rect 11670 -4004 11870 -3978
rect 11928 -4004 12128 -3978
rect 12380 -4004 12580 -3978
rect 12638 -4004 12838 -3978
rect 12896 -4004 13096 -3978
rect 13154 -4004 13354 -3978
rect 13606 -4004 13806 -3978
rect 5374 -4251 5574 -4204
rect 5374 -4285 5423 -4251
rect 5457 -4285 5491 -4251
rect 5525 -4285 5574 -4251
rect 5374 -4301 5574 -4285
rect 5826 -4251 6026 -4204
rect 5826 -4285 5875 -4251
rect 5909 -4285 5943 -4251
rect 5977 -4285 6026 -4251
rect 5826 -4301 6026 -4285
rect 6084 -4251 6284 -4204
rect 6084 -4285 6133 -4251
rect 6167 -4285 6201 -4251
rect 6235 -4285 6284 -4251
rect 6084 -4301 6284 -4285
rect 6342 -4251 6542 -4204
rect 6342 -4285 6391 -4251
rect 6425 -4285 6459 -4251
rect 6493 -4285 6542 -4251
rect 6342 -4301 6542 -4285
rect 6600 -4251 6800 -4204
rect 6600 -4285 6649 -4251
rect 6683 -4285 6717 -4251
rect 6751 -4285 6800 -4251
rect 6600 -4301 6800 -4285
rect 7052 -4251 7252 -4204
rect 7052 -4285 7101 -4251
rect 7135 -4285 7169 -4251
rect 7203 -4285 7252 -4251
rect 7052 -4301 7252 -4285
rect 7310 -4251 7510 -4204
rect 7310 -4285 7359 -4251
rect 7393 -4285 7427 -4251
rect 7461 -4285 7510 -4251
rect 7310 -4301 7510 -4285
rect 7568 -4251 7768 -4204
rect 7568 -4285 7617 -4251
rect 7651 -4285 7685 -4251
rect 7719 -4285 7768 -4251
rect 7568 -4301 7768 -4285
rect 8020 -4251 8220 -4204
rect 8020 -4285 8069 -4251
rect 8103 -4285 8137 -4251
rect 8171 -4285 8220 -4251
rect 8020 -4301 8220 -4285
rect 8278 -4251 8478 -4204
rect 8278 -4285 8327 -4251
rect 8361 -4285 8395 -4251
rect 8429 -4285 8478 -4251
rect 8278 -4301 8478 -4285
rect 8536 -4251 8736 -4204
rect 8536 -4285 8585 -4251
rect 8619 -4285 8653 -4251
rect 8687 -4285 8736 -4251
rect 8536 -4301 8736 -4285
rect 8794 -4251 8994 -4204
rect 8794 -4285 8843 -4251
rect 8877 -4285 8911 -4251
rect 8945 -4285 8994 -4251
rect 8794 -4301 8994 -4285
rect 9246 -4251 9446 -4204
rect 9246 -4285 9295 -4251
rect 9329 -4285 9363 -4251
rect 9397 -4285 9446 -4251
rect 9246 -4301 9446 -4285
rect 14092 -4004 14292 -3978
rect 14543 -4004 14743 -3978
rect 14801 -4004 15001 -3978
rect 15059 -4004 15259 -3978
rect 15317 -4004 15517 -3978
rect 15769 -4004 15969 -3978
rect 16027 -4004 16227 -3978
rect 16285 -4004 16485 -3978
rect 16737 -4004 16937 -3978
rect 16995 -4004 17195 -3978
rect 17253 -4004 17453 -3978
rect 17511 -4004 17711 -3978
rect 17963 -4004 18163 -3978
rect 9734 -4251 9934 -4204
rect 9734 -4285 9783 -4251
rect 9817 -4285 9851 -4251
rect 9885 -4285 9934 -4251
rect 9734 -4301 9934 -4285
rect 10186 -4251 10386 -4204
rect 10186 -4285 10235 -4251
rect 10269 -4285 10303 -4251
rect 10337 -4285 10386 -4251
rect 10186 -4301 10386 -4285
rect 10444 -4251 10644 -4204
rect 10444 -4285 10493 -4251
rect 10527 -4285 10561 -4251
rect 10595 -4285 10644 -4251
rect 10444 -4301 10644 -4285
rect 10702 -4251 10902 -4204
rect 10702 -4285 10751 -4251
rect 10785 -4285 10819 -4251
rect 10853 -4285 10902 -4251
rect 10702 -4301 10902 -4285
rect 10960 -4251 11160 -4204
rect 10960 -4285 11009 -4251
rect 11043 -4285 11077 -4251
rect 11111 -4285 11160 -4251
rect 10960 -4301 11160 -4285
rect 11412 -4251 11612 -4204
rect 11412 -4285 11461 -4251
rect 11495 -4285 11529 -4251
rect 11563 -4285 11612 -4251
rect 11412 -4301 11612 -4285
rect 11670 -4251 11870 -4204
rect 11670 -4285 11719 -4251
rect 11753 -4285 11787 -4251
rect 11821 -4285 11870 -4251
rect 11670 -4301 11870 -4285
rect 11928 -4251 12128 -4204
rect 11928 -4285 11977 -4251
rect 12011 -4285 12045 -4251
rect 12079 -4285 12128 -4251
rect 11928 -4301 12128 -4285
rect 12380 -4251 12580 -4204
rect 12380 -4285 12429 -4251
rect 12463 -4285 12497 -4251
rect 12531 -4285 12580 -4251
rect 12380 -4301 12580 -4285
rect 12638 -4251 12838 -4204
rect 12638 -4285 12687 -4251
rect 12721 -4285 12755 -4251
rect 12789 -4285 12838 -4251
rect 12638 -4301 12838 -4285
rect 12896 -4251 13096 -4204
rect 12896 -4285 12945 -4251
rect 12979 -4285 13013 -4251
rect 13047 -4285 13096 -4251
rect 12896 -4301 13096 -4285
rect 13154 -4251 13354 -4204
rect 13154 -4285 13203 -4251
rect 13237 -4285 13271 -4251
rect 13305 -4285 13354 -4251
rect 13154 -4301 13354 -4285
rect 13606 -4251 13806 -4204
rect 13606 -4285 13655 -4251
rect 13689 -4285 13723 -4251
rect 13757 -4285 13806 -4251
rect 13606 -4301 13806 -4285
rect 14092 -4251 14292 -4204
rect 14092 -4285 14141 -4251
rect 14175 -4285 14209 -4251
rect 14243 -4285 14292 -4251
rect 14092 -4301 14292 -4285
rect 14543 -4251 14743 -4204
rect 14543 -4285 14592 -4251
rect 14626 -4285 14660 -4251
rect 14694 -4285 14743 -4251
rect 14543 -4301 14743 -4285
rect 14801 -4251 15001 -4204
rect 14801 -4285 14850 -4251
rect 14884 -4285 14918 -4251
rect 14952 -4285 15001 -4251
rect 14801 -4301 15001 -4285
rect 15059 -4251 15259 -4204
rect 15059 -4285 15108 -4251
rect 15142 -4285 15176 -4251
rect 15210 -4285 15259 -4251
rect 15059 -4301 15259 -4285
rect 15317 -4251 15517 -4204
rect 15317 -4285 15366 -4251
rect 15400 -4285 15434 -4251
rect 15468 -4285 15517 -4251
rect 15317 -4301 15517 -4285
rect 15769 -4251 15969 -4204
rect 15769 -4285 15818 -4251
rect 15852 -4285 15886 -4251
rect 15920 -4285 15969 -4251
rect 15769 -4301 15969 -4285
rect 16027 -4251 16227 -4204
rect 16027 -4285 16076 -4251
rect 16110 -4285 16144 -4251
rect 16178 -4285 16227 -4251
rect 16027 -4301 16227 -4285
rect 16285 -4251 16485 -4204
rect 16285 -4285 16334 -4251
rect 16368 -4285 16402 -4251
rect 16436 -4285 16485 -4251
rect 16285 -4301 16485 -4285
rect 16737 -4251 16937 -4204
rect 16737 -4285 16786 -4251
rect 16820 -4285 16854 -4251
rect 16888 -4285 16937 -4251
rect 16737 -4301 16937 -4285
rect 16995 -4251 17195 -4204
rect 16995 -4285 17044 -4251
rect 17078 -4285 17112 -4251
rect 17146 -4285 17195 -4251
rect 16995 -4301 17195 -4285
rect 17253 -4251 17453 -4204
rect 17253 -4285 17302 -4251
rect 17336 -4285 17370 -4251
rect 17404 -4285 17453 -4251
rect 17253 -4301 17453 -4285
rect 17511 -4251 17711 -4204
rect 17511 -4285 17560 -4251
rect 17594 -4285 17628 -4251
rect 17662 -4285 17711 -4251
rect 17511 -4301 17711 -4285
rect 17963 -4251 18163 -4204
rect 17963 -4285 18012 -4251
rect 18046 -4285 18080 -4251
rect 18114 -4285 18163 -4251
rect 17963 -4301 18163 -4285
rect 1017 -4479 1217 -4463
rect 1017 -4513 1066 -4479
rect 1100 -4513 1134 -4479
rect 1168 -4513 1217 -4479
rect 1017 -4560 1217 -4513
rect 1469 -4479 1669 -4463
rect 1469 -4513 1518 -4479
rect 1552 -4513 1586 -4479
rect 1620 -4513 1669 -4479
rect 1469 -4560 1669 -4513
rect 1727 -4479 1927 -4463
rect 1727 -4513 1776 -4479
rect 1810 -4513 1844 -4479
rect 1878 -4513 1927 -4479
rect 1727 -4560 1927 -4513
rect 1985 -4479 2185 -4463
rect 1985 -4513 2034 -4479
rect 2068 -4513 2102 -4479
rect 2136 -4513 2185 -4479
rect 1985 -4560 2185 -4513
rect 2243 -4479 2443 -4463
rect 2243 -4513 2292 -4479
rect 2326 -4513 2360 -4479
rect 2394 -4513 2443 -4479
rect 2243 -4560 2443 -4513
rect 2695 -4479 2895 -4463
rect 2695 -4513 2744 -4479
rect 2778 -4513 2812 -4479
rect 2846 -4513 2895 -4479
rect 2695 -4560 2895 -4513
rect 2953 -4479 3153 -4463
rect 2953 -4513 3002 -4479
rect 3036 -4513 3070 -4479
rect 3104 -4513 3153 -4479
rect 2953 -4560 3153 -4513
rect 3211 -4479 3411 -4463
rect 3211 -4513 3260 -4479
rect 3294 -4513 3328 -4479
rect 3362 -4513 3411 -4479
rect 3211 -4560 3411 -4513
rect 3663 -4479 3863 -4463
rect 3663 -4513 3712 -4479
rect 3746 -4513 3780 -4479
rect 3814 -4513 3863 -4479
rect 3663 -4560 3863 -4513
rect 3921 -4479 4121 -4463
rect 3921 -4513 3970 -4479
rect 4004 -4513 4038 -4479
rect 4072 -4513 4121 -4479
rect 3921 -4560 4121 -4513
rect 4179 -4479 4379 -4463
rect 4179 -4513 4228 -4479
rect 4262 -4513 4296 -4479
rect 4330 -4513 4379 -4479
rect 4179 -4560 4379 -4513
rect 4437 -4479 4637 -4463
rect 4437 -4513 4486 -4479
rect 4520 -4513 4554 -4479
rect 4588 -4513 4637 -4479
rect 4437 -4560 4637 -4513
rect 4888 -4479 5088 -4463
rect 4888 -4513 4937 -4479
rect 4971 -4513 5005 -4479
rect 5039 -4513 5088 -4479
rect 4888 -4560 5088 -4513
rect 5374 -4479 5574 -4463
rect 5374 -4513 5423 -4479
rect 5457 -4513 5491 -4479
rect 5525 -4513 5574 -4479
rect 5374 -4560 5574 -4513
rect 5826 -4479 6026 -4463
rect 5826 -4513 5875 -4479
rect 5909 -4513 5943 -4479
rect 5977 -4513 6026 -4479
rect 5826 -4560 6026 -4513
rect 6084 -4479 6284 -4463
rect 6084 -4513 6133 -4479
rect 6167 -4513 6201 -4479
rect 6235 -4513 6284 -4479
rect 6084 -4560 6284 -4513
rect 6342 -4479 6542 -4463
rect 6342 -4513 6391 -4479
rect 6425 -4513 6459 -4479
rect 6493 -4513 6542 -4479
rect 6342 -4560 6542 -4513
rect 6600 -4479 6800 -4463
rect 6600 -4513 6649 -4479
rect 6683 -4513 6717 -4479
rect 6751 -4513 6800 -4479
rect 6600 -4560 6800 -4513
rect 7052 -4479 7252 -4463
rect 7052 -4513 7101 -4479
rect 7135 -4513 7169 -4479
rect 7203 -4513 7252 -4479
rect 7052 -4560 7252 -4513
rect 7310 -4479 7510 -4463
rect 7310 -4513 7359 -4479
rect 7393 -4513 7427 -4479
rect 7461 -4513 7510 -4479
rect 7310 -4560 7510 -4513
rect 7568 -4479 7768 -4463
rect 7568 -4513 7617 -4479
rect 7651 -4513 7685 -4479
rect 7719 -4513 7768 -4479
rect 7568 -4560 7768 -4513
rect 8020 -4479 8220 -4463
rect 8020 -4513 8069 -4479
rect 8103 -4513 8137 -4479
rect 8171 -4513 8220 -4479
rect 8020 -4560 8220 -4513
rect 8278 -4479 8478 -4463
rect 8278 -4513 8327 -4479
rect 8361 -4513 8395 -4479
rect 8429 -4513 8478 -4479
rect 8278 -4560 8478 -4513
rect 8536 -4479 8736 -4463
rect 8536 -4513 8585 -4479
rect 8619 -4513 8653 -4479
rect 8687 -4513 8736 -4479
rect 8536 -4560 8736 -4513
rect 8794 -4479 8994 -4463
rect 8794 -4513 8843 -4479
rect 8877 -4513 8911 -4479
rect 8945 -4513 8994 -4479
rect 8794 -4560 8994 -4513
rect 9246 -4479 9446 -4463
rect 9246 -4513 9295 -4479
rect 9329 -4513 9363 -4479
rect 9397 -4513 9446 -4479
rect 9246 -4560 9446 -4513
rect 1017 -4786 1217 -4760
rect 1469 -4786 1669 -4760
rect 1727 -4786 1927 -4760
rect 1985 -4786 2185 -4760
rect 2243 -4786 2443 -4760
rect 2695 -4786 2895 -4760
rect 2953 -4786 3153 -4760
rect 3211 -4786 3411 -4760
rect 3663 -4786 3863 -4760
rect 3921 -4786 4121 -4760
rect 4179 -4786 4379 -4760
rect 4437 -4786 4637 -4760
rect 4888 -4786 5088 -4760
rect 9734 -4479 9934 -4463
rect 9734 -4513 9783 -4479
rect 9817 -4513 9851 -4479
rect 9885 -4513 9934 -4479
rect 9734 -4560 9934 -4513
rect 10186 -4479 10386 -4463
rect 10186 -4513 10235 -4479
rect 10269 -4513 10303 -4479
rect 10337 -4513 10386 -4479
rect 10186 -4560 10386 -4513
rect 10444 -4479 10644 -4463
rect 10444 -4513 10493 -4479
rect 10527 -4513 10561 -4479
rect 10595 -4513 10644 -4479
rect 10444 -4560 10644 -4513
rect 10702 -4479 10902 -4463
rect 10702 -4513 10751 -4479
rect 10785 -4513 10819 -4479
rect 10853 -4513 10902 -4479
rect 10702 -4560 10902 -4513
rect 10960 -4479 11160 -4463
rect 10960 -4513 11009 -4479
rect 11043 -4513 11077 -4479
rect 11111 -4513 11160 -4479
rect 10960 -4560 11160 -4513
rect 11412 -4479 11612 -4463
rect 11412 -4513 11461 -4479
rect 11495 -4513 11529 -4479
rect 11563 -4513 11612 -4479
rect 11412 -4560 11612 -4513
rect 11670 -4479 11870 -4463
rect 11670 -4513 11719 -4479
rect 11753 -4513 11787 -4479
rect 11821 -4513 11870 -4479
rect 11670 -4560 11870 -4513
rect 11928 -4479 12128 -4463
rect 11928 -4513 11977 -4479
rect 12011 -4513 12045 -4479
rect 12079 -4513 12128 -4479
rect 11928 -4560 12128 -4513
rect 12380 -4479 12580 -4463
rect 12380 -4513 12429 -4479
rect 12463 -4513 12497 -4479
rect 12531 -4513 12580 -4479
rect 12380 -4560 12580 -4513
rect 12638 -4479 12838 -4463
rect 12638 -4513 12687 -4479
rect 12721 -4513 12755 -4479
rect 12789 -4513 12838 -4479
rect 12638 -4560 12838 -4513
rect 12896 -4479 13096 -4463
rect 12896 -4513 12945 -4479
rect 12979 -4513 13013 -4479
rect 13047 -4513 13096 -4479
rect 12896 -4560 13096 -4513
rect 13154 -4479 13354 -4463
rect 13154 -4513 13203 -4479
rect 13237 -4513 13271 -4479
rect 13305 -4513 13354 -4479
rect 13154 -4560 13354 -4513
rect 13606 -4479 13806 -4463
rect 13606 -4513 13655 -4479
rect 13689 -4513 13723 -4479
rect 13757 -4513 13806 -4479
rect 13606 -4560 13806 -4513
rect 5374 -4786 5574 -4760
rect 5826 -4786 6026 -4760
rect 6084 -4786 6284 -4760
rect 6342 -4786 6542 -4760
rect 6600 -4786 6800 -4760
rect 7052 -4786 7252 -4760
rect 7310 -4786 7510 -4760
rect 7568 -4786 7768 -4760
rect 8020 -4786 8220 -4760
rect 8278 -4786 8478 -4760
rect 8536 -4786 8736 -4760
rect 8794 -4786 8994 -4760
rect 9246 -4786 9446 -4760
rect 14092 -4479 14292 -4463
rect 14092 -4513 14141 -4479
rect 14175 -4513 14209 -4479
rect 14243 -4513 14292 -4479
rect 14092 -4560 14292 -4513
rect 14543 -4479 14743 -4463
rect 14543 -4513 14592 -4479
rect 14626 -4513 14660 -4479
rect 14694 -4513 14743 -4479
rect 14543 -4560 14743 -4513
rect 14801 -4479 15001 -4463
rect 14801 -4513 14850 -4479
rect 14884 -4513 14918 -4479
rect 14952 -4513 15001 -4479
rect 14801 -4560 15001 -4513
rect 15059 -4479 15259 -4463
rect 15059 -4513 15108 -4479
rect 15142 -4513 15176 -4479
rect 15210 -4513 15259 -4479
rect 15059 -4560 15259 -4513
rect 15317 -4479 15517 -4463
rect 15317 -4513 15366 -4479
rect 15400 -4513 15434 -4479
rect 15468 -4513 15517 -4479
rect 15317 -4560 15517 -4513
rect 15769 -4479 15969 -4463
rect 15769 -4513 15818 -4479
rect 15852 -4513 15886 -4479
rect 15920 -4513 15969 -4479
rect 15769 -4560 15969 -4513
rect 16027 -4479 16227 -4463
rect 16027 -4513 16076 -4479
rect 16110 -4513 16144 -4479
rect 16178 -4513 16227 -4479
rect 16027 -4560 16227 -4513
rect 16285 -4479 16485 -4463
rect 16285 -4513 16334 -4479
rect 16368 -4513 16402 -4479
rect 16436 -4513 16485 -4479
rect 16285 -4560 16485 -4513
rect 16737 -4479 16937 -4463
rect 16737 -4513 16786 -4479
rect 16820 -4513 16854 -4479
rect 16888 -4513 16937 -4479
rect 16737 -4560 16937 -4513
rect 16995 -4479 17195 -4463
rect 16995 -4513 17044 -4479
rect 17078 -4513 17112 -4479
rect 17146 -4513 17195 -4479
rect 16995 -4560 17195 -4513
rect 17253 -4479 17453 -4463
rect 17253 -4513 17302 -4479
rect 17336 -4513 17370 -4479
rect 17404 -4513 17453 -4479
rect 17253 -4560 17453 -4513
rect 17511 -4479 17711 -4463
rect 17511 -4513 17560 -4479
rect 17594 -4513 17628 -4479
rect 17662 -4513 17711 -4479
rect 17511 -4560 17711 -4513
rect 17963 -4479 18163 -4463
rect 17963 -4513 18012 -4479
rect 18046 -4513 18080 -4479
rect 18114 -4513 18163 -4479
rect 17963 -4560 18163 -4513
rect 9734 -4786 9934 -4760
rect 10186 -4786 10386 -4760
rect 10444 -4786 10644 -4760
rect 10702 -4786 10902 -4760
rect 10960 -4786 11160 -4760
rect 11412 -4786 11612 -4760
rect 11670 -4786 11870 -4760
rect 11928 -4786 12128 -4760
rect 12380 -4786 12580 -4760
rect 12638 -4786 12838 -4760
rect 12896 -4786 13096 -4760
rect 13154 -4786 13354 -4760
rect 13606 -4786 13806 -4760
rect 14092 -4786 14292 -4760
rect 14543 -4786 14743 -4760
rect 14801 -4786 15001 -4760
rect 15059 -4786 15259 -4760
rect 15317 -4786 15517 -4760
rect 15769 -4786 15969 -4760
rect 16027 -4786 16227 -4760
rect 16285 -4786 16485 -4760
rect 16737 -4786 16937 -4760
rect 16995 -4786 17195 -4760
rect 17253 -4786 17453 -4760
rect 17511 -4786 17711 -4760
rect 17963 -4786 18163 -4760
rect 1017 -5550 1217 -5524
rect 1469 -5550 1669 -5524
rect 1727 -5550 1927 -5524
rect 1985 -5550 2185 -5524
rect 2243 -5550 2443 -5524
rect 2695 -5550 2895 -5524
rect 2953 -5550 3153 -5524
rect 3211 -5550 3411 -5524
rect 3663 -5550 3863 -5524
rect 3921 -5550 4121 -5524
rect 4179 -5550 4379 -5524
rect 4437 -5550 4637 -5524
rect 4888 -5550 5088 -5524
rect 5374 -5550 5574 -5524
rect 5826 -5550 6026 -5524
rect 6084 -5550 6284 -5524
rect 6342 -5550 6542 -5524
rect 6600 -5550 6800 -5524
rect 7052 -5550 7252 -5524
rect 7310 -5550 7510 -5524
rect 7568 -5550 7768 -5524
rect 8020 -5550 8220 -5524
rect 8278 -5550 8478 -5524
rect 8536 -5550 8736 -5524
rect 8794 -5550 8994 -5524
rect 9246 -5550 9446 -5524
rect 9734 -5550 9934 -5524
rect 10186 -5550 10386 -5524
rect 10444 -5550 10644 -5524
rect 10702 -5550 10902 -5524
rect 10960 -5550 11160 -5524
rect 11412 -5550 11612 -5524
rect 11670 -5550 11870 -5524
rect 11928 -5550 12128 -5524
rect 12380 -5550 12580 -5524
rect 12638 -5550 12838 -5524
rect 12896 -5550 13096 -5524
rect 13154 -5550 13354 -5524
rect 13606 -5550 13806 -5524
rect 14092 -5550 14292 -5524
rect 14543 -5550 14743 -5524
rect 14801 -5550 15001 -5524
rect 15059 -5550 15259 -5524
rect 15317 -5550 15517 -5524
rect 15769 -5550 15969 -5524
rect 16027 -5550 16227 -5524
rect 16285 -5550 16485 -5524
rect 16737 -5550 16937 -5524
rect 16995 -5550 17195 -5524
rect 17253 -5550 17453 -5524
rect 17511 -5550 17711 -5524
rect 17963 -5550 18163 -5524
rect 1017 -5797 1217 -5750
rect 1017 -5831 1066 -5797
rect 1100 -5831 1134 -5797
rect 1168 -5831 1217 -5797
rect 1017 -5847 1217 -5831
rect 1469 -5797 1669 -5750
rect 1469 -5831 1518 -5797
rect 1552 -5831 1586 -5797
rect 1620 -5831 1669 -5797
rect 1469 -5847 1669 -5831
rect 1727 -5797 1927 -5750
rect 1727 -5831 1776 -5797
rect 1810 -5831 1844 -5797
rect 1878 -5831 1927 -5797
rect 1727 -5847 1927 -5831
rect 1985 -5797 2185 -5750
rect 1985 -5831 2034 -5797
rect 2068 -5831 2102 -5797
rect 2136 -5831 2185 -5797
rect 1985 -5847 2185 -5831
rect 2243 -5797 2443 -5750
rect 2243 -5831 2292 -5797
rect 2326 -5831 2360 -5797
rect 2394 -5831 2443 -5797
rect 2243 -5847 2443 -5831
rect 2695 -5797 2895 -5750
rect 2695 -5831 2744 -5797
rect 2778 -5831 2812 -5797
rect 2846 -5831 2895 -5797
rect 2695 -5847 2895 -5831
rect 2953 -5797 3153 -5750
rect 2953 -5831 3002 -5797
rect 3036 -5831 3070 -5797
rect 3104 -5831 3153 -5797
rect 2953 -5847 3153 -5831
rect 3211 -5797 3411 -5750
rect 3211 -5831 3260 -5797
rect 3294 -5831 3328 -5797
rect 3362 -5831 3411 -5797
rect 3211 -5847 3411 -5831
rect 3663 -5797 3863 -5750
rect 3663 -5831 3712 -5797
rect 3746 -5831 3780 -5797
rect 3814 -5831 3863 -5797
rect 3663 -5847 3863 -5831
rect 3921 -5797 4121 -5750
rect 3921 -5831 3970 -5797
rect 4004 -5831 4038 -5797
rect 4072 -5831 4121 -5797
rect 3921 -5847 4121 -5831
rect 4179 -5797 4379 -5750
rect 4179 -5831 4228 -5797
rect 4262 -5831 4296 -5797
rect 4330 -5831 4379 -5797
rect 4179 -5847 4379 -5831
rect 4437 -5797 4637 -5750
rect 4437 -5831 4486 -5797
rect 4520 -5831 4554 -5797
rect 4588 -5831 4637 -5797
rect 4437 -5847 4637 -5831
rect 4888 -5797 5088 -5750
rect 4888 -5831 4937 -5797
rect 4971 -5831 5005 -5797
rect 5039 -5831 5088 -5797
rect 4888 -5847 5088 -5831
rect 5374 -5797 5574 -5750
rect 5374 -5831 5423 -5797
rect 5457 -5831 5491 -5797
rect 5525 -5831 5574 -5797
rect 5374 -5847 5574 -5831
rect 5826 -5797 6026 -5750
rect 5826 -5831 5875 -5797
rect 5909 -5831 5943 -5797
rect 5977 -5831 6026 -5797
rect 5826 -5847 6026 -5831
rect 6084 -5797 6284 -5750
rect 6084 -5831 6133 -5797
rect 6167 -5831 6201 -5797
rect 6235 -5831 6284 -5797
rect 6084 -5847 6284 -5831
rect 6342 -5797 6542 -5750
rect 6342 -5831 6391 -5797
rect 6425 -5831 6459 -5797
rect 6493 -5831 6542 -5797
rect 6342 -5847 6542 -5831
rect 6600 -5797 6800 -5750
rect 6600 -5831 6649 -5797
rect 6683 -5831 6717 -5797
rect 6751 -5831 6800 -5797
rect 6600 -5847 6800 -5831
rect 7052 -5797 7252 -5750
rect 7052 -5831 7101 -5797
rect 7135 -5831 7169 -5797
rect 7203 -5831 7252 -5797
rect 7052 -5847 7252 -5831
rect 7310 -5797 7510 -5750
rect 7310 -5831 7359 -5797
rect 7393 -5831 7427 -5797
rect 7461 -5831 7510 -5797
rect 7310 -5847 7510 -5831
rect 7568 -5797 7768 -5750
rect 7568 -5831 7617 -5797
rect 7651 -5831 7685 -5797
rect 7719 -5831 7768 -5797
rect 7568 -5847 7768 -5831
rect 8020 -5797 8220 -5750
rect 8020 -5831 8069 -5797
rect 8103 -5831 8137 -5797
rect 8171 -5831 8220 -5797
rect 8020 -5847 8220 -5831
rect 8278 -5797 8478 -5750
rect 8278 -5831 8327 -5797
rect 8361 -5831 8395 -5797
rect 8429 -5831 8478 -5797
rect 8278 -5847 8478 -5831
rect 8536 -5797 8736 -5750
rect 8536 -5831 8585 -5797
rect 8619 -5831 8653 -5797
rect 8687 -5831 8736 -5797
rect 8536 -5847 8736 -5831
rect 8794 -5797 8994 -5750
rect 8794 -5831 8843 -5797
rect 8877 -5831 8911 -5797
rect 8945 -5831 8994 -5797
rect 8794 -5847 8994 -5831
rect 9246 -5797 9446 -5750
rect 9246 -5831 9295 -5797
rect 9329 -5831 9363 -5797
rect 9397 -5831 9446 -5797
rect 9246 -5847 9446 -5831
rect 1017 -6159 1217 -6143
rect 1017 -6193 1066 -6159
rect 1100 -6193 1134 -6159
rect 1168 -6193 1217 -6159
rect 1017 -6240 1217 -6193
rect 1469 -6159 1669 -6143
rect 1469 -6193 1518 -6159
rect 1552 -6193 1586 -6159
rect 1620 -6193 1669 -6159
rect 1469 -6240 1669 -6193
rect 1727 -6159 1927 -6143
rect 1727 -6193 1776 -6159
rect 1810 -6193 1844 -6159
rect 1878 -6193 1927 -6159
rect 1727 -6240 1927 -6193
rect 1985 -6159 2185 -6143
rect 1985 -6193 2034 -6159
rect 2068 -6193 2102 -6159
rect 2136 -6193 2185 -6159
rect 1985 -6240 2185 -6193
rect 2243 -6159 2443 -6143
rect 2243 -6193 2292 -6159
rect 2326 -6193 2360 -6159
rect 2394 -6193 2443 -6159
rect 2243 -6240 2443 -6193
rect 2695 -6159 2895 -6143
rect 2695 -6193 2744 -6159
rect 2778 -6193 2812 -6159
rect 2846 -6193 2895 -6159
rect 2695 -6240 2895 -6193
rect 2953 -6159 3153 -6143
rect 2953 -6193 3002 -6159
rect 3036 -6193 3070 -6159
rect 3104 -6193 3153 -6159
rect 2953 -6240 3153 -6193
rect 3211 -6159 3411 -6143
rect 3211 -6193 3260 -6159
rect 3294 -6193 3328 -6159
rect 3362 -6193 3411 -6159
rect 3211 -6240 3411 -6193
rect 3663 -6159 3863 -6143
rect 3663 -6193 3712 -6159
rect 3746 -6193 3780 -6159
rect 3814 -6193 3863 -6159
rect 3663 -6240 3863 -6193
rect 3921 -6159 4121 -6143
rect 3921 -6193 3970 -6159
rect 4004 -6193 4038 -6159
rect 4072 -6193 4121 -6159
rect 3921 -6240 4121 -6193
rect 4179 -6159 4379 -6143
rect 4179 -6193 4228 -6159
rect 4262 -6193 4296 -6159
rect 4330 -6193 4379 -6159
rect 4179 -6240 4379 -6193
rect 4437 -6159 4637 -6143
rect 4437 -6193 4486 -6159
rect 4520 -6193 4554 -6159
rect 4588 -6193 4637 -6159
rect 4437 -6240 4637 -6193
rect 4888 -6159 5088 -6143
rect 4888 -6193 4937 -6159
rect 4971 -6193 5005 -6159
rect 5039 -6193 5088 -6159
rect 4888 -6240 5088 -6193
rect 9734 -5797 9934 -5750
rect 9734 -5831 9783 -5797
rect 9817 -5831 9851 -5797
rect 9885 -5831 9934 -5797
rect 9734 -5847 9934 -5831
rect 10186 -5797 10386 -5750
rect 10186 -5831 10235 -5797
rect 10269 -5831 10303 -5797
rect 10337 -5831 10386 -5797
rect 10186 -5847 10386 -5831
rect 10444 -5797 10644 -5750
rect 10444 -5831 10493 -5797
rect 10527 -5831 10561 -5797
rect 10595 -5831 10644 -5797
rect 10444 -5847 10644 -5831
rect 10702 -5797 10902 -5750
rect 10702 -5831 10751 -5797
rect 10785 -5831 10819 -5797
rect 10853 -5831 10902 -5797
rect 10702 -5847 10902 -5831
rect 10960 -5797 11160 -5750
rect 10960 -5831 11009 -5797
rect 11043 -5831 11077 -5797
rect 11111 -5831 11160 -5797
rect 10960 -5847 11160 -5831
rect 11412 -5797 11612 -5750
rect 11412 -5831 11461 -5797
rect 11495 -5831 11529 -5797
rect 11563 -5831 11612 -5797
rect 11412 -5847 11612 -5831
rect 11670 -5797 11870 -5750
rect 11670 -5831 11719 -5797
rect 11753 -5831 11787 -5797
rect 11821 -5831 11870 -5797
rect 11670 -5847 11870 -5831
rect 11928 -5797 12128 -5750
rect 11928 -5831 11977 -5797
rect 12011 -5831 12045 -5797
rect 12079 -5831 12128 -5797
rect 11928 -5847 12128 -5831
rect 12380 -5797 12580 -5750
rect 12380 -5831 12429 -5797
rect 12463 -5831 12497 -5797
rect 12531 -5831 12580 -5797
rect 12380 -5847 12580 -5831
rect 12638 -5797 12838 -5750
rect 12638 -5831 12687 -5797
rect 12721 -5831 12755 -5797
rect 12789 -5831 12838 -5797
rect 12638 -5847 12838 -5831
rect 12896 -5797 13096 -5750
rect 12896 -5831 12945 -5797
rect 12979 -5831 13013 -5797
rect 13047 -5831 13096 -5797
rect 12896 -5847 13096 -5831
rect 13154 -5797 13354 -5750
rect 13154 -5831 13203 -5797
rect 13237 -5831 13271 -5797
rect 13305 -5831 13354 -5797
rect 13154 -5847 13354 -5831
rect 13606 -5797 13806 -5750
rect 13606 -5831 13655 -5797
rect 13689 -5831 13723 -5797
rect 13757 -5831 13806 -5797
rect 13606 -5847 13806 -5831
rect 5374 -6159 5574 -6143
rect 5374 -6193 5423 -6159
rect 5457 -6193 5491 -6159
rect 5525 -6193 5574 -6159
rect 5374 -6240 5574 -6193
rect 5826 -6159 6026 -6143
rect 5826 -6193 5875 -6159
rect 5909 -6193 5943 -6159
rect 5977 -6193 6026 -6159
rect 5826 -6240 6026 -6193
rect 6084 -6159 6284 -6143
rect 6084 -6193 6133 -6159
rect 6167 -6193 6201 -6159
rect 6235 -6193 6284 -6159
rect 6084 -6240 6284 -6193
rect 6342 -6159 6542 -6143
rect 6342 -6193 6391 -6159
rect 6425 -6193 6459 -6159
rect 6493 -6193 6542 -6159
rect 6342 -6240 6542 -6193
rect 6600 -6159 6800 -6143
rect 6600 -6193 6649 -6159
rect 6683 -6193 6717 -6159
rect 6751 -6193 6800 -6159
rect 6600 -6240 6800 -6193
rect 7052 -6159 7252 -6143
rect 7052 -6193 7101 -6159
rect 7135 -6193 7169 -6159
rect 7203 -6193 7252 -6159
rect 7052 -6240 7252 -6193
rect 7310 -6159 7510 -6143
rect 7310 -6193 7359 -6159
rect 7393 -6193 7427 -6159
rect 7461 -6193 7510 -6159
rect 7310 -6240 7510 -6193
rect 7568 -6159 7768 -6143
rect 7568 -6193 7617 -6159
rect 7651 -6193 7685 -6159
rect 7719 -6193 7768 -6159
rect 7568 -6240 7768 -6193
rect 8020 -6159 8220 -6143
rect 8020 -6193 8069 -6159
rect 8103 -6193 8137 -6159
rect 8171 -6193 8220 -6159
rect 8020 -6240 8220 -6193
rect 8278 -6159 8478 -6143
rect 8278 -6193 8327 -6159
rect 8361 -6193 8395 -6159
rect 8429 -6193 8478 -6159
rect 8278 -6240 8478 -6193
rect 8536 -6159 8736 -6143
rect 8536 -6193 8585 -6159
rect 8619 -6193 8653 -6159
rect 8687 -6193 8736 -6159
rect 8536 -6240 8736 -6193
rect 8794 -6159 8994 -6143
rect 8794 -6193 8843 -6159
rect 8877 -6193 8911 -6159
rect 8945 -6193 8994 -6159
rect 8794 -6240 8994 -6193
rect 9246 -6159 9446 -6143
rect 9246 -6193 9295 -6159
rect 9329 -6193 9363 -6159
rect 9397 -6193 9446 -6159
rect 9246 -6240 9446 -6193
rect 14092 -5797 14292 -5750
rect 14092 -5831 14141 -5797
rect 14175 -5831 14209 -5797
rect 14243 -5831 14292 -5797
rect 14092 -5847 14292 -5831
rect 14543 -5797 14743 -5750
rect 14543 -5831 14592 -5797
rect 14626 -5831 14660 -5797
rect 14694 -5831 14743 -5797
rect 14543 -5847 14743 -5831
rect 14801 -5797 15001 -5750
rect 14801 -5831 14850 -5797
rect 14884 -5831 14918 -5797
rect 14952 -5831 15001 -5797
rect 14801 -5847 15001 -5831
rect 15059 -5797 15259 -5750
rect 15059 -5831 15108 -5797
rect 15142 -5831 15176 -5797
rect 15210 -5831 15259 -5797
rect 15059 -5847 15259 -5831
rect 15317 -5797 15517 -5750
rect 15317 -5831 15366 -5797
rect 15400 -5831 15434 -5797
rect 15468 -5831 15517 -5797
rect 15317 -5847 15517 -5831
rect 15769 -5797 15969 -5750
rect 15769 -5831 15818 -5797
rect 15852 -5831 15886 -5797
rect 15920 -5831 15969 -5797
rect 15769 -5847 15969 -5831
rect 16027 -5797 16227 -5750
rect 16027 -5831 16076 -5797
rect 16110 -5831 16144 -5797
rect 16178 -5831 16227 -5797
rect 16027 -5847 16227 -5831
rect 16285 -5797 16485 -5750
rect 16285 -5831 16334 -5797
rect 16368 -5831 16402 -5797
rect 16436 -5831 16485 -5797
rect 16285 -5847 16485 -5831
rect 16737 -5797 16937 -5750
rect 16737 -5831 16786 -5797
rect 16820 -5831 16854 -5797
rect 16888 -5831 16937 -5797
rect 16737 -5847 16937 -5831
rect 16995 -5797 17195 -5750
rect 16995 -5831 17044 -5797
rect 17078 -5831 17112 -5797
rect 17146 -5831 17195 -5797
rect 16995 -5847 17195 -5831
rect 17253 -5797 17453 -5750
rect 17253 -5831 17302 -5797
rect 17336 -5831 17370 -5797
rect 17404 -5831 17453 -5797
rect 17253 -5847 17453 -5831
rect 17511 -5797 17711 -5750
rect 17511 -5831 17560 -5797
rect 17594 -5831 17628 -5797
rect 17662 -5831 17711 -5797
rect 17511 -5847 17711 -5831
rect 17963 -5797 18163 -5750
rect 17963 -5831 18012 -5797
rect 18046 -5831 18080 -5797
rect 18114 -5831 18163 -5797
rect 17963 -5847 18163 -5831
rect 1017 -6466 1217 -6440
rect 1469 -6466 1669 -6440
rect 1727 -6466 1927 -6440
rect 1985 -6466 2185 -6440
rect 2243 -6466 2443 -6440
rect 2695 -6466 2895 -6440
rect 2953 -6466 3153 -6440
rect 3211 -6466 3411 -6440
rect 3663 -6466 3863 -6440
rect 3921 -6466 4121 -6440
rect 4179 -6466 4379 -6440
rect 4437 -6466 4637 -6440
rect 4888 -6466 5088 -6440
rect 9734 -6159 9934 -6143
rect 9734 -6193 9783 -6159
rect 9817 -6193 9851 -6159
rect 9885 -6193 9934 -6159
rect 9734 -6240 9934 -6193
rect 10186 -6159 10386 -6143
rect 10186 -6193 10235 -6159
rect 10269 -6193 10303 -6159
rect 10337 -6193 10386 -6159
rect 10186 -6240 10386 -6193
rect 10444 -6159 10644 -6143
rect 10444 -6193 10493 -6159
rect 10527 -6193 10561 -6159
rect 10595 -6193 10644 -6159
rect 10444 -6240 10644 -6193
rect 10702 -6159 10902 -6143
rect 10702 -6193 10751 -6159
rect 10785 -6193 10819 -6159
rect 10853 -6193 10902 -6159
rect 10702 -6240 10902 -6193
rect 10960 -6159 11160 -6143
rect 10960 -6193 11009 -6159
rect 11043 -6193 11077 -6159
rect 11111 -6193 11160 -6159
rect 10960 -6240 11160 -6193
rect 11412 -6159 11612 -6143
rect 11412 -6193 11461 -6159
rect 11495 -6193 11529 -6159
rect 11563 -6193 11612 -6159
rect 11412 -6240 11612 -6193
rect 11670 -6159 11870 -6143
rect 11670 -6193 11719 -6159
rect 11753 -6193 11787 -6159
rect 11821 -6193 11870 -6159
rect 11670 -6240 11870 -6193
rect 11928 -6159 12128 -6143
rect 11928 -6193 11977 -6159
rect 12011 -6193 12045 -6159
rect 12079 -6193 12128 -6159
rect 11928 -6240 12128 -6193
rect 12380 -6159 12580 -6143
rect 12380 -6193 12429 -6159
rect 12463 -6193 12497 -6159
rect 12531 -6193 12580 -6159
rect 12380 -6240 12580 -6193
rect 12638 -6159 12838 -6143
rect 12638 -6193 12687 -6159
rect 12721 -6193 12755 -6159
rect 12789 -6193 12838 -6159
rect 12638 -6240 12838 -6193
rect 12896 -6159 13096 -6143
rect 12896 -6193 12945 -6159
rect 12979 -6193 13013 -6159
rect 13047 -6193 13096 -6159
rect 12896 -6240 13096 -6193
rect 13154 -6159 13354 -6143
rect 13154 -6193 13203 -6159
rect 13237 -6193 13271 -6159
rect 13305 -6193 13354 -6159
rect 13154 -6240 13354 -6193
rect 13606 -6159 13806 -6143
rect 13606 -6193 13655 -6159
rect 13689 -6193 13723 -6159
rect 13757 -6193 13806 -6159
rect 13606 -6240 13806 -6193
rect 5374 -6466 5574 -6440
rect 5826 -6466 6026 -6440
rect 6084 -6466 6284 -6440
rect 6342 -6466 6542 -6440
rect 6600 -6466 6800 -6440
rect 7052 -6466 7252 -6440
rect 7310 -6466 7510 -6440
rect 7568 -6466 7768 -6440
rect 8020 -6466 8220 -6440
rect 8278 -6466 8478 -6440
rect 8536 -6466 8736 -6440
rect 8794 -6466 8994 -6440
rect 9246 -6466 9446 -6440
rect 14092 -6159 14292 -6143
rect 14092 -6193 14141 -6159
rect 14175 -6193 14209 -6159
rect 14243 -6193 14292 -6159
rect 14092 -6240 14292 -6193
rect 14543 -6159 14743 -6143
rect 14543 -6193 14592 -6159
rect 14626 -6193 14660 -6159
rect 14694 -6193 14743 -6159
rect 14543 -6240 14743 -6193
rect 14801 -6159 15001 -6143
rect 14801 -6193 14850 -6159
rect 14884 -6193 14918 -6159
rect 14952 -6193 15001 -6159
rect 14801 -6240 15001 -6193
rect 15059 -6159 15259 -6143
rect 15059 -6193 15108 -6159
rect 15142 -6193 15176 -6159
rect 15210 -6193 15259 -6159
rect 15059 -6240 15259 -6193
rect 15317 -6159 15517 -6143
rect 15317 -6193 15366 -6159
rect 15400 -6193 15434 -6159
rect 15468 -6193 15517 -6159
rect 15317 -6240 15517 -6193
rect 15769 -6159 15969 -6143
rect 15769 -6193 15818 -6159
rect 15852 -6193 15886 -6159
rect 15920 -6193 15969 -6159
rect 15769 -6240 15969 -6193
rect 16027 -6159 16227 -6143
rect 16027 -6193 16076 -6159
rect 16110 -6193 16144 -6159
rect 16178 -6193 16227 -6159
rect 16027 -6240 16227 -6193
rect 16285 -6159 16485 -6143
rect 16285 -6193 16334 -6159
rect 16368 -6193 16402 -6159
rect 16436 -6193 16485 -6159
rect 16285 -6240 16485 -6193
rect 16737 -6159 16937 -6143
rect 16737 -6193 16786 -6159
rect 16820 -6193 16854 -6159
rect 16888 -6193 16937 -6159
rect 16737 -6240 16937 -6193
rect 16995 -6159 17195 -6143
rect 16995 -6193 17044 -6159
rect 17078 -6193 17112 -6159
rect 17146 -6193 17195 -6159
rect 16995 -6240 17195 -6193
rect 17253 -6159 17453 -6143
rect 17253 -6193 17302 -6159
rect 17336 -6193 17370 -6159
rect 17404 -6193 17453 -6159
rect 17253 -6240 17453 -6193
rect 17511 -6159 17711 -6143
rect 17511 -6193 17560 -6159
rect 17594 -6193 17628 -6159
rect 17662 -6193 17711 -6159
rect 17511 -6240 17711 -6193
rect 17963 -6159 18163 -6143
rect 17963 -6193 18012 -6159
rect 18046 -6193 18080 -6159
rect 18114 -6193 18163 -6159
rect 17963 -6240 18163 -6193
rect 9734 -6466 9934 -6440
rect 10186 -6466 10386 -6440
rect 10444 -6466 10644 -6440
rect 10702 -6466 10902 -6440
rect 10960 -6466 11160 -6440
rect 11412 -6466 11612 -6440
rect 11670 -6466 11870 -6440
rect 11928 -6466 12128 -6440
rect 12380 -6466 12580 -6440
rect 12638 -6466 12838 -6440
rect 12896 -6466 13096 -6440
rect 13154 -6466 13354 -6440
rect 13606 -6466 13806 -6440
rect 14092 -6466 14292 -6440
rect 14543 -6466 14743 -6440
rect 14801 -6466 15001 -6440
rect 15059 -6466 15259 -6440
rect 15317 -6466 15517 -6440
rect 15769 -6466 15969 -6440
rect 16027 -6466 16227 -6440
rect 16285 -6466 16485 -6440
rect 16737 -6466 16937 -6440
rect 16995 -6466 17195 -6440
rect 17253 -6466 17453 -6440
rect 17511 -6466 17711 -6440
rect 17963 -6466 18163 -6440
rect 1017 -7197 1217 -7171
rect 1469 -7197 1669 -7171
rect 1727 -7197 1927 -7171
rect 1985 -7197 2185 -7171
rect 2243 -7197 2443 -7171
rect 2695 -7197 2895 -7171
rect 2953 -7197 3153 -7171
rect 3211 -7197 3411 -7171
rect 3663 -7197 3863 -7171
rect 3921 -7197 4121 -7171
rect 4179 -7197 4379 -7171
rect 4437 -7197 4637 -7171
rect 4888 -7197 5088 -7171
rect 5374 -7197 5574 -7171
rect 5826 -7197 6026 -7171
rect 6084 -7197 6284 -7171
rect 6342 -7197 6542 -7171
rect 6600 -7197 6800 -7171
rect 7052 -7197 7252 -7171
rect 7310 -7197 7510 -7171
rect 7568 -7197 7768 -7171
rect 8020 -7197 8220 -7171
rect 8278 -7197 8478 -7171
rect 8536 -7197 8736 -7171
rect 8794 -7197 8994 -7171
rect 9246 -7197 9446 -7171
rect 1017 -7444 1217 -7397
rect 1017 -7478 1066 -7444
rect 1100 -7478 1134 -7444
rect 1168 -7478 1217 -7444
rect 1017 -7494 1217 -7478
rect 1469 -7444 1669 -7397
rect 1469 -7478 1518 -7444
rect 1552 -7478 1586 -7444
rect 1620 -7478 1669 -7444
rect 1469 -7494 1669 -7478
rect 1727 -7444 1927 -7397
rect 1727 -7478 1776 -7444
rect 1810 -7478 1844 -7444
rect 1878 -7478 1927 -7444
rect 1727 -7494 1927 -7478
rect 1985 -7444 2185 -7397
rect 1985 -7478 2034 -7444
rect 2068 -7478 2102 -7444
rect 2136 -7478 2185 -7444
rect 1985 -7494 2185 -7478
rect 2243 -7444 2443 -7397
rect 2243 -7478 2292 -7444
rect 2326 -7478 2360 -7444
rect 2394 -7478 2443 -7444
rect 2243 -7494 2443 -7478
rect 2695 -7444 2895 -7397
rect 2695 -7478 2744 -7444
rect 2778 -7478 2812 -7444
rect 2846 -7478 2895 -7444
rect 2695 -7494 2895 -7478
rect 2953 -7444 3153 -7397
rect 2953 -7478 3002 -7444
rect 3036 -7478 3070 -7444
rect 3104 -7478 3153 -7444
rect 2953 -7494 3153 -7478
rect 3211 -7444 3411 -7397
rect 3211 -7478 3260 -7444
rect 3294 -7478 3328 -7444
rect 3362 -7478 3411 -7444
rect 3211 -7494 3411 -7478
rect 3663 -7444 3863 -7397
rect 3663 -7478 3712 -7444
rect 3746 -7478 3780 -7444
rect 3814 -7478 3863 -7444
rect 3663 -7494 3863 -7478
rect 3921 -7444 4121 -7397
rect 3921 -7478 3970 -7444
rect 4004 -7478 4038 -7444
rect 4072 -7478 4121 -7444
rect 3921 -7494 4121 -7478
rect 4179 -7444 4379 -7397
rect 4179 -7478 4228 -7444
rect 4262 -7478 4296 -7444
rect 4330 -7478 4379 -7444
rect 4179 -7494 4379 -7478
rect 4437 -7444 4637 -7397
rect 4437 -7478 4486 -7444
rect 4520 -7478 4554 -7444
rect 4588 -7478 4637 -7444
rect 4437 -7494 4637 -7478
rect 4888 -7444 5088 -7397
rect 4888 -7478 4937 -7444
rect 4971 -7478 5005 -7444
rect 5039 -7478 5088 -7444
rect 4888 -7494 5088 -7478
rect 9734 -7197 9934 -7171
rect 10186 -7197 10386 -7171
rect 10444 -7197 10644 -7171
rect 10702 -7197 10902 -7171
rect 10960 -7197 11160 -7171
rect 11412 -7197 11612 -7171
rect 11670 -7197 11870 -7171
rect 11928 -7197 12128 -7171
rect 12380 -7197 12580 -7171
rect 12638 -7197 12838 -7171
rect 12896 -7197 13096 -7171
rect 13154 -7197 13354 -7171
rect 13606 -7197 13806 -7171
rect 5374 -7444 5574 -7397
rect 5374 -7478 5423 -7444
rect 5457 -7478 5491 -7444
rect 5525 -7478 5574 -7444
rect 5374 -7494 5574 -7478
rect 5826 -7444 6026 -7397
rect 5826 -7478 5875 -7444
rect 5909 -7478 5943 -7444
rect 5977 -7478 6026 -7444
rect 5826 -7494 6026 -7478
rect 6084 -7444 6284 -7397
rect 6084 -7478 6133 -7444
rect 6167 -7478 6201 -7444
rect 6235 -7478 6284 -7444
rect 6084 -7494 6284 -7478
rect 6342 -7444 6542 -7397
rect 6342 -7478 6391 -7444
rect 6425 -7478 6459 -7444
rect 6493 -7478 6542 -7444
rect 6342 -7494 6542 -7478
rect 6600 -7444 6800 -7397
rect 6600 -7478 6649 -7444
rect 6683 -7478 6717 -7444
rect 6751 -7478 6800 -7444
rect 6600 -7494 6800 -7478
rect 7052 -7444 7252 -7397
rect 7052 -7478 7101 -7444
rect 7135 -7478 7169 -7444
rect 7203 -7478 7252 -7444
rect 7052 -7494 7252 -7478
rect 7310 -7444 7510 -7397
rect 7310 -7478 7359 -7444
rect 7393 -7478 7427 -7444
rect 7461 -7478 7510 -7444
rect 7310 -7494 7510 -7478
rect 7568 -7444 7768 -7397
rect 7568 -7478 7617 -7444
rect 7651 -7478 7685 -7444
rect 7719 -7478 7768 -7444
rect 7568 -7494 7768 -7478
rect 8020 -7444 8220 -7397
rect 8020 -7478 8069 -7444
rect 8103 -7478 8137 -7444
rect 8171 -7478 8220 -7444
rect 8020 -7494 8220 -7478
rect 8278 -7444 8478 -7397
rect 8278 -7478 8327 -7444
rect 8361 -7478 8395 -7444
rect 8429 -7478 8478 -7444
rect 8278 -7494 8478 -7478
rect 8536 -7444 8736 -7397
rect 8536 -7478 8585 -7444
rect 8619 -7478 8653 -7444
rect 8687 -7478 8736 -7444
rect 8536 -7494 8736 -7478
rect 8794 -7444 8994 -7397
rect 8794 -7478 8843 -7444
rect 8877 -7478 8911 -7444
rect 8945 -7478 8994 -7444
rect 8794 -7494 8994 -7478
rect 9246 -7444 9446 -7397
rect 9246 -7478 9295 -7444
rect 9329 -7478 9363 -7444
rect 9397 -7478 9446 -7444
rect 9246 -7494 9446 -7478
rect 14092 -7197 14292 -7171
rect 14543 -7197 14743 -7171
rect 14801 -7197 15001 -7171
rect 15059 -7197 15259 -7171
rect 15317 -7197 15517 -7171
rect 15769 -7197 15969 -7171
rect 16027 -7197 16227 -7171
rect 16285 -7197 16485 -7171
rect 16737 -7197 16937 -7171
rect 16995 -7197 17195 -7171
rect 17253 -7197 17453 -7171
rect 17511 -7197 17711 -7171
rect 17963 -7197 18163 -7171
rect 9734 -7444 9934 -7397
rect 9734 -7478 9783 -7444
rect 9817 -7478 9851 -7444
rect 9885 -7478 9934 -7444
rect 9734 -7494 9934 -7478
rect 10186 -7444 10386 -7397
rect 10186 -7478 10235 -7444
rect 10269 -7478 10303 -7444
rect 10337 -7478 10386 -7444
rect 10186 -7494 10386 -7478
rect 10444 -7444 10644 -7397
rect 10444 -7478 10493 -7444
rect 10527 -7478 10561 -7444
rect 10595 -7478 10644 -7444
rect 10444 -7494 10644 -7478
rect 10702 -7444 10902 -7397
rect 10702 -7478 10751 -7444
rect 10785 -7478 10819 -7444
rect 10853 -7478 10902 -7444
rect 10702 -7494 10902 -7478
rect 10960 -7444 11160 -7397
rect 10960 -7478 11009 -7444
rect 11043 -7478 11077 -7444
rect 11111 -7478 11160 -7444
rect 10960 -7494 11160 -7478
rect 11412 -7444 11612 -7397
rect 11412 -7478 11461 -7444
rect 11495 -7478 11529 -7444
rect 11563 -7478 11612 -7444
rect 11412 -7494 11612 -7478
rect 11670 -7444 11870 -7397
rect 11670 -7478 11719 -7444
rect 11753 -7478 11787 -7444
rect 11821 -7478 11870 -7444
rect 11670 -7494 11870 -7478
rect 11928 -7444 12128 -7397
rect 11928 -7478 11977 -7444
rect 12011 -7478 12045 -7444
rect 12079 -7478 12128 -7444
rect 11928 -7494 12128 -7478
rect 12380 -7444 12580 -7397
rect 12380 -7478 12429 -7444
rect 12463 -7478 12497 -7444
rect 12531 -7478 12580 -7444
rect 12380 -7494 12580 -7478
rect 12638 -7444 12838 -7397
rect 12638 -7478 12687 -7444
rect 12721 -7478 12755 -7444
rect 12789 -7478 12838 -7444
rect 12638 -7494 12838 -7478
rect 12896 -7444 13096 -7397
rect 12896 -7478 12945 -7444
rect 12979 -7478 13013 -7444
rect 13047 -7478 13096 -7444
rect 12896 -7494 13096 -7478
rect 13154 -7444 13354 -7397
rect 13154 -7478 13203 -7444
rect 13237 -7478 13271 -7444
rect 13305 -7478 13354 -7444
rect 13154 -7494 13354 -7478
rect 13606 -7444 13806 -7397
rect 13606 -7478 13655 -7444
rect 13689 -7478 13723 -7444
rect 13757 -7478 13806 -7444
rect 13606 -7494 13806 -7478
rect 14092 -7444 14292 -7397
rect 14092 -7478 14141 -7444
rect 14175 -7478 14209 -7444
rect 14243 -7478 14292 -7444
rect 14092 -7494 14292 -7478
rect 14543 -7444 14743 -7397
rect 14543 -7478 14592 -7444
rect 14626 -7478 14660 -7444
rect 14694 -7478 14743 -7444
rect 14543 -7494 14743 -7478
rect 14801 -7444 15001 -7397
rect 14801 -7478 14850 -7444
rect 14884 -7478 14918 -7444
rect 14952 -7478 15001 -7444
rect 14801 -7494 15001 -7478
rect 15059 -7444 15259 -7397
rect 15059 -7478 15108 -7444
rect 15142 -7478 15176 -7444
rect 15210 -7478 15259 -7444
rect 15059 -7494 15259 -7478
rect 15317 -7444 15517 -7397
rect 15317 -7478 15366 -7444
rect 15400 -7478 15434 -7444
rect 15468 -7478 15517 -7444
rect 15317 -7494 15517 -7478
rect 15769 -7444 15969 -7397
rect 15769 -7478 15818 -7444
rect 15852 -7478 15886 -7444
rect 15920 -7478 15969 -7444
rect 15769 -7494 15969 -7478
rect 16027 -7444 16227 -7397
rect 16027 -7478 16076 -7444
rect 16110 -7478 16144 -7444
rect 16178 -7478 16227 -7444
rect 16027 -7494 16227 -7478
rect 16285 -7444 16485 -7397
rect 16285 -7478 16334 -7444
rect 16368 -7478 16402 -7444
rect 16436 -7478 16485 -7444
rect 16285 -7494 16485 -7478
rect 16737 -7444 16937 -7397
rect 16737 -7478 16786 -7444
rect 16820 -7478 16854 -7444
rect 16888 -7478 16937 -7444
rect 16737 -7494 16937 -7478
rect 16995 -7444 17195 -7397
rect 16995 -7478 17044 -7444
rect 17078 -7478 17112 -7444
rect 17146 -7478 17195 -7444
rect 16995 -7494 17195 -7478
rect 17253 -7444 17453 -7397
rect 17253 -7478 17302 -7444
rect 17336 -7478 17370 -7444
rect 17404 -7478 17453 -7444
rect 17253 -7494 17453 -7478
rect 17511 -7444 17711 -7397
rect 17511 -7478 17560 -7444
rect 17594 -7478 17628 -7444
rect 17662 -7478 17711 -7444
rect 17511 -7494 17711 -7478
rect 17963 -7444 18163 -7397
rect 17963 -7478 18012 -7444
rect 18046 -7478 18080 -7444
rect 18114 -7478 18163 -7444
rect 17963 -7494 18163 -7478
rect 1017 -7806 1217 -7790
rect 1017 -7840 1066 -7806
rect 1100 -7840 1134 -7806
rect 1168 -7840 1217 -7806
rect 1017 -7887 1217 -7840
rect 1469 -7806 1669 -7790
rect 1469 -7840 1518 -7806
rect 1552 -7840 1586 -7806
rect 1620 -7840 1669 -7806
rect 1469 -7887 1669 -7840
rect 1727 -7806 1927 -7790
rect 1727 -7840 1776 -7806
rect 1810 -7840 1844 -7806
rect 1878 -7840 1927 -7806
rect 1727 -7887 1927 -7840
rect 1985 -7806 2185 -7790
rect 1985 -7840 2034 -7806
rect 2068 -7840 2102 -7806
rect 2136 -7840 2185 -7806
rect 1985 -7887 2185 -7840
rect 2243 -7806 2443 -7790
rect 2243 -7840 2292 -7806
rect 2326 -7840 2360 -7806
rect 2394 -7840 2443 -7806
rect 2243 -7887 2443 -7840
rect 2695 -7806 2895 -7790
rect 2695 -7840 2744 -7806
rect 2778 -7840 2812 -7806
rect 2846 -7840 2895 -7806
rect 2695 -7887 2895 -7840
rect 2953 -7806 3153 -7790
rect 2953 -7840 3002 -7806
rect 3036 -7840 3070 -7806
rect 3104 -7840 3153 -7806
rect 2953 -7887 3153 -7840
rect 3211 -7806 3411 -7790
rect 3211 -7840 3260 -7806
rect 3294 -7840 3328 -7806
rect 3362 -7840 3411 -7806
rect 3211 -7887 3411 -7840
rect 3663 -7806 3863 -7790
rect 3663 -7840 3712 -7806
rect 3746 -7840 3780 -7806
rect 3814 -7840 3863 -7806
rect 3663 -7887 3863 -7840
rect 3921 -7806 4121 -7790
rect 3921 -7840 3970 -7806
rect 4004 -7840 4038 -7806
rect 4072 -7840 4121 -7806
rect 3921 -7887 4121 -7840
rect 4179 -7806 4379 -7790
rect 4179 -7840 4228 -7806
rect 4262 -7840 4296 -7806
rect 4330 -7840 4379 -7806
rect 4179 -7887 4379 -7840
rect 4437 -7806 4637 -7790
rect 4437 -7840 4486 -7806
rect 4520 -7840 4554 -7806
rect 4588 -7840 4637 -7806
rect 4437 -7887 4637 -7840
rect 4888 -7806 5088 -7790
rect 4888 -7840 4937 -7806
rect 4971 -7840 5005 -7806
rect 5039 -7840 5088 -7806
rect 4888 -7887 5088 -7840
rect 5374 -7806 5574 -7790
rect 5374 -7840 5423 -7806
rect 5457 -7840 5491 -7806
rect 5525 -7840 5574 -7806
rect 5374 -7887 5574 -7840
rect 5826 -7806 6026 -7790
rect 5826 -7840 5875 -7806
rect 5909 -7840 5943 -7806
rect 5977 -7840 6026 -7806
rect 5826 -7887 6026 -7840
rect 6084 -7806 6284 -7790
rect 6084 -7840 6133 -7806
rect 6167 -7840 6201 -7806
rect 6235 -7840 6284 -7806
rect 6084 -7887 6284 -7840
rect 6342 -7806 6542 -7790
rect 6342 -7840 6391 -7806
rect 6425 -7840 6459 -7806
rect 6493 -7840 6542 -7806
rect 6342 -7887 6542 -7840
rect 6600 -7806 6800 -7790
rect 6600 -7840 6649 -7806
rect 6683 -7840 6717 -7806
rect 6751 -7840 6800 -7806
rect 6600 -7887 6800 -7840
rect 7052 -7806 7252 -7790
rect 7052 -7840 7101 -7806
rect 7135 -7840 7169 -7806
rect 7203 -7840 7252 -7806
rect 7052 -7887 7252 -7840
rect 7310 -7806 7510 -7790
rect 7310 -7840 7359 -7806
rect 7393 -7840 7427 -7806
rect 7461 -7840 7510 -7806
rect 7310 -7887 7510 -7840
rect 7568 -7806 7768 -7790
rect 7568 -7840 7617 -7806
rect 7651 -7840 7685 -7806
rect 7719 -7840 7768 -7806
rect 7568 -7887 7768 -7840
rect 8020 -7806 8220 -7790
rect 8020 -7840 8069 -7806
rect 8103 -7840 8137 -7806
rect 8171 -7840 8220 -7806
rect 8020 -7887 8220 -7840
rect 8278 -7806 8478 -7790
rect 8278 -7840 8327 -7806
rect 8361 -7840 8395 -7806
rect 8429 -7840 8478 -7806
rect 8278 -7887 8478 -7840
rect 8536 -7806 8736 -7790
rect 8536 -7840 8585 -7806
rect 8619 -7840 8653 -7806
rect 8687 -7840 8736 -7806
rect 8536 -7887 8736 -7840
rect 8794 -7806 8994 -7790
rect 8794 -7840 8843 -7806
rect 8877 -7840 8911 -7806
rect 8945 -7840 8994 -7806
rect 8794 -7887 8994 -7840
rect 9246 -7806 9446 -7790
rect 9246 -7840 9295 -7806
rect 9329 -7840 9363 -7806
rect 9397 -7840 9446 -7806
rect 9246 -7887 9446 -7840
rect 1017 -8113 1217 -8087
rect 1469 -8113 1669 -8087
rect 1727 -8113 1927 -8087
rect 1985 -8113 2185 -8087
rect 2243 -8113 2443 -8087
rect 2695 -8113 2895 -8087
rect 2953 -8113 3153 -8087
rect 3211 -8113 3411 -8087
rect 3663 -8113 3863 -8087
rect 3921 -8113 4121 -8087
rect 4179 -8113 4379 -8087
rect 4437 -8113 4637 -8087
rect 4888 -8113 5088 -8087
rect 9734 -7806 9934 -7790
rect 9734 -7840 9783 -7806
rect 9817 -7840 9851 -7806
rect 9885 -7840 9934 -7806
rect 9734 -7887 9934 -7840
rect 10186 -7806 10386 -7790
rect 10186 -7840 10235 -7806
rect 10269 -7840 10303 -7806
rect 10337 -7840 10386 -7806
rect 10186 -7887 10386 -7840
rect 10444 -7806 10644 -7790
rect 10444 -7840 10493 -7806
rect 10527 -7840 10561 -7806
rect 10595 -7840 10644 -7806
rect 10444 -7887 10644 -7840
rect 10702 -7806 10902 -7790
rect 10702 -7840 10751 -7806
rect 10785 -7840 10819 -7806
rect 10853 -7840 10902 -7806
rect 10702 -7887 10902 -7840
rect 10960 -7806 11160 -7790
rect 10960 -7840 11009 -7806
rect 11043 -7840 11077 -7806
rect 11111 -7840 11160 -7806
rect 10960 -7887 11160 -7840
rect 11412 -7806 11612 -7790
rect 11412 -7840 11461 -7806
rect 11495 -7840 11529 -7806
rect 11563 -7840 11612 -7806
rect 11412 -7887 11612 -7840
rect 11670 -7806 11870 -7790
rect 11670 -7840 11719 -7806
rect 11753 -7840 11787 -7806
rect 11821 -7840 11870 -7806
rect 11670 -7887 11870 -7840
rect 11928 -7806 12128 -7790
rect 11928 -7840 11977 -7806
rect 12011 -7840 12045 -7806
rect 12079 -7840 12128 -7806
rect 11928 -7887 12128 -7840
rect 12380 -7806 12580 -7790
rect 12380 -7840 12429 -7806
rect 12463 -7840 12497 -7806
rect 12531 -7840 12580 -7806
rect 12380 -7887 12580 -7840
rect 12638 -7806 12838 -7790
rect 12638 -7840 12687 -7806
rect 12721 -7840 12755 -7806
rect 12789 -7840 12838 -7806
rect 12638 -7887 12838 -7840
rect 12896 -7806 13096 -7790
rect 12896 -7840 12945 -7806
rect 12979 -7840 13013 -7806
rect 13047 -7840 13096 -7806
rect 12896 -7887 13096 -7840
rect 13154 -7806 13354 -7790
rect 13154 -7840 13203 -7806
rect 13237 -7840 13271 -7806
rect 13305 -7840 13354 -7806
rect 13154 -7887 13354 -7840
rect 13606 -7806 13806 -7790
rect 13606 -7840 13655 -7806
rect 13689 -7840 13723 -7806
rect 13757 -7840 13806 -7806
rect 13606 -7887 13806 -7840
rect 5374 -8113 5574 -8087
rect 5826 -8113 6026 -8087
rect 6084 -8113 6284 -8087
rect 6342 -8113 6542 -8087
rect 6600 -8113 6800 -8087
rect 7052 -8113 7252 -8087
rect 7310 -8113 7510 -8087
rect 7568 -8113 7768 -8087
rect 8020 -8113 8220 -8087
rect 8278 -8113 8478 -8087
rect 8536 -8113 8736 -8087
rect 8794 -8113 8994 -8087
rect 9246 -8113 9446 -8087
rect 14092 -7806 14292 -7790
rect 14092 -7840 14141 -7806
rect 14175 -7840 14209 -7806
rect 14243 -7840 14292 -7806
rect 14092 -7887 14292 -7840
rect 14543 -7806 14743 -7790
rect 14543 -7840 14592 -7806
rect 14626 -7840 14660 -7806
rect 14694 -7840 14743 -7806
rect 14543 -7887 14743 -7840
rect 14801 -7806 15001 -7790
rect 14801 -7840 14850 -7806
rect 14884 -7840 14918 -7806
rect 14952 -7840 15001 -7806
rect 14801 -7887 15001 -7840
rect 15059 -7806 15259 -7790
rect 15059 -7840 15108 -7806
rect 15142 -7840 15176 -7806
rect 15210 -7840 15259 -7806
rect 15059 -7887 15259 -7840
rect 15317 -7806 15517 -7790
rect 15317 -7840 15366 -7806
rect 15400 -7840 15434 -7806
rect 15468 -7840 15517 -7806
rect 15317 -7887 15517 -7840
rect 15769 -7806 15969 -7790
rect 15769 -7840 15818 -7806
rect 15852 -7840 15886 -7806
rect 15920 -7840 15969 -7806
rect 15769 -7887 15969 -7840
rect 16027 -7806 16227 -7790
rect 16027 -7840 16076 -7806
rect 16110 -7840 16144 -7806
rect 16178 -7840 16227 -7806
rect 16027 -7887 16227 -7840
rect 16285 -7806 16485 -7790
rect 16285 -7840 16334 -7806
rect 16368 -7840 16402 -7806
rect 16436 -7840 16485 -7806
rect 16285 -7887 16485 -7840
rect 16737 -7806 16937 -7790
rect 16737 -7840 16786 -7806
rect 16820 -7840 16854 -7806
rect 16888 -7840 16937 -7806
rect 16737 -7887 16937 -7840
rect 16995 -7806 17195 -7790
rect 16995 -7840 17044 -7806
rect 17078 -7840 17112 -7806
rect 17146 -7840 17195 -7806
rect 16995 -7887 17195 -7840
rect 17253 -7806 17453 -7790
rect 17253 -7840 17302 -7806
rect 17336 -7840 17370 -7806
rect 17404 -7840 17453 -7806
rect 17253 -7887 17453 -7840
rect 17511 -7806 17711 -7790
rect 17511 -7840 17560 -7806
rect 17594 -7840 17628 -7806
rect 17662 -7840 17711 -7806
rect 17511 -7887 17711 -7840
rect 17963 -7806 18163 -7790
rect 17963 -7840 18012 -7806
rect 18046 -7840 18080 -7806
rect 18114 -7840 18163 -7806
rect 17963 -7887 18163 -7840
rect 9734 -8113 9934 -8087
rect 10186 -8113 10386 -8087
rect 10444 -8113 10644 -8087
rect 10702 -8113 10902 -8087
rect 10960 -8113 11160 -8087
rect 11412 -8113 11612 -8087
rect 11670 -8113 11870 -8087
rect 11928 -8113 12128 -8087
rect 12380 -8113 12580 -8087
rect 12638 -8113 12838 -8087
rect 12896 -8113 13096 -8087
rect 13154 -8113 13354 -8087
rect 13606 -8113 13806 -8087
rect 14092 -8113 14292 -8087
rect 14543 -8113 14743 -8087
rect 14801 -8113 15001 -8087
rect 15059 -8113 15259 -8087
rect 15317 -8113 15517 -8087
rect 15769 -8113 15969 -8087
rect 16027 -8113 16227 -8087
rect 16285 -8113 16485 -8087
rect 16737 -8113 16937 -8087
rect 16995 -8113 17195 -8087
rect 17253 -8113 17453 -8087
rect 17511 -8113 17711 -8087
rect 17963 -8113 18163 -8087
rect 1017 -8831 1217 -8805
rect 1469 -8831 1669 -8805
rect 1727 -8831 1927 -8805
rect 1985 -8831 2185 -8805
rect 2243 -8831 2443 -8805
rect 2695 -8831 2895 -8805
rect 2953 -8831 3153 -8805
rect 3211 -8831 3411 -8805
rect 3663 -8831 3863 -8805
rect 3921 -8831 4121 -8805
rect 4179 -8831 4379 -8805
rect 4437 -8831 4637 -8805
rect 4888 -8831 5088 -8805
rect 5374 -8831 5574 -8805
rect 5826 -8831 6026 -8805
rect 6084 -8831 6284 -8805
rect 6342 -8831 6542 -8805
rect 6600 -8831 6800 -8805
rect 7052 -8831 7252 -8805
rect 7310 -8831 7510 -8805
rect 7568 -8831 7768 -8805
rect 8020 -8831 8220 -8805
rect 8278 -8831 8478 -8805
rect 8536 -8831 8736 -8805
rect 8794 -8831 8994 -8805
rect 9246 -8831 9446 -8805
rect 1017 -9078 1217 -9031
rect 1017 -9112 1066 -9078
rect 1100 -9112 1134 -9078
rect 1168 -9112 1217 -9078
rect 1017 -9128 1217 -9112
rect 1469 -9078 1669 -9031
rect 1469 -9112 1518 -9078
rect 1552 -9112 1586 -9078
rect 1620 -9112 1669 -9078
rect 1469 -9128 1669 -9112
rect 1727 -9078 1927 -9031
rect 1727 -9112 1776 -9078
rect 1810 -9112 1844 -9078
rect 1878 -9112 1927 -9078
rect 1727 -9128 1927 -9112
rect 1985 -9078 2185 -9031
rect 1985 -9112 2034 -9078
rect 2068 -9112 2102 -9078
rect 2136 -9112 2185 -9078
rect 1985 -9128 2185 -9112
rect 2243 -9078 2443 -9031
rect 2243 -9112 2292 -9078
rect 2326 -9112 2360 -9078
rect 2394 -9112 2443 -9078
rect 2243 -9128 2443 -9112
rect 2695 -9078 2895 -9031
rect 2695 -9112 2744 -9078
rect 2778 -9112 2812 -9078
rect 2846 -9112 2895 -9078
rect 2695 -9128 2895 -9112
rect 2953 -9078 3153 -9031
rect 2953 -9112 3002 -9078
rect 3036 -9112 3070 -9078
rect 3104 -9112 3153 -9078
rect 2953 -9128 3153 -9112
rect 3211 -9078 3411 -9031
rect 3211 -9112 3260 -9078
rect 3294 -9112 3328 -9078
rect 3362 -9112 3411 -9078
rect 3211 -9128 3411 -9112
rect 3663 -9078 3863 -9031
rect 3663 -9112 3712 -9078
rect 3746 -9112 3780 -9078
rect 3814 -9112 3863 -9078
rect 3663 -9128 3863 -9112
rect 3921 -9078 4121 -9031
rect 3921 -9112 3970 -9078
rect 4004 -9112 4038 -9078
rect 4072 -9112 4121 -9078
rect 3921 -9128 4121 -9112
rect 4179 -9078 4379 -9031
rect 4179 -9112 4228 -9078
rect 4262 -9112 4296 -9078
rect 4330 -9112 4379 -9078
rect 4179 -9128 4379 -9112
rect 4437 -9078 4637 -9031
rect 4437 -9112 4486 -9078
rect 4520 -9112 4554 -9078
rect 4588 -9112 4637 -9078
rect 4437 -9128 4637 -9112
rect 4888 -9078 5088 -9031
rect 4888 -9112 4937 -9078
rect 4971 -9112 5005 -9078
rect 5039 -9112 5088 -9078
rect 4888 -9128 5088 -9112
rect 9734 -8831 9934 -8805
rect 10186 -8831 10386 -8805
rect 10444 -8831 10644 -8805
rect 10702 -8831 10902 -8805
rect 10960 -8831 11160 -8805
rect 11412 -8831 11612 -8805
rect 11670 -8831 11870 -8805
rect 11928 -8831 12128 -8805
rect 12380 -8831 12580 -8805
rect 12638 -8831 12838 -8805
rect 12896 -8831 13096 -8805
rect 13154 -8831 13354 -8805
rect 13606 -8831 13806 -8805
rect 5374 -9078 5574 -9031
rect 5374 -9112 5423 -9078
rect 5457 -9112 5491 -9078
rect 5525 -9112 5574 -9078
rect 5374 -9128 5574 -9112
rect 5826 -9078 6026 -9031
rect 5826 -9112 5875 -9078
rect 5909 -9112 5943 -9078
rect 5977 -9112 6026 -9078
rect 5826 -9128 6026 -9112
rect 6084 -9078 6284 -9031
rect 6084 -9112 6133 -9078
rect 6167 -9112 6201 -9078
rect 6235 -9112 6284 -9078
rect 6084 -9128 6284 -9112
rect 6342 -9078 6542 -9031
rect 6342 -9112 6391 -9078
rect 6425 -9112 6459 -9078
rect 6493 -9112 6542 -9078
rect 6342 -9128 6542 -9112
rect 6600 -9078 6800 -9031
rect 6600 -9112 6649 -9078
rect 6683 -9112 6717 -9078
rect 6751 -9112 6800 -9078
rect 6600 -9128 6800 -9112
rect 7052 -9078 7252 -9031
rect 7052 -9112 7101 -9078
rect 7135 -9112 7169 -9078
rect 7203 -9112 7252 -9078
rect 7052 -9128 7252 -9112
rect 7310 -9078 7510 -9031
rect 7310 -9112 7359 -9078
rect 7393 -9112 7427 -9078
rect 7461 -9112 7510 -9078
rect 7310 -9128 7510 -9112
rect 7568 -9078 7768 -9031
rect 7568 -9112 7617 -9078
rect 7651 -9112 7685 -9078
rect 7719 -9112 7768 -9078
rect 7568 -9128 7768 -9112
rect 8020 -9078 8220 -9031
rect 8020 -9112 8069 -9078
rect 8103 -9112 8137 -9078
rect 8171 -9112 8220 -9078
rect 8020 -9128 8220 -9112
rect 8278 -9078 8478 -9031
rect 8278 -9112 8327 -9078
rect 8361 -9112 8395 -9078
rect 8429 -9112 8478 -9078
rect 8278 -9128 8478 -9112
rect 8536 -9078 8736 -9031
rect 8536 -9112 8585 -9078
rect 8619 -9112 8653 -9078
rect 8687 -9112 8736 -9078
rect 8536 -9128 8736 -9112
rect 8794 -9078 8994 -9031
rect 8794 -9112 8843 -9078
rect 8877 -9112 8911 -9078
rect 8945 -9112 8994 -9078
rect 8794 -9128 8994 -9112
rect 9246 -9078 9446 -9031
rect 9246 -9112 9295 -9078
rect 9329 -9112 9363 -9078
rect 9397 -9112 9446 -9078
rect 9246 -9128 9446 -9112
rect 14092 -8831 14292 -8805
rect 14543 -8831 14743 -8805
rect 14801 -8831 15001 -8805
rect 15059 -8831 15259 -8805
rect 15317 -8831 15517 -8805
rect 15769 -8831 15969 -8805
rect 16027 -8831 16227 -8805
rect 16285 -8831 16485 -8805
rect 16737 -8831 16937 -8805
rect 16995 -8831 17195 -8805
rect 17253 -8831 17453 -8805
rect 17511 -8831 17711 -8805
rect 17963 -8831 18163 -8805
rect 9734 -9078 9934 -9031
rect 9734 -9112 9783 -9078
rect 9817 -9112 9851 -9078
rect 9885 -9112 9934 -9078
rect 9734 -9128 9934 -9112
rect 10186 -9078 10386 -9031
rect 10186 -9112 10235 -9078
rect 10269 -9112 10303 -9078
rect 10337 -9112 10386 -9078
rect 10186 -9128 10386 -9112
rect 10444 -9078 10644 -9031
rect 10444 -9112 10493 -9078
rect 10527 -9112 10561 -9078
rect 10595 -9112 10644 -9078
rect 10444 -9128 10644 -9112
rect 10702 -9078 10902 -9031
rect 10702 -9112 10751 -9078
rect 10785 -9112 10819 -9078
rect 10853 -9112 10902 -9078
rect 10702 -9128 10902 -9112
rect 10960 -9078 11160 -9031
rect 10960 -9112 11009 -9078
rect 11043 -9112 11077 -9078
rect 11111 -9112 11160 -9078
rect 10960 -9128 11160 -9112
rect 11412 -9078 11612 -9031
rect 11412 -9112 11461 -9078
rect 11495 -9112 11529 -9078
rect 11563 -9112 11612 -9078
rect 11412 -9128 11612 -9112
rect 11670 -9078 11870 -9031
rect 11670 -9112 11719 -9078
rect 11753 -9112 11787 -9078
rect 11821 -9112 11870 -9078
rect 11670 -9128 11870 -9112
rect 11928 -9078 12128 -9031
rect 11928 -9112 11977 -9078
rect 12011 -9112 12045 -9078
rect 12079 -9112 12128 -9078
rect 11928 -9128 12128 -9112
rect 12380 -9078 12580 -9031
rect 12380 -9112 12429 -9078
rect 12463 -9112 12497 -9078
rect 12531 -9112 12580 -9078
rect 12380 -9128 12580 -9112
rect 12638 -9078 12838 -9031
rect 12638 -9112 12687 -9078
rect 12721 -9112 12755 -9078
rect 12789 -9112 12838 -9078
rect 12638 -9128 12838 -9112
rect 12896 -9078 13096 -9031
rect 12896 -9112 12945 -9078
rect 12979 -9112 13013 -9078
rect 13047 -9112 13096 -9078
rect 12896 -9128 13096 -9112
rect 13154 -9078 13354 -9031
rect 13154 -9112 13203 -9078
rect 13237 -9112 13271 -9078
rect 13305 -9112 13354 -9078
rect 13154 -9128 13354 -9112
rect 13606 -9078 13806 -9031
rect 13606 -9112 13655 -9078
rect 13689 -9112 13723 -9078
rect 13757 -9112 13806 -9078
rect 13606 -9128 13806 -9112
rect 14092 -9078 14292 -9031
rect 14092 -9112 14141 -9078
rect 14175 -9112 14209 -9078
rect 14243 -9112 14292 -9078
rect 14092 -9128 14292 -9112
rect 14543 -9078 14743 -9031
rect 14543 -9112 14592 -9078
rect 14626 -9112 14660 -9078
rect 14694 -9112 14743 -9078
rect 14543 -9128 14743 -9112
rect 14801 -9078 15001 -9031
rect 14801 -9112 14850 -9078
rect 14884 -9112 14918 -9078
rect 14952 -9112 15001 -9078
rect 14801 -9128 15001 -9112
rect 15059 -9078 15259 -9031
rect 15059 -9112 15108 -9078
rect 15142 -9112 15176 -9078
rect 15210 -9112 15259 -9078
rect 15059 -9128 15259 -9112
rect 15317 -9078 15517 -9031
rect 15317 -9112 15366 -9078
rect 15400 -9112 15434 -9078
rect 15468 -9112 15517 -9078
rect 15317 -9128 15517 -9112
rect 15769 -9078 15969 -9031
rect 15769 -9112 15818 -9078
rect 15852 -9112 15886 -9078
rect 15920 -9112 15969 -9078
rect 15769 -9128 15969 -9112
rect 16027 -9078 16227 -9031
rect 16027 -9112 16076 -9078
rect 16110 -9112 16144 -9078
rect 16178 -9112 16227 -9078
rect 16027 -9128 16227 -9112
rect 16285 -9078 16485 -9031
rect 16285 -9112 16334 -9078
rect 16368 -9112 16402 -9078
rect 16436 -9112 16485 -9078
rect 16285 -9128 16485 -9112
rect 16737 -9078 16937 -9031
rect 16737 -9112 16786 -9078
rect 16820 -9112 16854 -9078
rect 16888 -9112 16937 -9078
rect 16737 -9128 16937 -9112
rect 16995 -9078 17195 -9031
rect 16995 -9112 17044 -9078
rect 17078 -9112 17112 -9078
rect 17146 -9112 17195 -9078
rect 16995 -9128 17195 -9112
rect 17253 -9078 17453 -9031
rect 17253 -9112 17302 -9078
rect 17336 -9112 17370 -9078
rect 17404 -9112 17453 -9078
rect 17253 -9128 17453 -9112
rect 17511 -9078 17711 -9031
rect 17511 -9112 17560 -9078
rect 17594 -9112 17628 -9078
rect 17662 -9112 17711 -9078
rect 17511 -9128 17711 -9112
rect 17963 -9078 18163 -9031
rect 17963 -9112 18012 -9078
rect 18046 -9112 18080 -9078
rect 18114 -9112 18163 -9078
rect 17963 -9128 18163 -9112
<< polycont >>
rect 1066 315 1100 349
rect 1134 315 1168 349
rect 1518 315 1552 349
rect 1586 315 1620 349
rect 1776 315 1810 349
rect 1844 315 1878 349
rect 2034 315 2068 349
rect 2102 315 2136 349
rect 2292 315 2326 349
rect 2360 315 2394 349
rect 2744 315 2778 349
rect 2812 315 2846 349
rect 3002 315 3036 349
rect 3070 315 3104 349
rect 3260 315 3294 349
rect 3328 315 3362 349
rect 3712 315 3746 349
rect 3780 315 3814 349
rect 3970 315 4004 349
rect 4038 315 4072 349
rect 4228 315 4262 349
rect 4296 315 4330 349
rect 4486 315 4520 349
rect 4554 315 4588 349
rect 4937 315 4971 349
rect 5005 315 5039 349
rect 5423 315 5457 349
rect 5491 315 5525 349
rect 5875 315 5909 349
rect 5943 315 5977 349
rect 6133 315 6167 349
rect 6201 315 6235 349
rect 6391 315 6425 349
rect 6459 315 6493 349
rect 6649 315 6683 349
rect 6717 315 6751 349
rect 7101 315 7135 349
rect 7169 315 7203 349
rect 7359 315 7393 349
rect 7427 315 7461 349
rect 7617 315 7651 349
rect 7685 315 7719 349
rect 8069 315 8103 349
rect 8137 315 8171 349
rect 8327 315 8361 349
rect 8395 315 8429 349
rect 8585 315 8619 349
rect 8653 315 8687 349
rect 8843 315 8877 349
rect 8911 315 8945 349
rect 9295 315 9329 349
rect 9363 315 9397 349
rect 9783 315 9817 349
rect 9851 315 9885 349
rect 10235 315 10269 349
rect 10303 315 10337 349
rect 10493 315 10527 349
rect 10561 315 10595 349
rect 10751 315 10785 349
rect 10819 315 10853 349
rect 11009 315 11043 349
rect 11077 315 11111 349
rect 11461 315 11495 349
rect 11529 315 11563 349
rect 11719 315 11753 349
rect 11787 315 11821 349
rect 11977 315 12011 349
rect 12045 315 12079 349
rect 12429 315 12463 349
rect 12497 315 12531 349
rect 12687 315 12721 349
rect 12755 315 12789 349
rect 12945 315 12979 349
rect 13013 315 13047 349
rect 13203 315 13237 349
rect 13271 315 13305 349
rect 13655 315 13689 349
rect 13723 315 13757 349
rect 14141 315 14175 349
rect 14209 315 14243 349
rect 14592 315 14626 349
rect 14660 315 14694 349
rect 14850 315 14884 349
rect 14918 315 14952 349
rect 15108 315 15142 349
rect 15176 315 15210 349
rect 15366 315 15400 349
rect 15434 315 15468 349
rect 15818 315 15852 349
rect 15886 315 15920 349
rect 16076 315 16110 349
rect 16144 315 16178 349
rect 16334 315 16368 349
rect 16402 315 16436 349
rect 16786 315 16820 349
rect 16854 315 16888 349
rect 17044 315 17078 349
rect 17112 315 17146 349
rect 17302 315 17336 349
rect 17370 315 17404 349
rect 17560 315 17594 349
rect 17628 315 17662 349
rect 18012 315 18046 349
rect 18080 315 18114 349
rect 1066 -957 1100 -923
rect 1134 -957 1168 -923
rect 1518 -957 1552 -923
rect 1586 -957 1620 -923
rect 1776 -957 1810 -923
rect 1844 -957 1878 -923
rect 2034 -957 2068 -923
rect 2102 -957 2136 -923
rect 2292 -957 2326 -923
rect 2360 -957 2394 -923
rect 2744 -957 2778 -923
rect 2812 -957 2846 -923
rect 3002 -957 3036 -923
rect 3070 -957 3104 -923
rect 3260 -957 3294 -923
rect 3328 -957 3362 -923
rect 3712 -957 3746 -923
rect 3780 -957 3814 -923
rect 3970 -957 4004 -923
rect 4038 -957 4072 -923
rect 4228 -957 4262 -923
rect 4296 -957 4330 -923
rect 4486 -957 4520 -923
rect 4554 -957 4588 -923
rect 4937 -957 4971 -923
rect 5005 -957 5039 -923
rect 5423 -957 5457 -923
rect 5491 -957 5525 -923
rect 5875 -957 5909 -923
rect 5943 -957 5977 -923
rect 6133 -957 6167 -923
rect 6201 -957 6235 -923
rect 6391 -957 6425 -923
rect 6459 -957 6493 -923
rect 6649 -957 6683 -923
rect 6717 -957 6751 -923
rect 7101 -957 7135 -923
rect 7169 -957 7203 -923
rect 7359 -957 7393 -923
rect 7427 -957 7461 -923
rect 7617 -957 7651 -923
rect 7685 -957 7719 -923
rect 8069 -957 8103 -923
rect 8137 -957 8171 -923
rect 8327 -957 8361 -923
rect 8395 -957 8429 -923
rect 8585 -957 8619 -923
rect 8653 -957 8687 -923
rect 8843 -957 8877 -923
rect 8911 -957 8945 -923
rect 9295 -957 9329 -923
rect 9363 -957 9397 -923
rect 1066 -1320 1100 -1286
rect 1134 -1320 1168 -1286
rect 1518 -1320 1552 -1286
rect 1586 -1320 1620 -1286
rect 1776 -1320 1810 -1286
rect 1844 -1320 1878 -1286
rect 2034 -1320 2068 -1286
rect 2102 -1320 2136 -1286
rect 2292 -1320 2326 -1286
rect 2360 -1320 2394 -1286
rect 2744 -1320 2778 -1286
rect 2812 -1320 2846 -1286
rect 3002 -1320 3036 -1286
rect 3070 -1320 3104 -1286
rect 3260 -1320 3294 -1286
rect 3328 -1320 3362 -1286
rect 3712 -1320 3746 -1286
rect 3780 -1320 3814 -1286
rect 3970 -1320 4004 -1286
rect 4038 -1320 4072 -1286
rect 4228 -1320 4262 -1286
rect 4296 -1320 4330 -1286
rect 4486 -1320 4520 -1286
rect 4554 -1320 4588 -1286
rect 4937 -1320 4971 -1286
rect 5005 -1320 5039 -1286
rect 9783 -957 9817 -923
rect 9851 -957 9885 -923
rect 10235 -957 10269 -923
rect 10303 -957 10337 -923
rect 10493 -957 10527 -923
rect 10561 -957 10595 -923
rect 10751 -957 10785 -923
rect 10819 -957 10853 -923
rect 11009 -957 11043 -923
rect 11077 -957 11111 -923
rect 11461 -957 11495 -923
rect 11529 -957 11563 -923
rect 11719 -957 11753 -923
rect 11787 -957 11821 -923
rect 11977 -957 12011 -923
rect 12045 -957 12079 -923
rect 12429 -957 12463 -923
rect 12497 -957 12531 -923
rect 12687 -957 12721 -923
rect 12755 -957 12789 -923
rect 12945 -957 12979 -923
rect 13013 -957 13047 -923
rect 13203 -957 13237 -923
rect 13271 -957 13305 -923
rect 13655 -957 13689 -923
rect 13723 -957 13757 -923
rect 5423 -1320 5457 -1286
rect 5491 -1320 5525 -1286
rect 5875 -1320 5909 -1286
rect 5943 -1320 5977 -1286
rect 6133 -1320 6167 -1286
rect 6201 -1320 6235 -1286
rect 6391 -1320 6425 -1286
rect 6459 -1320 6493 -1286
rect 6649 -1320 6683 -1286
rect 6717 -1320 6751 -1286
rect 7101 -1320 7135 -1286
rect 7169 -1320 7203 -1286
rect 7359 -1320 7393 -1286
rect 7427 -1320 7461 -1286
rect 7617 -1320 7651 -1286
rect 7685 -1320 7719 -1286
rect 8069 -1320 8103 -1286
rect 8137 -1320 8171 -1286
rect 8327 -1320 8361 -1286
rect 8395 -1320 8429 -1286
rect 8585 -1320 8619 -1286
rect 8653 -1320 8687 -1286
rect 8843 -1320 8877 -1286
rect 8911 -1320 8945 -1286
rect 9295 -1320 9329 -1286
rect 9363 -1320 9397 -1286
rect 14141 -957 14175 -923
rect 14209 -957 14243 -923
rect 14592 -957 14626 -923
rect 14660 -957 14694 -923
rect 14850 -957 14884 -923
rect 14918 -957 14952 -923
rect 15108 -957 15142 -923
rect 15176 -957 15210 -923
rect 15366 -957 15400 -923
rect 15434 -957 15468 -923
rect 15818 -957 15852 -923
rect 15886 -957 15920 -923
rect 16076 -957 16110 -923
rect 16144 -957 16178 -923
rect 16334 -957 16368 -923
rect 16402 -957 16436 -923
rect 16786 -957 16820 -923
rect 16854 -957 16888 -923
rect 17044 -957 17078 -923
rect 17112 -957 17146 -923
rect 17302 -957 17336 -923
rect 17370 -957 17404 -923
rect 17560 -957 17594 -923
rect 17628 -957 17662 -923
rect 18012 -957 18046 -923
rect 18080 -957 18114 -923
rect 9783 -1320 9817 -1286
rect 9851 -1320 9885 -1286
rect 10235 -1320 10269 -1286
rect 10303 -1320 10337 -1286
rect 10493 -1320 10527 -1286
rect 10561 -1320 10595 -1286
rect 10751 -1320 10785 -1286
rect 10819 -1320 10853 -1286
rect 11009 -1320 11043 -1286
rect 11077 -1320 11111 -1286
rect 11461 -1320 11495 -1286
rect 11529 -1320 11563 -1286
rect 11719 -1320 11753 -1286
rect 11787 -1320 11821 -1286
rect 11977 -1320 12011 -1286
rect 12045 -1320 12079 -1286
rect 12429 -1320 12463 -1286
rect 12497 -1320 12531 -1286
rect 12687 -1320 12721 -1286
rect 12755 -1320 12789 -1286
rect 12945 -1320 12979 -1286
rect 13013 -1320 13047 -1286
rect 13203 -1320 13237 -1286
rect 13271 -1320 13305 -1286
rect 13655 -1320 13689 -1286
rect 13723 -1320 13757 -1286
rect 14141 -1320 14175 -1286
rect 14209 -1320 14243 -1286
rect 14592 -1320 14626 -1286
rect 14660 -1320 14694 -1286
rect 14850 -1320 14884 -1286
rect 14918 -1320 14952 -1286
rect 15108 -1320 15142 -1286
rect 15176 -1320 15210 -1286
rect 15366 -1320 15400 -1286
rect 15434 -1320 15468 -1286
rect 15818 -1320 15852 -1286
rect 15886 -1320 15920 -1286
rect 16076 -1320 16110 -1286
rect 16144 -1320 16178 -1286
rect 16334 -1320 16368 -1286
rect 16402 -1320 16436 -1286
rect 16786 -1320 16820 -1286
rect 16854 -1320 16888 -1286
rect 17044 -1320 17078 -1286
rect 17112 -1320 17146 -1286
rect 17302 -1320 17336 -1286
rect 17370 -1320 17404 -1286
rect 17560 -1320 17594 -1286
rect 17628 -1320 17662 -1286
rect 18012 -1320 18046 -1286
rect 18080 -1320 18114 -1286
rect 1066 -2604 1100 -2570
rect 1134 -2604 1168 -2570
rect 1518 -2604 1552 -2570
rect 1586 -2604 1620 -2570
rect 1776 -2604 1810 -2570
rect 1844 -2604 1878 -2570
rect 2034 -2604 2068 -2570
rect 2102 -2604 2136 -2570
rect 2292 -2604 2326 -2570
rect 2360 -2604 2394 -2570
rect 2744 -2604 2778 -2570
rect 2812 -2604 2846 -2570
rect 3002 -2604 3036 -2570
rect 3070 -2604 3104 -2570
rect 3260 -2604 3294 -2570
rect 3328 -2604 3362 -2570
rect 3712 -2604 3746 -2570
rect 3780 -2604 3814 -2570
rect 3970 -2604 4004 -2570
rect 4038 -2604 4072 -2570
rect 4228 -2604 4262 -2570
rect 4296 -2604 4330 -2570
rect 4486 -2604 4520 -2570
rect 4554 -2604 4588 -2570
rect 4937 -2604 4971 -2570
rect 5005 -2604 5039 -2570
rect 5423 -2604 5457 -2570
rect 5491 -2604 5525 -2570
rect 5875 -2604 5909 -2570
rect 5943 -2604 5977 -2570
rect 6133 -2604 6167 -2570
rect 6201 -2604 6235 -2570
rect 6391 -2604 6425 -2570
rect 6459 -2604 6493 -2570
rect 6649 -2604 6683 -2570
rect 6717 -2604 6751 -2570
rect 7101 -2604 7135 -2570
rect 7169 -2604 7203 -2570
rect 7359 -2604 7393 -2570
rect 7427 -2604 7461 -2570
rect 7617 -2604 7651 -2570
rect 7685 -2604 7719 -2570
rect 8069 -2604 8103 -2570
rect 8137 -2604 8171 -2570
rect 8327 -2604 8361 -2570
rect 8395 -2604 8429 -2570
rect 8585 -2604 8619 -2570
rect 8653 -2604 8687 -2570
rect 8843 -2604 8877 -2570
rect 8911 -2604 8945 -2570
rect 9295 -2604 9329 -2570
rect 9363 -2604 9397 -2570
rect 1066 -2967 1100 -2933
rect 1134 -2967 1168 -2933
rect 1518 -2967 1552 -2933
rect 1586 -2967 1620 -2933
rect 1776 -2967 1810 -2933
rect 1844 -2967 1878 -2933
rect 2034 -2967 2068 -2933
rect 2102 -2967 2136 -2933
rect 2292 -2967 2326 -2933
rect 2360 -2967 2394 -2933
rect 2744 -2967 2778 -2933
rect 2812 -2967 2846 -2933
rect 3002 -2967 3036 -2933
rect 3070 -2967 3104 -2933
rect 3260 -2967 3294 -2933
rect 3328 -2967 3362 -2933
rect 3712 -2967 3746 -2933
rect 3780 -2967 3814 -2933
rect 3970 -2967 4004 -2933
rect 4038 -2967 4072 -2933
rect 4228 -2967 4262 -2933
rect 4296 -2967 4330 -2933
rect 4486 -2967 4520 -2933
rect 4554 -2967 4588 -2933
rect 4937 -2967 4971 -2933
rect 5005 -2967 5039 -2933
rect 9783 -2604 9817 -2570
rect 9851 -2604 9885 -2570
rect 10235 -2604 10269 -2570
rect 10303 -2604 10337 -2570
rect 10493 -2604 10527 -2570
rect 10561 -2604 10595 -2570
rect 10751 -2604 10785 -2570
rect 10819 -2604 10853 -2570
rect 11009 -2604 11043 -2570
rect 11077 -2604 11111 -2570
rect 11461 -2604 11495 -2570
rect 11529 -2604 11563 -2570
rect 11719 -2604 11753 -2570
rect 11787 -2604 11821 -2570
rect 11977 -2604 12011 -2570
rect 12045 -2604 12079 -2570
rect 12429 -2604 12463 -2570
rect 12497 -2604 12531 -2570
rect 12687 -2604 12721 -2570
rect 12755 -2604 12789 -2570
rect 12945 -2604 12979 -2570
rect 13013 -2604 13047 -2570
rect 13203 -2604 13237 -2570
rect 13271 -2604 13305 -2570
rect 13655 -2604 13689 -2570
rect 13723 -2604 13757 -2570
rect 5423 -2967 5457 -2933
rect 5491 -2967 5525 -2933
rect 5875 -2967 5909 -2933
rect 5943 -2967 5977 -2933
rect 6133 -2967 6167 -2933
rect 6201 -2967 6235 -2933
rect 6391 -2967 6425 -2933
rect 6459 -2967 6493 -2933
rect 6649 -2967 6683 -2933
rect 6717 -2967 6751 -2933
rect 7101 -2967 7135 -2933
rect 7169 -2967 7203 -2933
rect 7359 -2967 7393 -2933
rect 7427 -2967 7461 -2933
rect 7617 -2967 7651 -2933
rect 7685 -2967 7719 -2933
rect 8069 -2967 8103 -2933
rect 8137 -2967 8171 -2933
rect 8327 -2967 8361 -2933
rect 8395 -2967 8429 -2933
rect 8585 -2967 8619 -2933
rect 8653 -2967 8687 -2933
rect 8843 -2967 8877 -2933
rect 8911 -2967 8945 -2933
rect 9295 -2967 9329 -2933
rect 9363 -2967 9397 -2933
rect 14141 -2604 14175 -2570
rect 14209 -2604 14243 -2570
rect 14592 -2604 14626 -2570
rect 14660 -2604 14694 -2570
rect 14850 -2604 14884 -2570
rect 14918 -2604 14952 -2570
rect 15108 -2604 15142 -2570
rect 15176 -2604 15210 -2570
rect 15366 -2604 15400 -2570
rect 15434 -2604 15468 -2570
rect 15818 -2604 15852 -2570
rect 15886 -2604 15920 -2570
rect 16076 -2604 16110 -2570
rect 16144 -2604 16178 -2570
rect 16334 -2604 16368 -2570
rect 16402 -2604 16436 -2570
rect 16786 -2604 16820 -2570
rect 16854 -2604 16888 -2570
rect 17044 -2604 17078 -2570
rect 17112 -2604 17146 -2570
rect 17302 -2604 17336 -2570
rect 17370 -2604 17404 -2570
rect 17560 -2604 17594 -2570
rect 17628 -2604 17662 -2570
rect 18012 -2604 18046 -2570
rect 18080 -2604 18114 -2570
rect 9783 -2967 9817 -2933
rect 9851 -2967 9885 -2933
rect 10235 -2967 10269 -2933
rect 10303 -2967 10337 -2933
rect 10493 -2967 10527 -2933
rect 10561 -2967 10595 -2933
rect 10751 -2967 10785 -2933
rect 10819 -2967 10853 -2933
rect 11009 -2967 11043 -2933
rect 11077 -2967 11111 -2933
rect 11461 -2967 11495 -2933
rect 11529 -2967 11563 -2933
rect 11719 -2967 11753 -2933
rect 11787 -2967 11821 -2933
rect 11977 -2967 12011 -2933
rect 12045 -2967 12079 -2933
rect 12429 -2967 12463 -2933
rect 12497 -2967 12531 -2933
rect 12687 -2967 12721 -2933
rect 12755 -2967 12789 -2933
rect 12945 -2967 12979 -2933
rect 13013 -2967 13047 -2933
rect 13203 -2967 13237 -2933
rect 13271 -2967 13305 -2933
rect 13655 -2967 13689 -2933
rect 13723 -2967 13757 -2933
rect 14141 -2967 14175 -2933
rect 14209 -2967 14243 -2933
rect 14592 -2967 14626 -2933
rect 14660 -2967 14694 -2933
rect 14850 -2967 14884 -2933
rect 14918 -2967 14952 -2933
rect 15108 -2967 15142 -2933
rect 15176 -2967 15210 -2933
rect 15366 -2967 15400 -2933
rect 15434 -2967 15468 -2933
rect 15818 -2967 15852 -2933
rect 15886 -2967 15920 -2933
rect 16076 -2967 16110 -2933
rect 16144 -2967 16178 -2933
rect 16334 -2967 16368 -2933
rect 16402 -2967 16436 -2933
rect 16786 -2967 16820 -2933
rect 16854 -2967 16888 -2933
rect 17044 -2967 17078 -2933
rect 17112 -2967 17146 -2933
rect 17302 -2967 17336 -2933
rect 17370 -2967 17404 -2933
rect 17560 -2967 17594 -2933
rect 17628 -2967 17662 -2933
rect 18012 -2967 18046 -2933
rect 18080 -2967 18114 -2933
rect 1066 -4285 1100 -4251
rect 1134 -4285 1168 -4251
rect 1518 -4285 1552 -4251
rect 1586 -4285 1620 -4251
rect 1776 -4285 1810 -4251
rect 1844 -4285 1878 -4251
rect 2034 -4285 2068 -4251
rect 2102 -4285 2136 -4251
rect 2292 -4285 2326 -4251
rect 2360 -4285 2394 -4251
rect 2744 -4285 2778 -4251
rect 2812 -4285 2846 -4251
rect 3002 -4285 3036 -4251
rect 3070 -4285 3104 -4251
rect 3260 -4285 3294 -4251
rect 3328 -4285 3362 -4251
rect 3712 -4285 3746 -4251
rect 3780 -4285 3814 -4251
rect 3970 -4285 4004 -4251
rect 4038 -4285 4072 -4251
rect 4228 -4285 4262 -4251
rect 4296 -4285 4330 -4251
rect 4486 -4285 4520 -4251
rect 4554 -4285 4588 -4251
rect 4937 -4285 4971 -4251
rect 5005 -4285 5039 -4251
rect 5423 -4285 5457 -4251
rect 5491 -4285 5525 -4251
rect 5875 -4285 5909 -4251
rect 5943 -4285 5977 -4251
rect 6133 -4285 6167 -4251
rect 6201 -4285 6235 -4251
rect 6391 -4285 6425 -4251
rect 6459 -4285 6493 -4251
rect 6649 -4285 6683 -4251
rect 6717 -4285 6751 -4251
rect 7101 -4285 7135 -4251
rect 7169 -4285 7203 -4251
rect 7359 -4285 7393 -4251
rect 7427 -4285 7461 -4251
rect 7617 -4285 7651 -4251
rect 7685 -4285 7719 -4251
rect 8069 -4285 8103 -4251
rect 8137 -4285 8171 -4251
rect 8327 -4285 8361 -4251
rect 8395 -4285 8429 -4251
rect 8585 -4285 8619 -4251
rect 8653 -4285 8687 -4251
rect 8843 -4285 8877 -4251
rect 8911 -4285 8945 -4251
rect 9295 -4285 9329 -4251
rect 9363 -4285 9397 -4251
rect 9783 -4285 9817 -4251
rect 9851 -4285 9885 -4251
rect 10235 -4285 10269 -4251
rect 10303 -4285 10337 -4251
rect 10493 -4285 10527 -4251
rect 10561 -4285 10595 -4251
rect 10751 -4285 10785 -4251
rect 10819 -4285 10853 -4251
rect 11009 -4285 11043 -4251
rect 11077 -4285 11111 -4251
rect 11461 -4285 11495 -4251
rect 11529 -4285 11563 -4251
rect 11719 -4285 11753 -4251
rect 11787 -4285 11821 -4251
rect 11977 -4285 12011 -4251
rect 12045 -4285 12079 -4251
rect 12429 -4285 12463 -4251
rect 12497 -4285 12531 -4251
rect 12687 -4285 12721 -4251
rect 12755 -4285 12789 -4251
rect 12945 -4285 12979 -4251
rect 13013 -4285 13047 -4251
rect 13203 -4285 13237 -4251
rect 13271 -4285 13305 -4251
rect 13655 -4285 13689 -4251
rect 13723 -4285 13757 -4251
rect 14141 -4285 14175 -4251
rect 14209 -4285 14243 -4251
rect 14592 -4285 14626 -4251
rect 14660 -4285 14694 -4251
rect 14850 -4285 14884 -4251
rect 14918 -4285 14952 -4251
rect 15108 -4285 15142 -4251
rect 15176 -4285 15210 -4251
rect 15366 -4285 15400 -4251
rect 15434 -4285 15468 -4251
rect 15818 -4285 15852 -4251
rect 15886 -4285 15920 -4251
rect 16076 -4285 16110 -4251
rect 16144 -4285 16178 -4251
rect 16334 -4285 16368 -4251
rect 16402 -4285 16436 -4251
rect 16786 -4285 16820 -4251
rect 16854 -4285 16888 -4251
rect 17044 -4285 17078 -4251
rect 17112 -4285 17146 -4251
rect 17302 -4285 17336 -4251
rect 17370 -4285 17404 -4251
rect 17560 -4285 17594 -4251
rect 17628 -4285 17662 -4251
rect 18012 -4285 18046 -4251
rect 18080 -4285 18114 -4251
rect 1066 -4513 1100 -4479
rect 1134 -4513 1168 -4479
rect 1518 -4513 1552 -4479
rect 1586 -4513 1620 -4479
rect 1776 -4513 1810 -4479
rect 1844 -4513 1878 -4479
rect 2034 -4513 2068 -4479
rect 2102 -4513 2136 -4479
rect 2292 -4513 2326 -4479
rect 2360 -4513 2394 -4479
rect 2744 -4513 2778 -4479
rect 2812 -4513 2846 -4479
rect 3002 -4513 3036 -4479
rect 3070 -4513 3104 -4479
rect 3260 -4513 3294 -4479
rect 3328 -4513 3362 -4479
rect 3712 -4513 3746 -4479
rect 3780 -4513 3814 -4479
rect 3970 -4513 4004 -4479
rect 4038 -4513 4072 -4479
rect 4228 -4513 4262 -4479
rect 4296 -4513 4330 -4479
rect 4486 -4513 4520 -4479
rect 4554 -4513 4588 -4479
rect 4937 -4513 4971 -4479
rect 5005 -4513 5039 -4479
rect 5423 -4513 5457 -4479
rect 5491 -4513 5525 -4479
rect 5875 -4513 5909 -4479
rect 5943 -4513 5977 -4479
rect 6133 -4513 6167 -4479
rect 6201 -4513 6235 -4479
rect 6391 -4513 6425 -4479
rect 6459 -4513 6493 -4479
rect 6649 -4513 6683 -4479
rect 6717 -4513 6751 -4479
rect 7101 -4513 7135 -4479
rect 7169 -4513 7203 -4479
rect 7359 -4513 7393 -4479
rect 7427 -4513 7461 -4479
rect 7617 -4513 7651 -4479
rect 7685 -4513 7719 -4479
rect 8069 -4513 8103 -4479
rect 8137 -4513 8171 -4479
rect 8327 -4513 8361 -4479
rect 8395 -4513 8429 -4479
rect 8585 -4513 8619 -4479
rect 8653 -4513 8687 -4479
rect 8843 -4513 8877 -4479
rect 8911 -4513 8945 -4479
rect 9295 -4513 9329 -4479
rect 9363 -4513 9397 -4479
rect 9783 -4513 9817 -4479
rect 9851 -4513 9885 -4479
rect 10235 -4513 10269 -4479
rect 10303 -4513 10337 -4479
rect 10493 -4513 10527 -4479
rect 10561 -4513 10595 -4479
rect 10751 -4513 10785 -4479
rect 10819 -4513 10853 -4479
rect 11009 -4513 11043 -4479
rect 11077 -4513 11111 -4479
rect 11461 -4513 11495 -4479
rect 11529 -4513 11563 -4479
rect 11719 -4513 11753 -4479
rect 11787 -4513 11821 -4479
rect 11977 -4513 12011 -4479
rect 12045 -4513 12079 -4479
rect 12429 -4513 12463 -4479
rect 12497 -4513 12531 -4479
rect 12687 -4513 12721 -4479
rect 12755 -4513 12789 -4479
rect 12945 -4513 12979 -4479
rect 13013 -4513 13047 -4479
rect 13203 -4513 13237 -4479
rect 13271 -4513 13305 -4479
rect 13655 -4513 13689 -4479
rect 13723 -4513 13757 -4479
rect 14141 -4513 14175 -4479
rect 14209 -4513 14243 -4479
rect 14592 -4513 14626 -4479
rect 14660 -4513 14694 -4479
rect 14850 -4513 14884 -4479
rect 14918 -4513 14952 -4479
rect 15108 -4513 15142 -4479
rect 15176 -4513 15210 -4479
rect 15366 -4513 15400 -4479
rect 15434 -4513 15468 -4479
rect 15818 -4513 15852 -4479
rect 15886 -4513 15920 -4479
rect 16076 -4513 16110 -4479
rect 16144 -4513 16178 -4479
rect 16334 -4513 16368 -4479
rect 16402 -4513 16436 -4479
rect 16786 -4513 16820 -4479
rect 16854 -4513 16888 -4479
rect 17044 -4513 17078 -4479
rect 17112 -4513 17146 -4479
rect 17302 -4513 17336 -4479
rect 17370 -4513 17404 -4479
rect 17560 -4513 17594 -4479
rect 17628 -4513 17662 -4479
rect 18012 -4513 18046 -4479
rect 18080 -4513 18114 -4479
rect 1066 -5831 1100 -5797
rect 1134 -5831 1168 -5797
rect 1518 -5831 1552 -5797
rect 1586 -5831 1620 -5797
rect 1776 -5831 1810 -5797
rect 1844 -5831 1878 -5797
rect 2034 -5831 2068 -5797
rect 2102 -5831 2136 -5797
rect 2292 -5831 2326 -5797
rect 2360 -5831 2394 -5797
rect 2744 -5831 2778 -5797
rect 2812 -5831 2846 -5797
rect 3002 -5831 3036 -5797
rect 3070 -5831 3104 -5797
rect 3260 -5831 3294 -5797
rect 3328 -5831 3362 -5797
rect 3712 -5831 3746 -5797
rect 3780 -5831 3814 -5797
rect 3970 -5831 4004 -5797
rect 4038 -5831 4072 -5797
rect 4228 -5831 4262 -5797
rect 4296 -5831 4330 -5797
rect 4486 -5831 4520 -5797
rect 4554 -5831 4588 -5797
rect 4937 -5831 4971 -5797
rect 5005 -5831 5039 -5797
rect 5423 -5831 5457 -5797
rect 5491 -5831 5525 -5797
rect 5875 -5831 5909 -5797
rect 5943 -5831 5977 -5797
rect 6133 -5831 6167 -5797
rect 6201 -5831 6235 -5797
rect 6391 -5831 6425 -5797
rect 6459 -5831 6493 -5797
rect 6649 -5831 6683 -5797
rect 6717 -5831 6751 -5797
rect 7101 -5831 7135 -5797
rect 7169 -5831 7203 -5797
rect 7359 -5831 7393 -5797
rect 7427 -5831 7461 -5797
rect 7617 -5831 7651 -5797
rect 7685 -5831 7719 -5797
rect 8069 -5831 8103 -5797
rect 8137 -5831 8171 -5797
rect 8327 -5831 8361 -5797
rect 8395 -5831 8429 -5797
rect 8585 -5831 8619 -5797
rect 8653 -5831 8687 -5797
rect 8843 -5831 8877 -5797
rect 8911 -5831 8945 -5797
rect 9295 -5831 9329 -5797
rect 9363 -5831 9397 -5797
rect 1066 -6193 1100 -6159
rect 1134 -6193 1168 -6159
rect 1518 -6193 1552 -6159
rect 1586 -6193 1620 -6159
rect 1776 -6193 1810 -6159
rect 1844 -6193 1878 -6159
rect 2034 -6193 2068 -6159
rect 2102 -6193 2136 -6159
rect 2292 -6193 2326 -6159
rect 2360 -6193 2394 -6159
rect 2744 -6193 2778 -6159
rect 2812 -6193 2846 -6159
rect 3002 -6193 3036 -6159
rect 3070 -6193 3104 -6159
rect 3260 -6193 3294 -6159
rect 3328 -6193 3362 -6159
rect 3712 -6193 3746 -6159
rect 3780 -6193 3814 -6159
rect 3970 -6193 4004 -6159
rect 4038 -6193 4072 -6159
rect 4228 -6193 4262 -6159
rect 4296 -6193 4330 -6159
rect 4486 -6193 4520 -6159
rect 4554 -6193 4588 -6159
rect 4937 -6193 4971 -6159
rect 5005 -6193 5039 -6159
rect 9783 -5831 9817 -5797
rect 9851 -5831 9885 -5797
rect 10235 -5831 10269 -5797
rect 10303 -5831 10337 -5797
rect 10493 -5831 10527 -5797
rect 10561 -5831 10595 -5797
rect 10751 -5831 10785 -5797
rect 10819 -5831 10853 -5797
rect 11009 -5831 11043 -5797
rect 11077 -5831 11111 -5797
rect 11461 -5831 11495 -5797
rect 11529 -5831 11563 -5797
rect 11719 -5831 11753 -5797
rect 11787 -5831 11821 -5797
rect 11977 -5831 12011 -5797
rect 12045 -5831 12079 -5797
rect 12429 -5831 12463 -5797
rect 12497 -5831 12531 -5797
rect 12687 -5831 12721 -5797
rect 12755 -5831 12789 -5797
rect 12945 -5831 12979 -5797
rect 13013 -5831 13047 -5797
rect 13203 -5831 13237 -5797
rect 13271 -5831 13305 -5797
rect 13655 -5831 13689 -5797
rect 13723 -5831 13757 -5797
rect 5423 -6193 5457 -6159
rect 5491 -6193 5525 -6159
rect 5875 -6193 5909 -6159
rect 5943 -6193 5977 -6159
rect 6133 -6193 6167 -6159
rect 6201 -6193 6235 -6159
rect 6391 -6193 6425 -6159
rect 6459 -6193 6493 -6159
rect 6649 -6193 6683 -6159
rect 6717 -6193 6751 -6159
rect 7101 -6193 7135 -6159
rect 7169 -6193 7203 -6159
rect 7359 -6193 7393 -6159
rect 7427 -6193 7461 -6159
rect 7617 -6193 7651 -6159
rect 7685 -6193 7719 -6159
rect 8069 -6193 8103 -6159
rect 8137 -6193 8171 -6159
rect 8327 -6193 8361 -6159
rect 8395 -6193 8429 -6159
rect 8585 -6193 8619 -6159
rect 8653 -6193 8687 -6159
rect 8843 -6193 8877 -6159
rect 8911 -6193 8945 -6159
rect 9295 -6193 9329 -6159
rect 9363 -6193 9397 -6159
rect 14141 -5831 14175 -5797
rect 14209 -5831 14243 -5797
rect 14592 -5831 14626 -5797
rect 14660 -5831 14694 -5797
rect 14850 -5831 14884 -5797
rect 14918 -5831 14952 -5797
rect 15108 -5831 15142 -5797
rect 15176 -5831 15210 -5797
rect 15366 -5831 15400 -5797
rect 15434 -5831 15468 -5797
rect 15818 -5831 15852 -5797
rect 15886 -5831 15920 -5797
rect 16076 -5831 16110 -5797
rect 16144 -5831 16178 -5797
rect 16334 -5831 16368 -5797
rect 16402 -5831 16436 -5797
rect 16786 -5831 16820 -5797
rect 16854 -5831 16888 -5797
rect 17044 -5831 17078 -5797
rect 17112 -5831 17146 -5797
rect 17302 -5831 17336 -5797
rect 17370 -5831 17404 -5797
rect 17560 -5831 17594 -5797
rect 17628 -5831 17662 -5797
rect 18012 -5831 18046 -5797
rect 18080 -5831 18114 -5797
rect 9783 -6193 9817 -6159
rect 9851 -6193 9885 -6159
rect 10235 -6193 10269 -6159
rect 10303 -6193 10337 -6159
rect 10493 -6193 10527 -6159
rect 10561 -6193 10595 -6159
rect 10751 -6193 10785 -6159
rect 10819 -6193 10853 -6159
rect 11009 -6193 11043 -6159
rect 11077 -6193 11111 -6159
rect 11461 -6193 11495 -6159
rect 11529 -6193 11563 -6159
rect 11719 -6193 11753 -6159
rect 11787 -6193 11821 -6159
rect 11977 -6193 12011 -6159
rect 12045 -6193 12079 -6159
rect 12429 -6193 12463 -6159
rect 12497 -6193 12531 -6159
rect 12687 -6193 12721 -6159
rect 12755 -6193 12789 -6159
rect 12945 -6193 12979 -6159
rect 13013 -6193 13047 -6159
rect 13203 -6193 13237 -6159
rect 13271 -6193 13305 -6159
rect 13655 -6193 13689 -6159
rect 13723 -6193 13757 -6159
rect 14141 -6193 14175 -6159
rect 14209 -6193 14243 -6159
rect 14592 -6193 14626 -6159
rect 14660 -6193 14694 -6159
rect 14850 -6193 14884 -6159
rect 14918 -6193 14952 -6159
rect 15108 -6193 15142 -6159
rect 15176 -6193 15210 -6159
rect 15366 -6193 15400 -6159
rect 15434 -6193 15468 -6159
rect 15818 -6193 15852 -6159
rect 15886 -6193 15920 -6159
rect 16076 -6193 16110 -6159
rect 16144 -6193 16178 -6159
rect 16334 -6193 16368 -6159
rect 16402 -6193 16436 -6159
rect 16786 -6193 16820 -6159
rect 16854 -6193 16888 -6159
rect 17044 -6193 17078 -6159
rect 17112 -6193 17146 -6159
rect 17302 -6193 17336 -6159
rect 17370 -6193 17404 -6159
rect 17560 -6193 17594 -6159
rect 17628 -6193 17662 -6159
rect 18012 -6193 18046 -6159
rect 18080 -6193 18114 -6159
rect 1066 -7478 1100 -7444
rect 1134 -7478 1168 -7444
rect 1518 -7478 1552 -7444
rect 1586 -7478 1620 -7444
rect 1776 -7478 1810 -7444
rect 1844 -7478 1878 -7444
rect 2034 -7478 2068 -7444
rect 2102 -7478 2136 -7444
rect 2292 -7478 2326 -7444
rect 2360 -7478 2394 -7444
rect 2744 -7478 2778 -7444
rect 2812 -7478 2846 -7444
rect 3002 -7478 3036 -7444
rect 3070 -7478 3104 -7444
rect 3260 -7478 3294 -7444
rect 3328 -7478 3362 -7444
rect 3712 -7478 3746 -7444
rect 3780 -7478 3814 -7444
rect 3970 -7478 4004 -7444
rect 4038 -7478 4072 -7444
rect 4228 -7478 4262 -7444
rect 4296 -7478 4330 -7444
rect 4486 -7478 4520 -7444
rect 4554 -7478 4588 -7444
rect 4937 -7478 4971 -7444
rect 5005 -7478 5039 -7444
rect 5423 -7478 5457 -7444
rect 5491 -7478 5525 -7444
rect 5875 -7478 5909 -7444
rect 5943 -7478 5977 -7444
rect 6133 -7478 6167 -7444
rect 6201 -7478 6235 -7444
rect 6391 -7478 6425 -7444
rect 6459 -7478 6493 -7444
rect 6649 -7478 6683 -7444
rect 6717 -7478 6751 -7444
rect 7101 -7478 7135 -7444
rect 7169 -7478 7203 -7444
rect 7359 -7478 7393 -7444
rect 7427 -7478 7461 -7444
rect 7617 -7478 7651 -7444
rect 7685 -7478 7719 -7444
rect 8069 -7478 8103 -7444
rect 8137 -7478 8171 -7444
rect 8327 -7478 8361 -7444
rect 8395 -7478 8429 -7444
rect 8585 -7478 8619 -7444
rect 8653 -7478 8687 -7444
rect 8843 -7478 8877 -7444
rect 8911 -7478 8945 -7444
rect 9295 -7478 9329 -7444
rect 9363 -7478 9397 -7444
rect 9783 -7478 9817 -7444
rect 9851 -7478 9885 -7444
rect 10235 -7478 10269 -7444
rect 10303 -7478 10337 -7444
rect 10493 -7478 10527 -7444
rect 10561 -7478 10595 -7444
rect 10751 -7478 10785 -7444
rect 10819 -7478 10853 -7444
rect 11009 -7478 11043 -7444
rect 11077 -7478 11111 -7444
rect 11461 -7478 11495 -7444
rect 11529 -7478 11563 -7444
rect 11719 -7478 11753 -7444
rect 11787 -7478 11821 -7444
rect 11977 -7478 12011 -7444
rect 12045 -7478 12079 -7444
rect 12429 -7478 12463 -7444
rect 12497 -7478 12531 -7444
rect 12687 -7478 12721 -7444
rect 12755 -7478 12789 -7444
rect 12945 -7478 12979 -7444
rect 13013 -7478 13047 -7444
rect 13203 -7478 13237 -7444
rect 13271 -7478 13305 -7444
rect 13655 -7478 13689 -7444
rect 13723 -7478 13757 -7444
rect 14141 -7478 14175 -7444
rect 14209 -7478 14243 -7444
rect 14592 -7478 14626 -7444
rect 14660 -7478 14694 -7444
rect 14850 -7478 14884 -7444
rect 14918 -7478 14952 -7444
rect 15108 -7478 15142 -7444
rect 15176 -7478 15210 -7444
rect 15366 -7478 15400 -7444
rect 15434 -7478 15468 -7444
rect 15818 -7478 15852 -7444
rect 15886 -7478 15920 -7444
rect 16076 -7478 16110 -7444
rect 16144 -7478 16178 -7444
rect 16334 -7478 16368 -7444
rect 16402 -7478 16436 -7444
rect 16786 -7478 16820 -7444
rect 16854 -7478 16888 -7444
rect 17044 -7478 17078 -7444
rect 17112 -7478 17146 -7444
rect 17302 -7478 17336 -7444
rect 17370 -7478 17404 -7444
rect 17560 -7478 17594 -7444
rect 17628 -7478 17662 -7444
rect 18012 -7478 18046 -7444
rect 18080 -7478 18114 -7444
rect 1066 -7840 1100 -7806
rect 1134 -7840 1168 -7806
rect 1518 -7840 1552 -7806
rect 1586 -7840 1620 -7806
rect 1776 -7840 1810 -7806
rect 1844 -7840 1878 -7806
rect 2034 -7840 2068 -7806
rect 2102 -7840 2136 -7806
rect 2292 -7840 2326 -7806
rect 2360 -7840 2394 -7806
rect 2744 -7840 2778 -7806
rect 2812 -7840 2846 -7806
rect 3002 -7840 3036 -7806
rect 3070 -7840 3104 -7806
rect 3260 -7840 3294 -7806
rect 3328 -7840 3362 -7806
rect 3712 -7840 3746 -7806
rect 3780 -7840 3814 -7806
rect 3970 -7840 4004 -7806
rect 4038 -7840 4072 -7806
rect 4228 -7840 4262 -7806
rect 4296 -7840 4330 -7806
rect 4486 -7840 4520 -7806
rect 4554 -7840 4588 -7806
rect 4937 -7840 4971 -7806
rect 5005 -7840 5039 -7806
rect 5423 -7840 5457 -7806
rect 5491 -7840 5525 -7806
rect 5875 -7840 5909 -7806
rect 5943 -7840 5977 -7806
rect 6133 -7840 6167 -7806
rect 6201 -7840 6235 -7806
rect 6391 -7840 6425 -7806
rect 6459 -7840 6493 -7806
rect 6649 -7840 6683 -7806
rect 6717 -7840 6751 -7806
rect 7101 -7840 7135 -7806
rect 7169 -7840 7203 -7806
rect 7359 -7840 7393 -7806
rect 7427 -7840 7461 -7806
rect 7617 -7840 7651 -7806
rect 7685 -7840 7719 -7806
rect 8069 -7840 8103 -7806
rect 8137 -7840 8171 -7806
rect 8327 -7840 8361 -7806
rect 8395 -7840 8429 -7806
rect 8585 -7840 8619 -7806
rect 8653 -7840 8687 -7806
rect 8843 -7840 8877 -7806
rect 8911 -7840 8945 -7806
rect 9295 -7840 9329 -7806
rect 9363 -7840 9397 -7806
rect 9783 -7840 9817 -7806
rect 9851 -7840 9885 -7806
rect 10235 -7840 10269 -7806
rect 10303 -7840 10337 -7806
rect 10493 -7840 10527 -7806
rect 10561 -7840 10595 -7806
rect 10751 -7840 10785 -7806
rect 10819 -7840 10853 -7806
rect 11009 -7840 11043 -7806
rect 11077 -7840 11111 -7806
rect 11461 -7840 11495 -7806
rect 11529 -7840 11563 -7806
rect 11719 -7840 11753 -7806
rect 11787 -7840 11821 -7806
rect 11977 -7840 12011 -7806
rect 12045 -7840 12079 -7806
rect 12429 -7840 12463 -7806
rect 12497 -7840 12531 -7806
rect 12687 -7840 12721 -7806
rect 12755 -7840 12789 -7806
rect 12945 -7840 12979 -7806
rect 13013 -7840 13047 -7806
rect 13203 -7840 13237 -7806
rect 13271 -7840 13305 -7806
rect 13655 -7840 13689 -7806
rect 13723 -7840 13757 -7806
rect 14141 -7840 14175 -7806
rect 14209 -7840 14243 -7806
rect 14592 -7840 14626 -7806
rect 14660 -7840 14694 -7806
rect 14850 -7840 14884 -7806
rect 14918 -7840 14952 -7806
rect 15108 -7840 15142 -7806
rect 15176 -7840 15210 -7806
rect 15366 -7840 15400 -7806
rect 15434 -7840 15468 -7806
rect 15818 -7840 15852 -7806
rect 15886 -7840 15920 -7806
rect 16076 -7840 16110 -7806
rect 16144 -7840 16178 -7806
rect 16334 -7840 16368 -7806
rect 16402 -7840 16436 -7806
rect 16786 -7840 16820 -7806
rect 16854 -7840 16888 -7806
rect 17044 -7840 17078 -7806
rect 17112 -7840 17146 -7806
rect 17302 -7840 17336 -7806
rect 17370 -7840 17404 -7806
rect 17560 -7840 17594 -7806
rect 17628 -7840 17662 -7806
rect 18012 -7840 18046 -7806
rect 18080 -7840 18114 -7806
rect 1066 -9112 1100 -9078
rect 1134 -9112 1168 -9078
rect 1518 -9112 1552 -9078
rect 1586 -9112 1620 -9078
rect 1776 -9112 1810 -9078
rect 1844 -9112 1878 -9078
rect 2034 -9112 2068 -9078
rect 2102 -9112 2136 -9078
rect 2292 -9112 2326 -9078
rect 2360 -9112 2394 -9078
rect 2744 -9112 2778 -9078
rect 2812 -9112 2846 -9078
rect 3002 -9112 3036 -9078
rect 3070 -9112 3104 -9078
rect 3260 -9112 3294 -9078
rect 3328 -9112 3362 -9078
rect 3712 -9112 3746 -9078
rect 3780 -9112 3814 -9078
rect 3970 -9112 4004 -9078
rect 4038 -9112 4072 -9078
rect 4228 -9112 4262 -9078
rect 4296 -9112 4330 -9078
rect 4486 -9112 4520 -9078
rect 4554 -9112 4588 -9078
rect 4937 -9112 4971 -9078
rect 5005 -9112 5039 -9078
rect 5423 -9112 5457 -9078
rect 5491 -9112 5525 -9078
rect 5875 -9112 5909 -9078
rect 5943 -9112 5977 -9078
rect 6133 -9112 6167 -9078
rect 6201 -9112 6235 -9078
rect 6391 -9112 6425 -9078
rect 6459 -9112 6493 -9078
rect 6649 -9112 6683 -9078
rect 6717 -9112 6751 -9078
rect 7101 -9112 7135 -9078
rect 7169 -9112 7203 -9078
rect 7359 -9112 7393 -9078
rect 7427 -9112 7461 -9078
rect 7617 -9112 7651 -9078
rect 7685 -9112 7719 -9078
rect 8069 -9112 8103 -9078
rect 8137 -9112 8171 -9078
rect 8327 -9112 8361 -9078
rect 8395 -9112 8429 -9078
rect 8585 -9112 8619 -9078
rect 8653 -9112 8687 -9078
rect 8843 -9112 8877 -9078
rect 8911 -9112 8945 -9078
rect 9295 -9112 9329 -9078
rect 9363 -9112 9397 -9078
rect 9783 -9112 9817 -9078
rect 9851 -9112 9885 -9078
rect 10235 -9112 10269 -9078
rect 10303 -9112 10337 -9078
rect 10493 -9112 10527 -9078
rect 10561 -9112 10595 -9078
rect 10751 -9112 10785 -9078
rect 10819 -9112 10853 -9078
rect 11009 -9112 11043 -9078
rect 11077 -9112 11111 -9078
rect 11461 -9112 11495 -9078
rect 11529 -9112 11563 -9078
rect 11719 -9112 11753 -9078
rect 11787 -9112 11821 -9078
rect 11977 -9112 12011 -9078
rect 12045 -9112 12079 -9078
rect 12429 -9112 12463 -9078
rect 12497 -9112 12531 -9078
rect 12687 -9112 12721 -9078
rect 12755 -9112 12789 -9078
rect 12945 -9112 12979 -9078
rect 13013 -9112 13047 -9078
rect 13203 -9112 13237 -9078
rect 13271 -9112 13305 -9078
rect 13655 -9112 13689 -9078
rect 13723 -9112 13757 -9078
rect 14141 -9112 14175 -9078
rect 14209 -9112 14243 -9078
rect 14592 -9112 14626 -9078
rect 14660 -9112 14694 -9078
rect 14850 -9112 14884 -9078
rect 14918 -9112 14952 -9078
rect 15108 -9112 15142 -9078
rect 15176 -9112 15210 -9078
rect 15366 -9112 15400 -9078
rect 15434 -9112 15468 -9078
rect 15818 -9112 15852 -9078
rect 15886 -9112 15920 -9078
rect 16076 -9112 16110 -9078
rect 16144 -9112 16178 -9078
rect 16334 -9112 16368 -9078
rect 16402 -9112 16436 -9078
rect 16786 -9112 16820 -9078
rect 16854 -9112 16888 -9078
rect 17044 -9112 17078 -9078
rect 17112 -9112 17146 -9078
rect 17302 -9112 17336 -9078
rect 17370 -9112 17404 -9078
rect 17560 -9112 17594 -9078
rect 17628 -9112 17662 -9078
rect 18012 -9112 18046 -9078
rect 18080 -9112 18114 -9078
<< locali >>
rect 856 429 930 463
rect 964 429 977 463
rect 1036 429 1045 463
rect 1108 429 1113 463
rect 1180 429 1181 463
rect 1215 429 1218 463
rect 1283 429 1290 463
rect 1351 429 1362 463
rect 1419 429 1434 463
rect 1487 429 1506 463
rect 1555 429 1578 463
rect 1623 429 1650 463
rect 1691 429 1722 463
rect 1759 429 1793 463
rect 1828 429 1861 463
rect 1900 429 1929 463
rect 1972 429 1997 463
rect 2044 429 2065 463
rect 2116 429 2133 463
rect 2188 429 2201 463
rect 2260 429 2269 463
rect 2332 429 2337 463
rect 2404 429 2405 463
rect 2439 429 2442 463
rect 2507 429 2514 463
rect 2575 429 2586 463
rect 2643 429 2658 463
rect 2711 429 2730 463
rect 2779 429 2802 463
rect 2847 429 2874 463
rect 2915 429 2946 463
rect 2983 429 3017 463
rect 3052 429 3085 463
rect 3124 429 3153 463
rect 3196 429 3221 463
rect 3268 429 3289 463
rect 3340 429 3357 463
rect 3412 429 3425 463
rect 3484 429 3493 463
rect 3556 429 3561 463
rect 3628 429 3629 463
rect 3663 429 3666 463
rect 3731 429 3738 463
rect 3799 429 3810 463
rect 3867 429 3882 463
rect 3935 429 3954 463
rect 4003 429 4026 463
rect 4071 429 4098 463
rect 4139 429 4170 463
rect 4207 429 4241 463
rect 4276 429 4309 463
rect 4348 429 4377 463
rect 4420 429 4445 463
rect 4492 429 4513 463
rect 4564 429 4581 463
rect 4636 429 4649 463
rect 4708 429 4717 463
rect 4780 429 4785 463
rect 4852 429 4853 463
rect 4887 429 4890 463
rect 4955 429 4962 463
rect 5023 429 5034 463
rect 5091 429 5106 463
rect 5140 429 5323 463
rect 5357 429 5372 463
rect 5429 429 5440 463
rect 5501 429 5508 463
rect 5573 429 5576 463
rect 5610 429 5611 463
rect 5678 429 5683 463
rect 5746 429 5755 463
rect 5814 429 5827 463
rect 5882 429 5899 463
rect 5950 429 5971 463
rect 6018 429 6043 463
rect 6086 429 6115 463
rect 6154 429 6187 463
rect 6222 429 6256 463
rect 6293 429 6324 463
rect 6365 429 6392 463
rect 6437 429 6460 463
rect 6509 429 6528 463
rect 6581 429 6596 463
rect 6653 429 6664 463
rect 6725 429 6732 463
rect 6797 429 6800 463
rect 6834 429 6835 463
rect 6902 429 6907 463
rect 6970 429 6979 463
rect 7038 429 7051 463
rect 7106 429 7123 463
rect 7174 429 7195 463
rect 7242 429 7267 463
rect 7310 429 7339 463
rect 7378 429 7411 463
rect 7446 429 7480 463
rect 7517 429 7548 463
rect 7589 429 7616 463
rect 7661 429 7684 463
rect 7733 429 7752 463
rect 7805 429 7820 463
rect 7877 429 7888 463
rect 7949 429 7956 463
rect 8021 429 8024 463
rect 8058 429 8059 463
rect 8126 429 8131 463
rect 8194 429 8203 463
rect 8262 429 8275 463
rect 8330 429 8347 463
rect 8398 429 8419 463
rect 8466 429 8491 463
rect 8534 429 8563 463
rect 8602 429 8635 463
rect 8670 429 8704 463
rect 8741 429 8772 463
rect 8813 429 8840 463
rect 8885 429 8908 463
rect 8957 429 8976 463
rect 9029 429 9044 463
rect 9101 429 9112 463
rect 9173 429 9180 463
rect 9245 429 9248 463
rect 9282 429 9283 463
rect 9350 429 9355 463
rect 9418 429 9427 463
rect 9486 429 9499 463
rect 9533 429 9647 463
rect 9681 429 9694 463
rect 9753 429 9762 463
rect 9825 429 9830 463
rect 9897 429 9898 463
rect 9932 429 9935 463
rect 10000 429 10007 463
rect 10068 429 10079 463
rect 10136 429 10151 463
rect 10204 429 10223 463
rect 10272 429 10295 463
rect 10340 429 10367 463
rect 10408 429 10439 463
rect 10476 429 10510 463
rect 10545 429 10578 463
rect 10617 429 10646 463
rect 10689 429 10714 463
rect 10761 429 10782 463
rect 10833 429 10850 463
rect 10905 429 10918 463
rect 10977 429 10986 463
rect 11049 429 11054 463
rect 11121 429 11122 463
rect 11156 429 11159 463
rect 11224 429 11231 463
rect 11292 429 11303 463
rect 11360 429 11375 463
rect 11428 429 11447 463
rect 11496 429 11519 463
rect 11564 429 11591 463
rect 11632 429 11663 463
rect 11700 429 11734 463
rect 11769 429 11802 463
rect 11841 429 11870 463
rect 11913 429 11938 463
rect 11985 429 12006 463
rect 12057 429 12074 463
rect 12129 429 12142 463
rect 12201 429 12210 463
rect 12273 429 12278 463
rect 12345 429 12346 463
rect 12380 429 12383 463
rect 12448 429 12455 463
rect 12516 429 12527 463
rect 12584 429 12599 463
rect 12652 429 12671 463
rect 12720 429 12743 463
rect 12788 429 12815 463
rect 12856 429 12887 463
rect 12924 429 12958 463
rect 12993 429 13026 463
rect 13065 429 13094 463
rect 13137 429 13162 463
rect 13209 429 13230 463
rect 13281 429 13298 463
rect 13353 429 13366 463
rect 13425 429 13434 463
rect 13497 429 13502 463
rect 13569 429 13570 463
rect 13604 429 13607 463
rect 13672 429 13679 463
rect 13740 429 13751 463
rect 13808 429 13823 463
rect 13857 429 14040 463
rect 14074 429 14089 463
rect 14146 429 14157 463
rect 14218 429 14225 463
rect 14290 429 14293 463
rect 14327 429 14328 463
rect 14395 429 14400 463
rect 14463 429 14472 463
rect 14531 429 14544 463
rect 14599 429 14616 463
rect 14667 429 14688 463
rect 14735 429 14760 463
rect 14803 429 14832 463
rect 14871 429 14904 463
rect 14939 429 14973 463
rect 15010 429 15041 463
rect 15082 429 15109 463
rect 15154 429 15177 463
rect 15226 429 15245 463
rect 15298 429 15313 463
rect 15370 429 15381 463
rect 15442 429 15449 463
rect 15514 429 15517 463
rect 15551 429 15552 463
rect 15619 429 15624 463
rect 15687 429 15696 463
rect 15755 429 15768 463
rect 15823 429 15840 463
rect 15891 429 15912 463
rect 15959 429 15984 463
rect 16027 429 16056 463
rect 16095 429 16128 463
rect 16163 429 16197 463
rect 16234 429 16265 463
rect 16306 429 16333 463
rect 16378 429 16401 463
rect 16450 429 16469 463
rect 16522 429 16537 463
rect 16594 429 16605 463
rect 16666 429 16673 463
rect 16738 429 16741 463
rect 16775 429 16776 463
rect 16843 429 16848 463
rect 16911 429 16920 463
rect 16979 429 16992 463
rect 17047 429 17064 463
rect 17115 429 17136 463
rect 17183 429 17208 463
rect 17251 429 17280 463
rect 17319 429 17352 463
rect 17387 429 17421 463
rect 17458 429 17489 463
rect 17530 429 17557 463
rect 17602 429 17625 463
rect 17674 429 17693 463
rect 17746 429 17761 463
rect 17818 429 17829 463
rect 17890 429 17897 463
rect 17962 429 17965 463
rect 17999 429 18000 463
rect 18067 429 18072 463
rect 18135 429 18144 463
rect 18203 429 18216 463
rect 18250 429 18324 463
rect 856 306 890 429
rect 1017 315 1064 349
rect 1100 315 1134 349
rect 1170 315 1217 349
rect 1469 315 1516 349
rect 1552 315 1586 349
rect 1622 315 1669 349
rect 1727 315 1774 349
rect 1810 315 1844 349
rect 1880 315 1927 349
rect 1985 315 2032 349
rect 2068 315 2102 349
rect 2138 315 2185 349
rect 2243 315 2290 349
rect 2326 315 2360 349
rect 2396 315 2443 349
rect 2695 315 2742 349
rect 2778 315 2812 349
rect 2848 315 2895 349
rect 2953 315 3000 349
rect 3036 315 3070 349
rect 3106 315 3153 349
rect 3211 315 3258 349
rect 3294 315 3328 349
rect 3364 315 3411 349
rect 3663 315 3710 349
rect 3746 315 3780 349
rect 3816 315 3863 349
rect 3921 315 3968 349
rect 4004 315 4038 349
rect 4074 315 4121 349
rect 4179 315 4226 349
rect 4262 315 4296 349
rect 4332 315 4379 349
rect 4437 315 4484 349
rect 4520 315 4554 349
rect 4590 315 4637 349
rect 4888 315 4935 349
rect 4971 315 5005 349
rect 5041 315 5088 349
rect 5214 306 5249 429
rect 5374 315 5421 349
rect 5457 315 5491 349
rect 5527 315 5574 349
rect 5826 315 5873 349
rect 5909 315 5943 349
rect 5979 315 6026 349
rect 6084 315 6131 349
rect 6167 315 6201 349
rect 6237 315 6284 349
rect 6342 315 6389 349
rect 6425 315 6459 349
rect 6495 315 6542 349
rect 6600 315 6647 349
rect 6683 315 6717 349
rect 6753 315 6800 349
rect 7052 315 7099 349
rect 7135 315 7169 349
rect 7205 315 7252 349
rect 7310 315 7357 349
rect 7393 315 7427 349
rect 7463 315 7510 349
rect 7568 315 7615 349
rect 7651 315 7685 349
rect 7721 315 7768 349
rect 8020 315 8067 349
rect 8103 315 8137 349
rect 8173 315 8220 349
rect 8278 315 8325 349
rect 8361 315 8395 349
rect 8431 315 8478 349
rect 8536 315 8583 349
rect 8619 315 8653 349
rect 8689 315 8736 349
rect 8794 315 8841 349
rect 8877 315 8911 349
rect 8947 315 8994 349
rect 9246 315 9293 349
rect 9329 315 9363 349
rect 9399 315 9446 349
rect 5248 272 5249 306
rect 9573 306 9607 429
rect 9734 315 9781 349
rect 9817 315 9851 349
rect 9887 315 9934 349
rect 10186 315 10233 349
rect 10269 315 10303 349
rect 10339 315 10386 349
rect 10444 315 10491 349
rect 10527 315 10561 349
rect 10597 315 10644 349
rect 10702 315 10749 349
rect 10785 315 10819 349
rect 10855 315 10902 349
rect 10960 315 11007 349
rect 11043 315 11077 349
rect 11113 315 11160 349
rect 11412 315 11459 349
rect 11495 315 11529 349
rect 11565 315 11612 349
rect 11670 315 11717 349
rect 11753 315 11787 349
rect 11823 315 11870 349
rect 11928 315 11975 349
rect 12011 315 12045 349
rect 12081 315 12128 349
rect 12380 315 12427 349
rect 12463 315 12497 349
rect 12533 315 12580 349
rect 12638 315 12685 349
rect 12721 315 12755 349
rect 12791 315 12838 349
rect 12896 315 12943 349
rect 12979 315 13013 349
rect 13049 315 13096 349
rect 13154 315 13201 349
rect 13237 315 13271 349
rect 13307 315 13354 349
rect 13606 315 13653 349
rect 13689 315 13723 349
rect 13759 315 13806 349
rect 13931 306 13966 429
rect 14092 315 14139 349
rect 14175 315 14209 349
rect 14245 315 14292 349
rect 14543 315 14590 349
rect 14626 315 14660 349
rect 14696 315 14743 349
rect 14801 315 14848 349
rect 14884 315 14918 349
rect 14954 315 15001 349
rect 15059 315 15106 349
rect 15142 315 15176 349
rect 15212 315 15259 349
rect 15317 315 15364 349
rect 15400 315 15434 349
rect 15470 315 15517 349
rect 15769 315 15816 349
rect 15852 315 15886 349
rect 15922 315 15969 349
rect 16027 315 16074 349
rect 16110 315 16144 349
rect 16180 315 16227 349
rect 16285 315 16332 349
rect 16368 315 16402 349
rect 16438 315 16485 349
rect 16737 315 16784 349
rect 16820 315 16854 349
rect 16890 315 16937 349
rect 16995 315 17042 349
rect 17078 315 17112 349
rect 17148 315 17195 349
rect 17253 315 17300 349
rect 17336 315 17370 349
rect 17406 315 17453 349
rect 17511 315 17558 349
rect 17594 315 17628 349
rect 17664 315 17711 349
rect 17963 315 18010 349
rect 18046 315 18080 349
rect 18116 315 18163 349
rect 13931 272 13932 306
rect 18290 306 18324 429
rect 856 250 890 272
rect 856 182 890 200
rect 856 114 890 128
rect 971 253 1005 272
rect 971 185 1005 187
rect 971 149 1005 151
rect 971 64 1005 83
rect 1229 253 1263 272
rect 1229 185 1263 187
rect 1229 149 1263 151
rect 1229 64 1263 83
rect 1423 253 1457 272
rect 1423 185 1457 187
rect 1423 149 1457 151
rect 1423 64 1457 83
rect 1681 253 1715 272
rect 1681 185 1715 187
rect 1681 149 1715 151
rect 1681 64 1715 83
rect 1939 253 1973 272
rect 1939 185 1973 187
rect 1939 149 1973 151
rect 1939 64 1973 83
rect 2197 253 2231 272
rect 2197 185 2231 187
rect 2197 149 2231 151
rect 2197 64 2231 83
rect 2455 253 2489 272
rect 2455 185 2489 187
rect 2455 149 2489 151
rect 2455 64 2489 83
rect 2649 253 2683 272
rect 2649 185 2683 187
rect 2649 149 2683 151
rect 2649 64 2683 83
rect 2907 253 2941 272
rect 2907 185 2941 187
rect 2907 149 2941 151
rect 2907 64 2941 83
rect 3165 253 3199 272
rect 3165 185 3199 187
rect 3165 149 3199 151
rect 3165 64 3199 83
rect 3423 253 3457 272
rect 3423 185 3457 187
rect 3423 149 3457 151
rect 3423 64 3457 83
rect 3617 253 3651 272
rect 3617 185 3651 187
rect 3617 149 3651 151
rect 3617 64 3651 83
rect 3875 253 3909 272
rect 3875 185 3909 187
rect 3875 149 3909 151
rect 3875 64 3909 83
rect 4133 253 4167 272
rect 4133 185 4167 187
rect 4133 149 4167 151
rect 4133 64 4167 83
rect 4391 253 4425 272
rect 4391 185 4425 187
rect 4391 149 4425 151
rect 4391 64 4425 83
rect 4649 253 4683 272
rect 4649 185 4683 187
rect 4649 149 4683 151
rect 4649 64 4683 83
rect 4842 253 4876 272
rect 4842 185 4876 187
rect 4842 149 4876 151
rect 4842 64 4876 83
rect 5100 253 5134 272
rect 5100 185 5134 187
rect 5100 149 5134 151
rect 5100 64 5134 83
rect 5214 250 5249 272
rect 5248 200 5249 250
rect 5214 182 5249 200
rect 5248 128 5249 182
rect 5214 114 5249 128
rect 856 46 890 56
rect 856 -22 890 -16
rect 856 -90 890 -88
rect 856 -126 890 -124
rect 856 -198 890 -192
rect 856 -270 890 -260
rect 5248 56 5249 114
rect 5328 253 5362 272
rect 5328 185 5362 187
rect 5328 149 5362 151
rect 5328 64 5362 83
rect 5586 253 5620 272
rect 5586 185 5620 187
rect 5586 149 5620 151
rect 5586 64 5620 83
rect 5780 253 5814 272
rect 5780 185 5814 187
rect 5780 149 5814 151
rect 5780 64 5814 83
rect 6038 253 6072 272
rect 6038 185 6072 187
rect 6038 149 6072 151
rect 6038 64 6072 83
rect 6296 253 6330 272
rect 6296 185 6330 187
rect 6296 149 6330 151
rect 6296 64 6330 83
rect 6554 253 6588 272
rect 6554 185 6588 187
rect 6554 149 6588 151
rect 6554 64 6588 83
rect 6812 253 6846 272
rect 6812 185 6846 187
rect 6812 149 6846 151
rect 6812 64 6846 83
rect 7006 253 7040 272
rect 7006 185 7040 187
rect 7006 149 7040 151
rect 7006 64 7040 83
rect 7264 253 7298 272
rect 7264 185 7298 187
rect 7264 149 7298 151
rect 7264 64 7298 83
rect 7522 253 7556 272
rect 7522 185 7556 187
rect 7522 149 7556 151
rect 7522 64 7556 83
rect 7780 253 7814 272
rect 7780 185 7814 187
rect 7780 149 7814 151
rect 7780 64 7814 83
rect 7974 253 8008 272
rect 7974 185 8008 187
rect 7974 149 8008 151
rect 7974 64 8008 83
rect 8232 253 8266 272
rect 8232 185 8266 187
rect 8232 149 8266 151
rect 8232 64 8266 83
rect 8490 253 8524 272
rect 8490 185 8524 187
rect 8490 149 8524 151
rect 8490 64 8524 83
rect 8748 253 8782 272
rect 8748 185 8782 187
rect 8748 149 8782 151
rect 8748 64 8782 83
rect 9006 253 9040 272
rect 9006 185 9040 187
rect 9006 149 9040 151
rect 9006 64 9040 83
rect 9200 253 9234 272
rect 9200 185 9234 187
rect 9200 149 9234 151
rect 9200 64 9234 83
rect 9458 253 9492 272
rect 9458 185 9492 187
rect 9458 149 9492 151
rect 9458 64 9492 83
rect 9573 250 9607 272
rect 9573 182 9607 200
rect 9573 114 9607 128
rect 5214 46 5249 56
rect 5248 -16 5249 46
rect 5214 -22 5249 -16
rect 5248 -88 5249 -22
rect 5214 -90 5249 -88
rect 5248 -124 5249 -90
rect 5214 -126 5249 -124
rect 5248 -192 5249 -126
rect 5214 -198 5249 -192
rect 5248 -260 5249 -198
rect 5214 -270 5249 -260
rect 5248 -328 5249 -270
rect 9688 253 9722 272
rect 9688 185 9722 187
rect 9688 149 9722 151
rect 9688 64 9722 83
rect 9946 253 9980 272
rect 9946 185 9980 187
rect 9946 149 9980 151
rect 9946 64 9980 83
rect 10140 253 10174 272
rect 10140 185 10174 187
rect 10140 149 10174 151
rect 10140 64 10174 83
rect 10398 253 10432 272
rect 10398 185 10432 187
rect 10398 149 10432 151
rect 10398 64 10432 83
rect 10656 253 10690 272
rect 10656 185 10690 187
rect 10656 149 10690 151
rect 10656 64 10690 83
rect 10914 253 10948 272
rect 10914 185 10948 187
rect 10914 149 10948 151
rect 10914 64 10948 83
rect 11172 253 11206 272
rect 11172 185 11206 187
rect 11172 149 11206 151
rect 11172 64 11206 83
rect 11366 253 11400 272
rect 11366 185 11400 187
rect 11366 149 11400 151
rect 11366 64 11400 83
rect 11624 253 11658 272
rect 11624 185 11658 187
rect 11624 149 11658 151
rect 11624 64 11658 83
rect 11882 253 11916 272
rect 11882 185 11916 187
rect 11882 149 11916 151
rect 11882 64 11916 83
rect 12140 253 12174 272
rect 12140 185 12174 187
rect 12140 149 12174 151
rect 12140 64 12174 83
rect 12334 253 12368 272
rect 12334 185 12368 187
rect 12334 149 12368 151
rect 12334 64 12368 83
rect 12592 253 12626 272
rect 12592 185 12626 187
rect 12592 149 12626 151
rect 12592 64 12626 83
rect 12850 253 12884 272
rect 12850 185 12884 187
rect 12850 149 12884 151
rect 12850 64 12884 83
rect 13108 253 13142 272
rect 13108 185 13142 187
rect 13108 149 13142 151
rect 13108 64 13142 83
rect 13366 253 13400 272
rect 13366 185 13400 187
rect 13366 149 13400 151
rect 13366 64 13400 83
rect 13560 253 13594 272
rect 13560 185 13594 187
rect 13560 149 13594 151
rect 13560 64 13594 83
rect 13818 253 13852 272
rect 13818 185 13852 187
rect 13818 149 13852 151
rect 13818 64 13852 83
rect 13931 250 13966 272
rect 13931 200 13932 250
rect 13931 182 13966 200
rect 13931 128 13932 182
rect 13931 114 13966 128
rect 9573 46 9607 56
rect 9573 -22 9607 -16
rect 9573 -90 9607 -88
rect 9573 -126 9607 -124
rect 9573 -198 9607 -192
rect 9573 -270 9607 -260
rect 13931 56 13932 114
rect 14046 253 14080 272
rect 14046 185 14080 187
rect 14046 149 14080 151
rect 14046 64 14080 83
rect 14304 253 14338 272
rect 14304 185 14338 187
rect 14304 149 14338 151
rect 14304 64 14338 83
rect 14497 253 14531 272
rect 14497 185 14531 187
rect 14497 149 14531 151
rect 14497 64 14531 83
rect 14755 253 14789 272
rect 14755 185 14789 187
rect 14755 149 14789 151
rect 14755 64 14789 83
rect 15013 253 15047 272
rect 15013 185 15047 187
rect 15013 149 15047 151
rect 15013 64 15047 83
rect 15271 253 15305 272
rect 15271 185 15305 187
rect 15271 149 15305 151
rect 15271 64 15305 83
rect 15529 253 15563 272
rect 15529 185 15563 187
rect 15529 149 15563 151
rect 15529 64 15563 83
rect 15723 253 15757 272
rect 15723 185 15757 187
rect 15723 149 15757 151
rect 15723 64 15757 83
rect 15981 253 16015 272
rect 15981 185 16015 187
rect 15981 149 16015 151
rect 15981 64 16015 83
rect 16239 253 16273 272
rect 16239 185 16273 187
rect 16239 149 16273 151
rect 16239 64 16273 83
rect 16497 253 16531 272
rect 16497 185 16531 187
rect 16497 149 16531 151
rect 16497 64 16531 83
rect 16691 253 16725 272
rect 16691 185 16725 187
rect 16691 149 16725 151
rect 16691 64 16725 83
rect 16949 253 16983 272
rect 16949 185 16983 187
rect 16949 149 16983 151
rect 16949 64 16983 83
rect 17207 253 17241 272
rect 17207 185 17241 187
rect 17207 149 17241 151
rect 17207 64 17241 83
rect 17465 253 17499 272
rect 17465 185 17499 187
rect 17465 149 17499 151
rect 17465 64 17499 83
rect 17723 253 17757 272
rect 17723 185 17757 187
rect 17723 149 17757 151
rect 17723 64 17757 83
rect 17917 253 17951 272
rect 17917 185 17951 187
rect 17917 149 17951 151
rect 17917 64 17951 83
rect 18175 253 18209 272
rect 18175 185 18209 187
rect 18175 149 18209 151
rect 18175 64 18209 83
rect 18290 250 18324 272
rect 18290 182 18324 200
rect 18290 114 18324 128
rect 13931 46 13966 56
rect 13931 -16 13932 46
rect 13931 -22 13966 -16
rect 13931 -88 13932 -22
rect 13931 -90 13966 -88
rect 13931 -124 13932 -90
rect 13931 -126 13966 -124
rect 13931 -192 13932 -126
rect 13931 -198 13966 -192
rect 13931 -260 13932 -198
rect 13931 -270 13966 -260
rect 13931 -328 13932 -270
rect 18290 46 18324 56
rect 18290 -22 18324 -16
rect 18290 -90 18324 -88
rect 18290 -126 18324 -124
rect 18290 -198 18324 -192
rect 18290 -270 18324 -260
rect 856 -342 977 -328
rect 890 -362 977 -342
rect 1011 -362 1045 -328
rect 1079 -362 1113 -328
rect 1147 -362 1181 -328
rect 1215 -362 1249 -328
rect 1283 -362 1317 -328
rect 1351 -362 1385 -328
rect 1419 -362 1453 -328
rect 1487 -362 1521 -328
rect 1555 -362 1589 -328
rect 1623 -362 1657 -328
rect 1691 -362 1725 -328
rect 1759 -362 1793 -328
rect 1827 -362 1861 -328
rect 1895 -362 1929 -328
rect 1963 -362 1997 -328
rect 2031 -362 2065 -328
rect 2099 -362 2133 -328
rect 2167 -362 2201 -328
rect 2235 -362 2269 -328
rect 2303 -362 2337 -328
rect 2371 -362 2405 -328
rect 2439 -362 2473 -328
rect 2507 -362 2541 -328
rect 2575 -362 2609 -328
rect 2643 -362 2677 -328
rect 2711 -362 2745 -328
rect 2779 -362 2813 -328
rect 2847 -362 2881 -328
rect 2915 -362 2949 -328
rect 2983 -362 3017 -328
rect 3051 -362 3085 -328
rect 3119 -362 3153 -328
rect 3187 -362 3221 -328
rect 3255 -362 3289 -328
rect 3323 -362 3357 -328
rect 3391 -362 3425 -328
rect 3459 -362 3493 -328
rect 3527 -362 3561 -328
rect 3595 -362 3629 -328
rect 3663 -362 3697 -328
rect 3731 -362 3765 -328
rect 3799 -362 3833 -328
rect 3867 -362 3901 -328
rect 3935 -362 3969 -328
rect 4003 -362 4037 -328
rect 4071 -362 4105 -328
rect 4139 -362 4173 -328
rect 4207 -362 4241 -328
rect 4275 -362 4309 -328
rect 4343 -362 4377 -328
rect 4411 -362 4445 -328
rect 4479 -362 4513 -328
rect 4547 -362 4581 -328
rect 4615 -362 4649 -328
rect 4683 -362 4717 -328
rect 4751 -362 4785 -328
rect 4819 -362 4853 -328
rect 4887 -362 4921 -328
rect 4955 -362 4989 -328
rect 5023 -362 5057 -328
rect 5091 -342 5372 -328
rect 5091 -362 5214 -342
rect 5248 -362 5372 -342
rect 5406 -362 5440 -328
rect 5474 -362 5508 -328
rect 5542 -362 5576 -328
rect 5610 -362 5644 -328
rect 5678 -362 5712 -328
rect 5746 -362 5780 -328
rect 5814 -362 5848 -328
rect 5882 -362 5916 -328
rect 5950 -362 5984 -328
rect 6018 -362 6052 -328
rect 6086 -362 6120 -328
rect 6154 -362 6188 -328
rect 6222 -362 6256 -328
rect 6290 -362 6324 -328
rect 6358 -362 6392 -328
rect 6426 -362 6460 -328
rect 6494 -362 6528 -328
rect 6562 -362 6596 -328
rect 6630 -362 6664 -328
rect 6698 -362 6732 -328
rect 6766 -362 6800 -328
rect 6834 -362 6868 -328
rect 6902 -362 6936 -328
rect 6970 -362 7004 -328
rect 7038 -362 7072 -328
rect 7106 -362 7140 -328
rect 7174 -362 7208 -328
rect 7242 -362 7276 -328
rect 7310 -362 7344 -328
rect 7378 -362 7412 -328
rect 7446 -362 7480 -328
rect 7514 -362 7548 -328
rect 7582 -362 7616 -328
rect 7650 -362 7684 -328
rect 7718 -362 7752 -328
rect 7786 -362 7820 -328
rect 7854 -362 7888 -328
rect 7922 -362 7956 -328
rect 7990 -362 8024 -328
rect 8058 -362 8092 -328
rect 8126 -362 8160 -328
rect 8194 -362 8228 -328
rect 8262 -362 8296 -328
rect 8330 -362 8364 -328
rect 8398 -362 8432 -328
rect 8466 -362 8500 -328
rect 8534 -362 8568 -328
rect 8602 -362 8636 -328
rect 8670 -362 8704 -328
rect 8738 -362 8772 -328
rect 8806 -362 8840 -328
rect 8874 -362 8908 -328
rect 8942 -362 8976 -328
rect 9010 -362 9044 -328
rect 9078 -362 9112 -328
rect 9146 -362 9180 -328
rect 9214 -362 9248 -328
rect 9282 -362 9316 -328
rect 9350 -362 9384 -328
rect 9418 -362 9452 -328
rect 9486 -342 9694 -328
rect 9486 -362 9573 -342
rect 9607 -362 9694 -342
rect 9728 -362 9762 -328
rect 9796 -362 9830 -328
rect 9864 -362 9898 -328
rect 9932 -362 9966 -328
rect 10000 -362 10034 -328
rect 10068 -362 10102 -328
rect 10136 -362 10170 -328
rect 10204 -362 10238 -328
rect 10272 -362 10306 -328
rect 10340 -362 10374 -328
rect 10408 -362 10442 -328
rect 10476 -362 10510 -328
rect 10544 -362 10578 -328
rect 10612 -362 10646 -328
rect 10680 -362 10714 -328
rect 10748 -362 10782 -328
rect 10816 -362 10850 -328
rect 10884 -362 10918 -328
rect 10952 -362 10986 -328
rect 11020 -362 11054 -328
rect 11088 -362 11122 -328
rect 11156 -362 11190 -328
rect 11224 -362 11258 -328
rect 11292 -362 11326 -328
rect 11360 -362 11394 -328
rect 11428 -362 11462 -328
rect 11496 -362 11530 -328
rect 11564 -362 11598 -328
rect 11632 -362 11666 -328
rect 11700 -362 11734 -328
rect 11768 -362 11802 -328
rect 11836 -362 11870 -328
rect 11904 -362 11938 -328
rect 11972 -362 12006 -328
rect 12040 -362 12074 -328
rect 12108 -362 12142 -328
rect 12176 -362 12210 -328
rect 12244 -362 12278 -328
rect 12312 -362 12346 -328
rect 12380 -362 12414 -328
rect 12448 -362 12482 -328
rect 12516 -362 12550 -328
rect 12584 -362 12618 -328
rect 12652 -362 12686 -328
rect 12720 -362 12754 -328
rect 12788 -362 12822 -328
rect 12856 -362 12890 -328
rect 12924 -362 12958 -328
rect 12992 -362 13026 -328
rect 13060 -362 13094 -328
rect 13128 -362 13162 -328
rect 13196 -362 13230 -328
rect 13264 -362 13298 -328
rect 13332 -362 13366 -328
rect 13400 -362 13434 -328
rect 13468 -362 13502 -328
rect 13536 -362 13570 -328
rect 13604 -362 13638 -328
rect 13672 -362 13706 -328
rect 13740 -362 13774 -328
rect 13808 -342 14089 -328
rect 13808 -362 13932 -342
rect 13966 -362 14089 -342
rect 14123 -362 14157 -328
rect 14191 -362 14225 -328
rect 14259 -362 14293 -328
rect 14327 -362 14361 -328
rect 14395 -362 14429 -328
rect 14463 -362 14497 -328
rect 14531 -362 14565 -328
rect 14599 -362 14633 -328
rect 14667 -362 14701 -328
rect 14735 -362 14769 -328
rect 14803 -362 14837 -328
rect 14871 -362 14905 -328
rect 14939 -362 14973 -328
rect 15007 -362 15041 -328
rect 15075 -362 15109 -328
rect 15143 -362 15177 -328
rect 15211 -362 15245 -328
rect 15279 -362 15313 -328
rect 15347 -362 15381 -328
rect 15415 -362 15449 -328
rect 15483 -362 15517 -328
rect 15551 -362 15585 -328
rect 15619 -362 15653 -328
rect 15687 -362 15721 -328
rect 15755 -362 15789 -328
rect 15823 -362 15857 -328
rect 15891 -362 15925 -328
rect 15959 -362 15993 -328
rect 16027 -362 16061 -328
rect 16095 -362 16129 -328
rect 16163 -362 16197 -328
rect 16231 -362 16265 -328
rect 16299 -362 16333 -328
rect 16367 -362 16401 -328
rect 16435 -362 16469 -328
rect 16503 -362 16537 -328
rect 16571 -362 16605 -328
rect 16639 -362 16673 -328
rect 16707 -362 16741 -328
rect 16775 -362 16809 -328
rect 16843 -362 16877 -328
rect 16911 -362 16945 -328
rect 16979 -362 17013 -328
rect 17047 -362 17081 -328
rect 17115 -362 17149 -328
rect 17183 -362 17217 -328
rect 17251 -362 17285 -328
rect 17319 -362 17353 -328
rect 17387 -362 17421 -328
rect 17455 -362 17489 -328
rect 17523 -362 17557 -328
rect 17591 -362 17625 -328
rect 17659 -362 17693 -328
rect 17727 -362 17761 -328
rect 17795 -362 17829 -328
rect 17863 -362 17897 -328
rect 17931 -362 17965 -328
rect 17999 -362 18033 -328
rect 18067 -362 18101 -328
rect 18135 -362 18169 -328
rect 18203 -342 18324 -328
rect 18203 -362 18290 -342
rect 856 -414 890 -396
rect 856 -486 890 -464
rect 856 -558 890 -532
rect 856 -630 890 -600
rect 856 -702 890 -668
rect 5248 -396 5249 -362
rect 5214 -414 5249 -396
rect 5248 -464 5249 -414
rect 5214 -486 5249 -464
rect 5248 -532 5249 -486
rect 5214 -558 5249 -532
rect 5248 -600 5249 -558
rect 5214 -630 5249 -600
rect 5248 -668 5249 -630
rect 856 -770 890 -736
rect 856 -838 890 -808
rect 971 -691 1005 -672
rect 971 -759 1005 -757
rect 971 -795 1005 -793
rect 971 -880 1005 -861
rect 1229 -691 1263 -672
rect 1229 -759 1263 -757
rect 1229 -795 1263 -793
rect 1229 -880 1263 -861
rect 1423 -691 1457 -672
rect 1423 -759 1457 -757
rect 1423 -795 1457 -793
rect 1423 -880 1457 -861
rect 1681 -691 1715 -672
rect 1681 -759 1715 -757
rect 1681 -795 1715 -793
rect 1681 -880 1715 -861
rect 1939 -691 1973 -672
rect 1939 -759 1973 -757
rect 1939 -795 1973 -793
rect 1939 -880 1973 -861
rect 2197 -691 2231 -672
rect 2197 -759 2231 -757
rect 2197 -795 2231 -793
rect 2197 -880 2231 -861
rect 2455 -691 2489 -672
rect 2455 -759 2489 -757
rect 2455 -795 2489 -793
rect 2455 -880 2489 -861
rect 2649 -691 2683 -672
rect 2649 -759 2683 -757
rect 2649 -795 2683 -793
rect 2649 -880 2683 -861
rect 2907 -691 2941 -672
rect 2907 -759 2941 -757
rect 2907 -795 2941 -793
rect 2907 -880 2941 -861
rect 3165 -691 3199 -672
rect 3165 -759 3199 -757
rect 3165 -795 3199 -793
rect 3165 -880 3199 -861
rect 3423 -691 3457 -672
rect 3423 -759 3457 -757
rect 3423 -795 3457 -793
rect 3423 -880 3457 -861
rect 3617 -691 3651 -672
rect 3617 -759 3651 -757
rect 3617 -795 3651 -793
rect 3617 -880 3651 -861
rect 3875 -691 3909 -672
rect 3875 -759 3909 -757
rect 3875 -795 3909 -793
rect 3875 -880 3909 -861
rect 4133 -691 4167 -672
rect 4133 -759 4167 -757
rect 4133 -795 4167 -793
rect 4133 -880 4167 -861
rect 4391 -691 4425 -672
rect 4391 -759 4425 -757
rect 4391 -795 4425 -793
rect 4391 -880 4425 -861
rect 4649 -691 4683 -672
rect 4649 -759 4683 -757
rect 4649 -795 4683 -793
rect 4649 -880 4683 -861
rect 4842 -691 4876 -672
rect 4842 -759 4876 -757
rect 4842 -795 4876 -793
rect 4842 -880 4876 -861
rect 5100 -691 5134 -672
rect 5100 -759 5134 -757
rect 5100 -795 5134 -793
rect 5100 -880 5134 -861
rect 5214 -702 5249 -668
rect 9573 -414 9607 -396
rect 9573 -486 9607 -464
rect 9573 -558 9607 -532
rect 9573 -630 9607 -600
rect 5248 -736 5249 -702
rect 5214 -770 5249 -736
rect 5248 -808 5249 -770
rect 5214 -838 5249 -808
rect 5248 -880 5249 -838
rect 5328 -691 5362 -672
rect 5328 -759 5362 -757
rect 5328 -795 5362 -793
rect 5328 -880 5362 -861
rect 5586 -691 5620 -672
rect 5586 -759 5620 -757
rect 5586 -795 5620 -793
rect 5586 -880 5620 -861
rect 5780 -691 5814 -672
rect 5780 -759 5814 -757
rect 5780 -795 5814 -793
rect 5780 -880 5814 -861
rect 6038 -691 6072 -672
rect 6038 -759 6072 -757
rect 6038 -795 6072 -793
rect 6038 -880 6072 -861
rect 6296 -691 6330 -672
rect 6296 -759 6330 -757
rect 6296 -795 6330 -793
rect 6296 -880 6330 -861
rect 6554 -691 6588 -672
rect 6554 -759 6588 -757
rect 6554 -795 6588 -793
rect 6554 -880 6588 -861
rect 6812 -691 6846 -672
rect 6812 -759 6846 -757
rect 6812 -795 6846 -793
rect 6812 -880 6846 -861
rect 7006 -691 7040 -672
rect 7006 -759 7040 -757
rect 7006 -795 7040 -793
rect 7006 -880 7040 -861
rect 7264 -691 7298 -672
rect 7264 -759 7298 -757
rect 7264 -795 7298 -793
rect 7264 -880 7298 -861
rect 7522 -691 7556 -672
rect 7522 -759 7556 -757
rect 7522 -795 7556 -793
rect 7522 -880 7556 -861
rect 7780 -691 7814 -672
rect 7780 -759 7814 -757
rect 7780 -795 7814 -793
rect 7780 -880 7814 -861
rect 7974 -691 8008 -672
rect 7974 -759 8008 -757
rect 7974 -795 8008 -793
rect 7974 -880 8008 -861
rect 8232 -691 8266 -672
rect 8232 -759 8266 -757
rect 8232 -795 8266 -793
rect 8232 -880 8266 -861
rect 8490 -691 8524 -672
rect 8490 -759 8524 -757
rect 8490 -795 8524 -793
rect 8490 -880 8524 -861
rect 8748 -691 8782 -672
rect 8748 -759 8782 -757
rect 8748 -795 8782 -793
rect 8748 -880 8782 -861
rect 9006 -691 9040 -672
rect 9006 -759 9040 -757
rect 9006 -795 9040 -793
rect 9006 -880 9040 -861
rect 9200 -691 9234 -672
rect 9200 -759 9234 -757
rect 9200 -795 9234 -793
rect 9200 -880 9234 -861
rect 9458 -691 9492 -672
rect 9458 -759 9492 -757
rect 9458 -795 9492 -793
rect 9458 -880 9492 -861
rect 9573 -702 9607 -668
rect 13931 -396 13932 -362
rect 13931 -414 13966 -396
rect 13931 -464 13932 -414
rect 13931 -486 13966 -464
rect 13931 -532 13932 -486
rect 13931 -558 13966 -532
rect 13931 -600 13932 -558
rect 13931 -630 13966 -600
rect 13931 -668 13932 -630
rect 9573 -770 9607 -736
rect 9573 -838 9607 -808
rect 9688 -691 9722 -672
rect 9688 -759 9722 -757
rect 9688 -795 9722 -793
rect 9688 -880 9722 -861
rect 9946 -691 9980 -672
rect 9946 -759 9980 -757
rect 9946 -795 9980 -793
rect 9946 -880 9980 -861
rect 10140 -691 10174 -672
rect 10140 -759 10174 -757
rect 10140 -795 10174 -793
rect 10140 -880 10174 -861
rect 10398 -691 10432 -672
rect 10398 -759 10432 -757
rect 10398 -795 10432 -793
rect 10398 -880 10432 -861
rect 10656 -691 10690 -672
rect 10656 -759 10690 -757
rect 10656 -795 10690 -793
rect 10656 -880 10690 -861
rect 10914 -691 10948 -672
rect 10914 -759 10948 -757
rect 10914 -795 10948 -793
rect 10914 -880 10948 -861
rect 11172 -691 11206 -672
rect 11172 -759 11206 -757
rect 11172 -795 11206 -793
rect 11172 -880 11206 -861
rect 11366 -691 11400 -672
rect 11366 -759 11400 -757
rect 11366 -795 11400 -793
rect 11366 -880 11400 -861
rect 11624 -691 11658 -672
rect 11624 -759 11658 -757
rect 11624 -795 11658 -793
rect 11624 -880 11658 -861
rect 11882 -691 11916 -672
rect 11882 -759 11916 -757
rect 11882 -795 11916 -793
rect 11882 -880 11916 -861
rect 12140 -691 12174 -672
rect 12140 -759 12174 -757
rect 12140 -795 12174 -793
rect 12140 -880 12174 -861
rect 12334 -691 12368 -672
rect 12334 -759 12368 -757
rect 12334 -795 12368 -793
rect 12334 -880 12368 -861
rect 12592 -691 12626 -672
rect 12592 -759 12626 -757
rect 12592 -795 12626 -793
rect 12592 -880 12626 -861
rect 12850 -691 12884 -672
rect 12850 -759 12884 -757
rect 12850 -795 12884 -793
rect 12850 -880 12884 -861
rect 13108 -691 13142 -672
rect 13108 -759 13142 -757
rect 13108 -795 13142 -793
rect 13108 -880 13142 -861
rect 13366 -691 13400 -672
rect 13366 -759 13400 -757
rect 13366 -795 13400 -793
rect 13366 -880 13400 -861
rect 13560 -691 13594 -672
rect 13560 -759 13594 -757
rect 13560 -795 13594 -793
rect 13560 -880 13594 -861
rect 13818 -691 13852 -672
rect 13818 -759 13852 -757
rect 13818 -795 13852 -793
rect 13818 -880 13852 -861
rect 13931 -702 13966 -668
rect 18290 -414 18324 -396
rect 18290 -486 18324 -464
rect 18290 -558 18324 -532
rect 18290 -630 18324 -600
rect 13931 -736 13932 -702
rect 13931 -770 13966 -736
rect 13931 -808 13932 -770
rect 13931 -838 13966 -808
rect 13931 -880 13932 -838
rect 14046 -691 14080 -672
rect 14046 -759 14080 -757
rect 14046 -795 14080 -793
rect 14046 -880 14080 -861
rect 14304 -691 14338 -672
rect 14304 -759 14338 -757
rect 14304 -795 14338 -793
rect 14304 -880 14338 -861
rect 14497 -691 14531 -672
rect 14497 -759 14531 -757
rect 14497 -795 14531 -793
rect 14497 -880 14531 -861
rect 14755 -691 14789 -672
rect 14755 -759 14789 -757
rect 14755 -795 14789 -793
rect 14755 -880 14789 -861
rect 15013 -691 15047 -672
rect 15013 -759 15047 -757
rect 15013 -795 15047 -793
rect 15013 -880 15047 -861
rect 15271 -691 15305 -672
rect 15271 -759 15305 -757
rect 15271 -795 15305 -793
rect 15271 -880 15305 -861
rect 15529 -691 15563 -672
rect 15529 -759 15563 -757
rect 15529 -795 15563 -793
rect 15529 -880 15563 -861
rect 15723 -691 15757 -672
rect 15723 -759 15757 -757
rect 15723 -795 15757 -793
rect 15723 -880 15757 -861
rect 15981 -691 16015 -672
rect 15981 -759 16015 -757
rect 15981 -795 16015 -793
rect 15981 -880 16015 -861
rect 16239 -691 16273 -672
rect 16239 -759 16273 -757
rect 16239 -795 16273 -793
rect 16239 -880 16273 -861
rect 16497 -691 16531 -672
rect 16497 -759 16531 -757
rect 16497 -795 16531 -793
rect 16497 -880 16531 -861
rect 16691 -691 16725 -672
rect 16691 -759 16725 -757
rect 16691 -795 16725 -793
rect 16691 -880 16725 -861
rect 16949 -691 16983 -672
rect 16949 -759 16983 -757
rect 16949 -795 16983 -793
rect 16949 -880 16983 -861
rect 17207 -691 17241 -672
rect 17207 -759 17241 -757
rect 17207 -795 17241 -793
rect 17207 -880 17241 -861
rect 17465 -691 17499 -672
rect 17465 -759 17499 -757
rect 17465 -795 17499 -793
rect 17465 -880 17499 -861
rect 17723 -691 17757 -672
rect 17723 -759 17757 -757
rect 17723 -795 17757 -793
rect 17723 -880 17757 -861
rect 17917 -691 17951 -672
rect 17917 -759 17951 -757
rect 17917 -795 17951 -793
rect 17917 -880 17951 -861
rect 18175 -691 18209 -672
rect 18175 -759 18209 -757
rect 18175 -795 18209 -793
rect 18175 -880 18209 -861
rect 18290 -702 18324 -668
rect 18290 -770 18324 -736
rect 18290 -838 18324 -808
rect 856 -906 890 -880
rect 5214 -906 5249 -880
rect 856 -974 890 -952
rect 1017 -957 1064 -923
rect 1100 -957 1134 -923
rect 1170 -957 1217 -923
rect 1469 -957 1516 -923
rect 1552 -957 1586 -923
rect 1622 -957 1669 -923
rect 1727 -957 1774 -923
rect 1810 -957 1844 -923
rect 1880 -957 1927 -923
rect 1985 -957 2032 -923
rect 2068 -957 2102 -923
rect 2138 -957 2185 -923
rect 2243 -957 2290 -923
rect 2326 -957 2360 -923
rect 2396 -957 2443 -923
rect 2695 -957 2742 -923
rect 2778 -957 2812 -923
rect 2848 -957 2895 -923
rect 2953 -957 3000 -923
rect 3036 -957 3070 -923
rect 3106 -957 3153 -923
rect 3211 -957 3258 -923
rect 3294 -957 3328 -923
rect 3364 -957 3411 -923
rect 3663 -957 3710 -923
rect 3746 -957 3780 -923
rect 3816 -957 3863 -923
rect 3921 -957 3968 -923
rect 4004 -957 4038 -923
rect 4074 -957 4121 -923
rect 4179 -957 4226 -923
rect 4262 -957 4296 -923
rect 4332 -957 4379 -923
rect 4437 -957 4484 -923
rect 4520 -957 4554 -923
rect 4590 -957 4637 -923
rect 4888 -957 4935 -923
rect 4971 -957 5005 -923
rect 5041 -957 5088 -923
rect 5248 -952 5249 -906
rect 9573 -906 9607 -880
rect 856 -1042 890 -1024
rect 856 -1110 890 -1096
rect 856 -1178 890 -1168
rect 856 -1246 890 -1240
rect 5214 -974 5249 -952
rect 5374 -957 5421 -923
rect 5457 -957 5491 -923
rect 5527 -957 5574 -923
rect 5826 -957 5873 -923
rect 5909 -957 5943 -923
rect 5979 -957 6026 -923
rect 6084 -957 6131 -923
rect 6167 -957 6201 -923
rect 6237 -957 6284 -923
rect 6342 -957 6389 -923
rect 6425 -957 6459 -923
rect 6495 -957 6542 -923
rect 6600 -957 6647 -923
rect 6683 -957 6717 -923
rect 6753 -957 6800 -923
rect 7052 -957 7099 -923
rect 7135 -957 7169 -923
rect 7205 -957 7252 -923
rect 7310 -957 7357 -923
rect 7393 -957 7427 -923
rect 7463 -957 7510 -923
rect 7568 -957 7615 -923
rect 7651 -957 7685 -923
rect 7721 -957 7768 -923
rect 8020 -957 8067 -923
rect 8103 -957 8137 -923
rect 8173 -957 8220 -923
rect 8278 -957 8325 -923
rect 8361 -957 8395 -923
rect 8431 -957 8478 -923
rect 8536 -957 8583 -923
rect 8619 -957 8653 -923
rect 8689 -957 8736 -923
rect 8794 -957 8841 -923
rect 8877 -957 8911 -923
rect 8947 -957 8994 -923
rect 9246 -957 9293 -923
rect 9329 -957 9363 -923
rect 9399 -957 9446 -923
rect 13931 -906 13966 -880
rect 5248 -1024 5249 -974
rect 5214 -1042 5249 -1024
rect 5248 -1096 5249 -1042
rect 5214 -1110 5249 -1096
rect 5248 -1168 5249 -1110
rect 5214 -1178 5249 -1168
rect 5248 -1240 5249 -1178
rect 5214 -1246 5249 -1240
rect 856 -1314 890 -1312
rect 1017 -1320 1064 -1286
rect 1100 -1320 1134 -1286
rect 1170 -1320 1217 -1286
rect 1469 -1320 1516 -1286
rect 1552 -1320 1586 -1286
rect 1622 -1320 1669 -1286
rect 1727 -1320 1774 -1286
rect 1810 -1320 1844 -1286
rect 1880 -1320 1927 -1286
rect 1985 -1320 2032 -1286
rect 2068 -1320 2102 -1286
rect 2138 -1320 2185 -1286
rect 2243 -1320 2290 -1286
rect 2326 -1320 2360 -1286
rect 2396 -1320 2443 -1286
rect 2695 -1320 2742 -1286
rect 2778 -1320 2812 -1286
rect 2848 -1320 2895 -1286
rect 2953 -1320 3000 -1286
rect 3036 -1320 3070 -1286
rect 3106 -1320 3153 -1286
rect 3211 -1320 3258 -1286
rect 3294 -1320 3328 -1286
rect 3364 -1320 3411 -1286
rect 3663 -1320 3710 -1286
rect 3746 -1320 3780 -1286
rect 3816 -1320 3863 -1286
rect 3921 -1320 3968 -1286
rect 4004 -1320 4038 -1286
rect 4074 -1320 4121 -1286
rect 4179 -1320 4226 -1286
rect 4262 -1320 4296 -1286
rect 4332 -1320 4379 -1286
rect 4437 -1320 4484 -1286
rect 4520 -1320 4554 -1286
rect 4590 -1320 4637 -1286
rect 4888 -1320 4935 -1286
rect 4971 -1320 5005 -1286
rect 5041 -1320 5088 -1286
rect 5248 -1312 5249 -1246
rect 9573 -974 9607 -952
rect 9734 -957 9781 -923
rect 9817 -957 9851 -923
rect 9887 -957 9934 -923
rect 10186 -957 10233 -923
rect 10269 -957 10303 -923
rect 10339 -957 10386 -923
rect 10444 -957 10491 -923
rect 10527 -957 10561 -923
rect 10597 -957 10644 -923
rect 10702 -957 10749 -923
rect 10785 -957 10819 -923
rect 10855 -957 10902 -923
rect 10960 -957 11007 -923
rect 11043 -957 11077 -923
rect 11113 -957 11160 -923
rect 11412 -957 11459 -923
rect 11495 -957 11529 -923
rect 11565 -957 11612 -923
rect 11670 -957 11717 -923
rect 11753 -957 11787 -923
rect 11823 -957 11870 -923
rect 11928 -957 11975 -923
rect 12011 -957 12045 -923
rect 12081 -957 12128 -923
rect 12380 -957 12427 -923
rect 12463 -957 12497 -923
rect 12533 -957 12580 -923
rect 12638 -957 12685 -923
rect 12721 -957 12755 -923
rect 12791 -957 12838 -923
rect 12896 -957 12943 -923
rect 12979 -957 13013 -923
rect 13049 -957 13096 -923
rect 13154 -957 13201 -923
rect 13237 -957 13271 -923
rect 13307 -957 13354 -923
rect 13606 -957 13653 -923
rect 13689 -957 13723 -923
rect 13759 -957 13806 -923
rect 13931 -952 13932 -906
rect 18290 -906 18324 -880
rect 9573 -1042 9607 -1024
rect 9573 -1110 9607 -1096
rect 9573 -1178 9607 -1168
rect 9573 -1246 9607 -1240
rect 5214 -1314 5249 -1312
rect 856 -1350 890 -1348
rect 5248 -1348 5249 -1314
rect 5374 -1320 5421 -1286
rect 5457 -1320 5491 -1286
rect 5527 -1320 5574 -1286
rect 5826 -1320 5873 -1286
rect 5909 -1320 5943 -1286
rect 5979 -1320 6026 -1286
rect 6084 -1320 6131 -1286
rect 6167 -1320 6201 -1286
rect 6237 -1320 6284 -1286
rect 6342 -1320 6389 -1286
rect 6425 -1320 6459 -1286
rect 6495 -1320 6542 -1286
rect 6600 -1320 6647 -1286
rect 6683 -1320 6717 -1286
rect 6753 -1320 6800 -1286
rect 7052 -1320 7099 -1286
rect 7135 -1320 7169 -1286
rect 7205 -1320 7252 -1286
rect 7310 -1320 7357 -1286
rect 7393 -1320 7427 -1286
rect 7463 -1320 7510 -1286
rect 7568 -1320 7615 -1286
rect 7651 -1320 7685 -1286
rect 7721 -1320 7768 -1286
rect 8020 -1320 8067 -1286
rect 8103 -1320 8137 -1286
rect 8173 -1320 8220 -1286
rect 8278 -1320 8325 -1286
rect 8361 -1320 8395 -1286
rect 8431 -1320 8478 -1286
rect 8536 -1320 8583 -1286
rect 8619 -1320 8653 -1286
rect 8689 -1320 8736 -1286
rect 8794 -1320 8841 -1286
rect 8877 -1320 8911 -1286
rect 8947 -1320 8994 -1286
rect 9246 -1320 9293 -1286
rect 9329 -1320 9363 -1286
rect 9399 -1320 9446 -1286
rect 13931 -974 13966 -952
rect 14092 -957 14139 -923
rect 14175 -957 14209 -923
rect 14245 -957 14292 -923
rect 14543 -957 14590 -923
rect 14626 -957 14660 -923
rect 14696 -957 14743 -923
rect 14801 -957 14848 -923
rect 14884 -957 14918 -923
rect 14954 -957 15001 -923
rect 15059 -957 15106 -923
rect 15142 -957 15176 -923
rect 15212 -957 15259 -923
rect 15317 -957 15364 -923
rect 15400 -957 15434 -923
rect 15470 -957 15517 -923
rect 15769 -957 15816 -923
rect 15852 -957 15886 -923
rect 15922 -957 15969 -923
rect 16027 -957 16074 -923
rect 16110 -957 16144 -923
rect 16180 -957 16227 -923
rect 16285 -957 16332 -923
rect 16368 -957 16402 -923
rect 16438 -957 16485 -923
rect 16737 -957 16784 -923
rect 16820 -957 16854 -923
rect 16890 -957 16937 -923
rect 16995 -957 17042 -923
rect 17078 -957 17112 -923
rect 17148 -957 17195 -923
rect 17253 -957 17300 -923
rect 17336 -957 17370 -923
rect 17406 -957 17453 -923
rect 17511 -957 17558 -923
rect 17594 -957 17628 -923
rect 17664 -957 17711 -923
rect 17963 -957 18010 -923
rect 18046 -957 18080 -923
rect 18116 -957 18163 -923
rect 13931 -1024 13932 -974
rect 13931 -1042 13966 -1024
rect 13931 -1096 13932 -1042
rect 13931 -1110 13966 -1096
rect 13931 -1168 13932 -1110
rect 13931 -1178 13966 -1168
rect 13931 -1240 13932 -1178
rect 13931 -1246 13966 -1240
rect 9573 -1314 9607 -1312
rect 5214 -1350 5249 -1348
rect 856 -1422 890 -1416
rect 856 -1494 890 -1484
rect 856 -1566 890 -1552
rect 971 -1382 1005 -1363
rect 971 -1450 1005 -1448
rect 971 -1486 1005 -1484
rect 971 -1571 1005 -1552
rect 1229 -1382 1263 -1363
rect 1229 -1450 1263 -1448
rect 1229 -1486 1263 -1484
rect 1229 -1571 1263 -1552
rect 1423 -1382 1457 -1363
rect 1423 -1450 1457 -1448
rect 1423 -1486 1457 -1484
rect 1423 -1571 1457 -1552
rect 1681 -1382 1715 -1363
rect 1681 -1450 1715 -1448
rect 1681 -1486 1715 -1484
rect 1681 -1571 1715 -1552
rect 1939 -1382 1973 -1363
rect 1939 -1450 1973 -1448
rect 1939 -1486 1973 -1484
rect 1939 -1571 1973 -1552
rect 2197 -1382 2231 -1363
rect 2197 -1450 2231 -1448
rect 2197 -1486 2231 -1484
rect 2197 -1571 2231 -1552
rect 2455 -1382 2489 -1363
rect 2455 -1450 2489 -1448
rect 2455 -1486 2489 -1484
rect 2455 -1571 2489 -1552
rect 2649 -1382 2683 -1363
rect 2649 -1450 2683 -1448
rect 2649 -1486 2683 -1484
rect 2649 -1571 2683 -1552
rect 2907 -1382 2941 -1363
rect 2907 -1450 2941 -1448
rect 2907 -1486 2941 -1484
rect 2907 -1571 2941 -1552
rect 3165 -1382 3199 -1363
rect 3165 -1450 3199 -1448
rect 3165 -1486 3199 -1484
rect 3165 -1571 3199 -1552
rect 3423 -1382 3457 -1363
rect 3423 -1450 3457 -1448
rect 3423 -1486 3457 -1484
rect 3423 -1571 3457 -1552
rect 3617 -1382 3651 -1363
rect 3617 -1450 3651 -1448
rect 3617 -1486 3651 -1484
rect 3617 -1571 3651 -1552
rect 3875 -1382 3909 -1363
rect 3875 -1450 3909 -1448
rect 3875 -1486 3909 -1484
rect 3875 -1571 3909 -1552
rect 4133 -1382 4167 -1363
rect 4133 -1450 4167 -1448
rect 4133 -1486 4167 -1484
rect 4133 -1571 4167 -1552
rect 4391 -1382 4425 -1363
rect 4391 -1450 4425 -1448
rect 4391 -1486 4425 -1484
rect 4391 -1571 4425 -1552
rect 4649 -1382 4683 -1363
rect 4649 -1450 4683 -1448
rect 4649 -1486 4683 -1484
rect 4649 -1571 4683 -1552
rect 4842 -1382 4876 -1363
rect 4842 -1450 4876 -1448
rect 4842 -1486 4876 -1484
rect 4842 -1571 4876 -1552
rect 5100 -1382 5134 -1363
rect 5100 -1450 5134 -1448
rect 5100 -1486 5134 -1484
rect 5100 -1571 5134 -1552
rect 5248 -1416 5249 -1350
rect 9734 -1320 9781 -1286
rect 9817 -1320 9851 -1286
rect 9887 -1320 9934 -1286
rect 10186 -1320 10233 -1286
rect 10269 -1320 10303 -1286
rect 10339 -1320 10386 -1286
rect 10444 -1320 10491 -1286
rect 10527 -1320 10561 -1286
rect 10597 -1320 10644 -1286
rect 10702 -1320 10749 -1286
rect 10785 -1320 10819 -1286
rect 10855 -1320 10902 -1286
rect 10960 -1320 11007 -1286
rect 11043 -1320 11077 -1286
rect 11113 -1320 11160 -1286
rect 11412 -1320 11459 -1286
rect 11495 -1320 11529 -1286
rect 11565 -1320 11612 -1286
rect 11670 -1320 11717 -1286
rect 11753 -1320 11787 -1286
rect 11823 -1320 11870 -1286
rect 11928 -1320 11975 -1286
rect 12011 -1320 12045 -1286
rect 12081 -1320 12128 -1286
rect 12380 -1320 12427 -1286
rect 12463 -1320 12497 -1286
rect 12533 -1320 12580 -1286
rect 12638 -1320 12685 -1286
rect 12721 -1320 12755 -1286
rect 12791 -1320 12838 -1286
rect 12896 -1320 12943 -1286
rect 12979 -1320 13013 -1286
rect 13049 -1320 13096 -1286
rect 13154 -1320 13201 -1286
rect 13237 -1320 13271 -1286
rect 13307 -1320 13354 -1286
rect 13606 -1320 13653 -1286
rect 13689 -1320 13723 -1286
rect 13759 -1320 13806 -1286
rect 13931 -1312 13932 -1246
rect 18290 -974 18324 -952
rect 18290 -1042 18324 -1024
rect 18290 -1110 18324 -1096
rect 18290 -1178 18324 -1168
rect 18290 -1246 18324 -1240
rect 13931 -1314 13966 -1312
rect 9573 -1350 9607 -1348
rect 5214 -1422 5249 -1416
rect 5248 -1484 5249 -1422
rect 5214 -1494 5249 -1484
rect 5248 -1552 5249 -1494
rect 5214 -1566 5249 -1552
rect 856 -1638 890 -1620
rect 856 -1710 890 -1688
rect 856 -1782 890 -1756
rect 856 -1854 890 -1824
rect 856 -1926 890 -1888
rect 5248 -1620 5249 -1566
rect 5328 -1382 5362 -1363
rect 5328 -1450 5362 -1448
rect 5328 -1486 5362 -1484
rect 5328 -1571 5362 -1552
rect 5586 -1382 5620 -1363
rect 5586 -1450 5620 -1448
rect 5586 -1486 5620 -1484
rect 5586 -1571 5620 -1552
rect 5780 -1382 5814 -1363
rect 5780 -1450 5814 -1448
rect 5780 -1486 5814 -1484
rect 5780 -1571 5814 -1552
rect 6038 -1382 6072 -1363
rect 6038 -1450 6072 -1448
rect 6038 -1486 6072 -1484
rect 6038 -1571 6072 -1552
rect 6296 -1382 6330 -1363
rect 6296 -1450 6330 -1448
rect 6296 -1486 6330 -1484
rect 6296 -1571 6330 -1552
rect 6554 -1382 6588 -1363
rect 6554 -1450 6588 -1448
rect 6554 -1486 6588 -1484
rect 6554 -1571 6588 -1552
rect 6812 -1382 6846 -1363
rect 6812 -1450 6846 -1448
rect 6812 -1486 6846 -1484
rect 6812 -1571 6846 -1552
rect 7006 -1382 7040 -1363
rect 7006 -1450 7040 -1448
rect 7006 -1486 7040 -1484
rect 7006 -1571 7040 -1552
rect 7264 -1382 7298 -1363
rect 7264 -1450 7298 -1448
rect 7264 -1486 7298 -1484
rect 7264 -1571 7298 -1552
rect 7522 -1382 7556 -1363
rect 7522 -1450 7556 -1448
rect 7522 -1486 7556 -1484
rect 7522 -1571 7556 -1552
rect 7780 -1382 7814 -1363
rect 7780 -1450 7814 -1448
rect 7780 -1486 7814 -1484
rect 7780 -1571 7814 -1552
rect 7974 -1382 8008 -1363
rect 7974 -1450 8008 -1448
rect 7974 -1486 8008 -1484
rect 7974 -1571 8008 -1552
rect 8232 -1382 8266 -1363
rect 8232 -1450 8266 -1448
rect 8232 -1486 8266 -1484
rect 8232 -1571 8266 -1552
rect 8490 -1382 8524 -1363
rect 8490 -1450 8524 -1448
rect 8490 -1486 8524 -1484
rect 8490 -1571 8524 -1552
rect 8748 -1382 8782 -1363
rect 8748 -1450 8782 -1448
rect 8748 -1486 8782 -1484
rect 8748 -1571 8782 -1552
rect 9006 -1382 9040 -1363
rect 9006 -1450 9040 -1448
rect 9006 -1486 9040 -1484
rect 9006 -1571 9040 -1552
rect 9200 -1382 9234 -1363
rect 9200 -1450 9234 -1448
rect 9200 -1486 9234 -1484
rect 9200 -1571 9234 -1552
rect 9458 -1382 9492 -1363
rect 9458 -1450 9492 -1448
rect 9458 -1486 9492 -1484
rect 9458 -1571 9492 -1552
rect 13931 -1348 13932 -1314
rect 14092 -1320 14139 -1286
rect 14175 -1320 14209 -1286
rect 14245 -1320 14292 -1286
rect 14543 -1320 14590 -1286
rect 14626 -1320 14660 -1286
rect 14696 -1320 14743 -1286
rect 14801 -1320 14848 -1286
rect 14884 -1320 14918 -1286
rect 14954 -1320 15001 -1286
rect 15059 -1320 15106 -1286
rect 15142 -1320 15176 -1286
rect 15212 -1320 15259 -1286
rect 15317 -1320 15364 -1286
rect 15400 -1320 15434 -1286
rect 15470 -1320 15517 -1286
rect 15769 -1320 15816 -1286
rect 15852 -1320 15886 -1286
rect 15922 -1320 15969 -1286
rect 16027 -1320 16074 -1286
rect 16110 -1320 16144 -1286
rect 16180 -1320 16227 -1286
rect 16285 -1320 16332 -1286
rect 16368 -1320 16402 -1286
rect 16438 -1320 16485 -1286
rect 16737 -1320 16784 -1286
rect 16820 -1320 16854 -1286
rect 16890 -1320 16937 -1286
rect 16995 -1320 17042 -1286
rect 17078 -1320 17112 -1286
rect 17148 -1320 17195 -1286
rect 17253 -1320 17300 -1286
rect 17336 -1320 17370 -1286
rect 17406 -1320 17453 -1286
rect 17511 -1320 17558 -1286
rect 17594 -1320 17628 -1286
rect 17664 -1320 17711 -1286
rect 17963 -1320 18010 -1286
rect 18046 -1320 18080 -1286
rect 18116 -1320 18163 -1286
rect 18290 -1314 18324 -1312
rect 13931 -1350 13966 -1348
rect 9573 -1422 9607 -1416
rect 9573 -1494 9607 -1484
rect 9573 -1566 9607 -1552
rect 5214 -1638 5249 -1620
rect 5248 -1688 5249 -1638
rect 5214 -1710 5249 -1688
rect 5248 -1756 5249 -1710
rect 5214 -1782 5249 -1756
rect 5248 -1824 5249 -1782
rect 5214 -1854 5249 -1824
rect 5248 -1888 5249 -1854
rect 5214 -1926 5249 -1888
rect 9688 -1382 9722 -1363
rect 9688 -1450 9722 -1448
rect 9688 -1486 9722 -1484
rect 9688 -1571 9722 -1552
rect 9946 -1382 9980 -1363
rect 9946 -1450 9980 -1448
rect 9946 -1486 9980 -1484
rect 9946 -1571 9980 -1552
rect 10140 -1382 10174 -1363
rect 10140 -1450 10174 -1448
rect 10140 -1486 10174 -1484
rect 10140 -1571 10174 -1552
rect 10398 -1382 10432 -1363
rect 10398 -1450 10432 -1448
rect 10398 -1486 10432 -1484
rect 10398 -1571 10432 -1552
rect 10656 -1382 10690 -1363
rect 10656 -1450 10690 -1448
rect 10656 -1486 10690 -1484
rect 10656 -1571 10690 -1552
rect 10914 -1382 10948 -1363
rect 10914 -1450 10948 -1448
rect 10914 -1486 10948 -1484
rect 10914 -1571 10948 -1552
rect 11172 -1382 11206 -1363
rect 11172 -1450 11206 -1448
rect 11172 -1486 11206 -1484
rect 11172 -1571 11206 -1552
rect 11366 -1382 11400 -1363
rect 11366 -1450 11400 -1448
rect 11366 -1486 11400 -1484
rect 11366 -1571 11400 -1552
rect 11624 -1382 11658 -1363
rect 11624 -1450 11658 -1448
rect 11624 -1486 11658 -1484
rect 11624 -1571 11658 -1552
rect 11882 -1382 11916 -1363
rect 11882 -1450 11916 -1448
rect 11882 -1486 11916 -1484
rect 11882 -1571 11916 -1552
rect 12140 -1382 12174 -1363
rect 12140 -1450 12174 -1448
rect 12140 -1486 12174 -1484
rect 12140 -1571 12174 -1552
rect 12334 -1382 12368 -1363
rect 12334 -1450 12368 -1448
rect 12334 -1486 12368 -1484
rect 12334 -1571 12368 -1552
rect 12592 -1382 12626 -1363
rect 12592 -1450 12626 -1448
rect 12592 -1486 12626 -1484
rect 12592 -1571 12626 -1552
rect 12850 -1382 12884 -1363
rect 12850 -1450 12884 -1448
rect 12850 -1486 12884 -1484
rect 12850 -1571 12884 -1552
rect 13108 -1382 13142 -1363
rect 13108 -1450 13142 -1448
rect 13108 -1486 13142 -1484
rect 13108 -1571 13142 -1552
rect 13366 -1382 13400 -1363
rect 13366 -1450 13400 -1448
rect 13366 -1486 13400 -1484
rect 13366 -1571 13400 -1552
rect 13560 -1382 13594 -1363
rect 13560 -1450 13594 -1448
rect 13560 -1486 13594 -1484
rect 13560 -1571 13594 -1552
rect 13818 -1382 13852 -1363
rect 13818 -1450 13852 -1448
rect 13818 -1486 13852 -1484
rect 13818 -1571 13852 -1552
rect 13931 -1416 13932 -1350
rect 18290 -1350 18324 -1348
rect 13931 -1422 13966 -1416
rect 13931 -1484 13932 -1422
rect 13931 -1494 13966 -1484
rect 13931 -1552 13932 -1494
rect 13931 -1566 13966 -1552
rect 9573 -1638 9607 -1620
rect 9573 -1710 9607 -1688
rect 9573 -1782 9607 -1756
rect 9573 -1854 9607 -1824
rect 9573 -1926 9607 -1888
rect 13931 -1620 13932 -1566
rect 14046 -1382 14080 -1363
rect 14046 -1450 14080 -1448
rect 14046 -1486 14080 -1484
rect 14046 -1571 14080 -1552
rect 14304 -1382 14338 -1363
rect 14304 -1450 14338 -1448
rect 14304 -1486 14338 -1484
rect 14304 -1571 14338 -1552
rect 14497 -1382 14531 -1363
rect 14497 -1450 14531 -1448
rect 14497 -1486 14531 -1484
rect 14497 -1571 14531 -1552
rect 14755 -1382 14789 -1363
rect 14755 -1450 14789 -1448
rect 14755 -1486 14789 -1484
rect 14755 -1571 14789 -1552
rect 15013 -1382 15047 -1363
rect 15013 -1450 15047 -1448
rect 15013 -1486 15047 -1484
rect 15013 -1571 15047 -1552
rect 15271 -1382 15305 -1363
rect 15271 -1450 15305 -1448
rect 15271 -1486 15305 -1484
rect 15271 -1571 15305 -1552
rect 15529 -1382 15563 -1363
rect 15529 -1450 15563 -1448
rect 15529 -1486 15563 -1484
rect 15529 -1571 15563 -1552
rect 15723 -1382 15757 -1363
rect 15723 -1450 15757 -1448
rect 15723 -1486 15757 -1484
rect 15723 -1571 15757 -1552
rect 15981 -1382 16015 -1363
rect 15981 -1450 16015 -1448
rect 15981 -1486 16015 -1484
rect 15981 -1571 16015 -1552
rect 16239 -1382 16273 -1363
rect 16239 -1450 16273 -1448
rect 16239 -1486 16273 -1484
rect 16239 -1571 16273 -1552
rect 16497 -1382 16531 -1363
rect 16497 -1450 16531 -1448
rect 16497 -1486 16531 -1484
rect 16497 -1571 16531 -1552
rect 16691 -1382 16725 -1363
rect 16691 -1450 16725 -1448
rect 16691 -1486 16725 -1484
rect 16691 -1571 16725 -1552
rect 16949 -1382 16983 -1363
rect 16949 -1450 16983 -1448
rect 16949 -1486 16983 -1484
rect 16949 -1571 16983 -1552
rect 17207 -1382 17241 -1363
rect 17207 -1450 17241 -1448
rect 17207 -1486 17241 -1484
rect 17207 -1571 17241 -1552
rect 17465 -1382 17499 -1363
rect 17465 -1450 17499 -1448
rect 17465 -1486 17499 -1484
rect 17465 -1571 17499 -1552
rect 17723 -1382 17757 -1363
rect 17723 -1450 17757 -1448
rect 17723 -1486 17757 -1484
rect 17723 -1571 17757 -1552
rect 17917 -1382 17951 -1363
rect 17917 -1450 17951 -1448
rect 17917 -1486 17951 -1484
rect 17917 -1571 17951 -1552
rect 18175 -1382 18209 -1363
rect 18175 -1450 18209 -1448
rect 18175 -1486 18209 -1484
rect 18175 -1571 18209 -1552
rect 18290 -1422 18324 -1416
rect 18290 -1494 18324 -1484
rect 18290 -1566 18324 -1552
rect 13931 -1638 13966 -1620
rect 13931 -1688 13932 -1638
rect 13931 -1710 13966 -1688
rect 13931 -1756 13932 -1710
rect 13931 -1782 13966 -1756
rect 13931 -1824 13932 -1782
rect 13931 -1854 13966 -1824
rect 13931 -1888 13932 -1854
rect 13931 -1926 13966 -1888
rect 18290 -1638 18324 -1620
rect 18290 -1710 18324 -1688
rect 18290 -1782 18324 -1756
rect 18290 -1854 18324 -1824
rect 18290 -1926 18324 -1888
rect 890 -1960 977 -1926
rect 1011 -1960 1045 -1926
rect 1079 -1960 1113 -1926
rect 1147 -1960 1181 -1926
rect 1215 -1960 1249 -1926
rect 1283 -1960 1317 -1926
rect 1351 -1960 1385 -1926
rect 1419 -1960 1453 -1926
rect 1487 -1960 1521 -1926
rect 1555 -1960 1589 -1926
rect 1623 -1960 1657 -1926
rect 1691 -1960 1725 -1926
rect 1759 -1960 1793 -1926
rect 1827 -1960 1861 -1926
rect 1895 -1960 1929 -1926
rect 1963 -1960 1997 -1926
rect 2031 -1960 2065 -1926
rect 2099 -1960 2133 -1926
rect 2167 -1960 2201 -1926
rect 2235 -1960 2269 -1926
rect 2303 -1960 2337 -1926
rect 2371 -1960 2405 -1926
rect 2439 -1960 2473 -1926
rect 2507 -1960 2541 -1926
rect 2575 -1960 2609 -1926
rect 2643 -1960 2677 -1926
rect 2711 -1960 2745 -1926
rect 2779 -1960 2813 -1926
rect 2847 -1960 2881 -1926
rect 2915 -1960 2949 -1926
rect 2983 -1960 3017 -1926
rect 3051 -1960 3085 -1926
rect 3119 -1960 3153 -1926
rect 3187 -1960 3221 -1926
rect 3255 -1960 3289 -1926
rect 3323 -1960 3357 -1926
rect 3391 -1960 3425 -1926
rect 3459 -1960 3493 -1926
rect 3527 -1960 3561 -1926
rect 3595 -1960 3629 -1926
rect 3663 -1960 3697 -1926
rect 3731 -1960 3765 -1926
rect 3799 -1960 3833 -1926
rect 3867 -1960 3901 -1926
rect 3935 -1960 3969 -1926
rect 4003 -1960 4037 -1926
rect 4071 -1960 4105 -1926
rect 4139 -1960 4173 -1926
rect 4207 -1960 4241 -1926
rect 4275 -1960 4309 -1926
rect 4343 -1960 4377 -1926
rect 4411 -1960 4445 -1926
rect 4479 -1960 4513 -1926
rect 4547 -1960 4581 -1926
rect 4615 -1960 4649 -1926
rect 4683 -1960 4717 -1926
rect 4751 -1960 4785 -1926
rect 4819 -1960 4853 -1926
rect 4887 -1960 4921 -1926
rect 4955 -1960 4989 -1926
rect 5023 -1960 5057 -1926
rect 5091 -1960 5214 -1926
rect 5248 -1960 5372 -1926
rect 5406 -1960 5440 -1926
rect 5474 -1960 5508 -1926
rect 5542 -1960 5576 -1926
rect 5610 -1960 5644 -1926
rect 5678 -1960 5712 -1926
rect 5746 -1960 5780 -1926
rect 5814 -1960 5848 -1926
rect 5882 -1960 5916 -1926
rect 5950 -1960 5984 -1926
rect 6018 -1960 6052 -1926
rect 6086 -1960 6120 -1926
rect 6154 -1960 6188 -1926
rect 6222 -1960 6256 -1926
rect 6290 -1960 6324 -1926
rect 6358 -1960 6392 -1926
rect 6426 -1960 6460 -1926
rect 6494 -1960 6528 -1926
rect 6562 -1960 6596 -1926
rect 6630 -1960 6664 -1926
rect 6698 -1960 6732 -1926
rect 6766 -1960 6800 -1926
rect 6834 -1960 6868 -1926
rect 6902 -1960 6936 -1926
rect 6970 -1960 7004 -1926
rect 7038 -1960 7072 -1926
rect 7106 -1960 7140 -1926
rect 7174 -1960 7208 -1926
rect 7242 -1960 7276 -1926
rect 7310 -1960 7344 -1926
rect 7378 -1960 7412 -1926
rect 7446 -1960 7480 -1926
rect 7514 -1960 7548 -1926
rect 7582 -1960 7616 -1926
rect 7650 -1960 7684 -1926
rect 7718 -1960 7752 -1926
rect 7786 -1960 7820 -1926
rect 7854 -1960 7888 -1926
rect 7922 -1960 7956 -1926
rect 7990 -1960 8024 -1926
rect 8058 -1960 8092 -1926
rect 8126 -1960 8160 -1926
rect 8194 -1960 8228 -1926
rect 8262 -1960 8296 -1926
rect 8330 -1960 8364 -1926
rect 8398 -1960 8432 -1926
rect 8466 -1960 8500 -1926
rect 8534 -1960 8568 -1926
rect 8602 -1960 8636 -1926
rect 8670 -1960 8704 -1926
rect 8738 -1960 8772 -1926
rect 8806 -1960 8840 -1926
rect 8874 -1960 8908 -1926
rect 8942 -1960 8976 -1926
rect 9010 -1960 9044 -1926
rect 9078 -1960 9112 -1926
rect 9146 -1960 9180 -1926
rect 9214 -1960 9248 -1926
rect 9282 -1960 9316 -1926
rect 9350 -1960 9384 -1926
rect 9418 -1960 9452 -1926
rect 9486 -1960 9573 -1926
rect 9607 -1960 9694 -1926
rect 9728 -1960 9762 -1926
rect 9796 -1960 9830 -1926
rect 9864 -1960 9898 -1926
rect 9932 -1960 9966 -1926
rect 10000 -1960 10034 -1926
rect 10068 -1960 10102 -1926
rect 10136 -1960 10170 -1926
rect 10204 -1960 10238 -1926
rect 10272 -1960 10306 -1926
rect 10340 -1960 10374 -1926
rect 10408 -1960 10442 -1926
rect 10476 -1960 10510 -1926
rect 10544 -1960 10578 -1926
rect 10612 -1960 10646 -1926
rect 10680 -1960 10714 -1926
rect 10748 -1960 10782 -1926
rect 10816 -1960 10850 -1926
rect 10884 -1960 10918 -1926
rect 10952 -1960 10986 -1926
rect 11020 -1960 11054 -1926
rect 11088 -1960 11122 -1926
rect 11156 -1960 11190 -1926
rect 11224 -1960 11258 -1926
rect 11292 -1960 11326 -1926
rect 11360 -1960 11394 -1926
rect 11428 -1960 11462 -1926
rect 11496 -1960 11530 -1926
rect 11564 -1960 11598 -1926
rect 11632 -1960 11666 -1926
rect 11700 -1960 11734 -1926
rect 11768 -1960 11802 -1926
rect 11836 -1960 11870 -1926
rect 11904 -1960 11938 -1926
rect 11972 -1960 12006 -1926
rect 12040 -1960 12074 -1926
rect 12108 -1960 12142 -1926
rect 12176 -1960 12210 -1926
rect 12244 -1960 12278 -1926
rect 12312 -1960 12346 -1926
rect 12380 -1960 12414 -1926
rect 12448 -1960 12482 -1926
rect 12516 -1960 12550 -1926
rect 12584 -1960 12618 -1926
rect 12652 -1960 12686 -1926
rect 12720 -1960 12754 -1926
rect 12788 -1960 12822 -1926
rect 12856 -1960 12890 -1926
rect 12924 -1960 12958 -1926
rect 12992 -1960 13026 -1926
rect 13060 -1960 13094 -1926
rect 13128 -1960 13162 -1926
rect 13196 -1960 13230 -1926
rect 13264 -1960 13298 -1926
rect 13332 -1960 13366 -1926
rect 13400 -1960 13434 -1926
rect 13468 -1960 13502 -1926
rect 13536 -1960 13570 -1926
rect 13604 -1960 13638 -1926
rect 13672 -1960 13706 -1926
rect 13740 -1960 13774 -1926
rect 13808 -1960 13932 -1926
rect 13966 -1960 14089 -1926
rect 14123 -1960 14157 -1926
rect 14191 -1960 14225 -1926
rect 14259 -1960 14293 -1926
rect 14327 -1960 14361 -1926
rect 14395 -1960 14429 -1926
rect 14463 -1960 14497 -1926
rect 14531 -1960 14565 -1926
rect 14599 -1960 14633 -1926
rect 14667 -1960 14701 -1926
rect 14735 -1960 14769 -1926
rect 14803 -1960 14837 -1926
rect 14871 -1960 14905 -1926
rect 14939 -1960 14973 -1926
rect 15007 -1960 15041 -1926
rect 15075 -1960 15109 -1926
rect 15143 -1960 15177 -1926
rect 15211 -1960 15245 -1926
rect 15279 -1960 15313 -1926
rect 15347 -1960 15381 -1926
rect 15415 -1960 15449 -1926
rect 15483 -1960 15517 -1926
rect 15551 -1960 15585 -1926
rect 15619 -1960 15653 -1926
rect 15687 -1960 15721 -1926
rect 15755 -1960 15789 -1926
rect 15823 -1960 15857 -1926
rect 15891 -1960 15925 -1926
rect 15959 -1960 15993 -1926
rect 16027 -1960 16061 -1926
rect 16095 -1960 16129 -1926
rect 16163 -1960 16197 -1926
rect 16231 -1960 16265 -1926
rect 16299 -1960 16333 -1926
rect 16367 -1960 16401 -1926
rect 16435 -1960 16469 -1926
rect 16503 -1960 16537 -1926
rect 16571 -1960 16605 -1926
rect 16639 -1960 16673 -1926
rect 16707 -1960 16741 -1926
rect 16775 -1960 16809 -1926
rect 16843 -1960 16877 -1926
rect 16911 -1960 16945 -1926
rect 16979 -1960 17013 -1926
rect 17047 -1960 17081 -1926
rect 17115 -1960 17149 -1926
rect 17183 -1960 17217 -1926
rect 17251 -1960 17285 -1926
rect 17319 -1960 17353 -1926
rect 17387 -1960 17421 -1926
rect 17455 -1960 17489 -1926
rect 17523 -1960 17557 -1926
rect 17591 -1960 17625 -1926
rect 17659 -1960 17693 -1926
rect 17727 -1960 17761 -1926
rect 17795 -1960 17829 -1926
rect 17863 -1960 17897 -1926
rect 17931 -1960 17965 -1926
rect 17999 -1960 18033 -1926
rect 18067 -1960 18101 -1926
rect 18135 -1960 18169 -1926
rect 18203 -1960 18290 -1926
rect 856 -1998 890 -1960
rect 856 -2062 890 -2032
rect 856 -2130 890 -2104
rect 856 -2198 890 -2176
rect 856 -2266 890 -2248
rect 5214 -1998 5249 -1960
rect 5248 -2032 5249 -1998
rect 5214 -2062 5249 -2032
rect 5248 -2104 5249 -2062
rect 5214 -2130 5249 -2104
rect 5248 -2176 5249 -2130
rect 5214 -2198 5249 -2176
rect 5248 -2248 5249 -2198
rect 5214 -2266 5249 -2248
rect 856 -2334 890 -2320
rect 856 -2402 890 -2392
rect 856 -2470 890 -2464
rect 971 -2338 1005 -2319
rect 971 -2406 1005 -2404
rect 971 -2442 1005 -2440
rect 971 -2527 1005 -2508
rect 1229 -2338 1263 -2319
rect 1229 -2406 1263 -2404
rect 1229 -2442 1263 -2440
rect 1229 -2527 1263 -2508
rect 1423 -2338 1457 -2319
rect 1423 -2406 1457 -2404
rect 1423 -2442 1457 -2440
rect 1423 -2527 1457 -2508
rect 1681 -2338 1715 -2319
rect 1681 -2406 1715 -2404
rect 1681 -2442 1715 -2440
rect 1681 -2527 1715 -2508
rect 1939 -2338 1973 -2319
rect 1939 -2406 1973 -2404
rect 1939 -2442 1973 -2440
rect 1939 -2527 1973 -2508
rect 2197 -2338 2231 -2319
rect 2197 -2406 2231 -2404
rect 2197 -2442 2231 -2440
rect 2197 -2527 2231 -2508
rect 2455 -2338 2489 -2319
rect 2455 -2406 2489 -2404
rect 2455 -2442 2489 -2440
rect 2455 -2527 2489 -2508
rect 2649 -2338 2683 -2319
rect 2649 -2406 2683 -2404
rect 2649 -2442 2683 -2440
rect 2649 -2527 2683 -2508
rect 2907 -2338 2941 -2319
rect 2907 -2406 2941 -2404
rect 2907 -2442 2941 -2440
rect 2907 -2527 2941 -2508
rect 3165 -2338 3199 -2319
rect 3165 -2406 3199 -2404
rect 3165 -2442 3199 -2440
rect 3165 -2527 3199 -2508
rect 3423 -2338 3457 -2319
rect 3423 -2406 3457 -2404
rect 3423 -2442 3457 -2440
rect 3423 -2527 3457 -2508
rect 3617 -2338 3651 -2319
rect 3617 -2406 3651 -2404
rect 3617 -2442 3651 -2440
rect 3617 -2527 3651 -2508
rect 3875 -2338 3909 -2319
rect 3875 -2406 3909 -2404
rect 3875 -2442 3909 -2440
rect 3875 -2527 3909 -2508
rect 4133 -2338 4167 -2319
rect 4133 -2406 4167 -2404
rect 4133 -2442 4167 -2440
rect 4133 -2527 4167 -2508
rect 4391 -2338 4425 -2319
rect 4391 -2406 4425 -2404
rect 4391 -2442 4425 -2440
rect 4391 -2527 4425 -2508
rect 4649 -2338 4683 -2319
rect 4649 -2406 4683 -2404
rect 4649 -2442 4683 -2440
rect 4649 -2527 4683 -2508
rect 4842 -2338 4876 -2319
rect 4842 -2406 4876 -2404
rect 4842 -2442 4876 -2440
rect 4842 -2527 4876 -2508
rect 5100 -2338 5134 -2319
rect 5100 -2406 5134 -2404
rect 5100 -2442 5134 -2440
rect 5100 -2527 5134 -2508
rect 5248 -2320 5249 -2266
rect 9573 -1998 9607 -1960
rect 9573 -2062 9607 -2032
rect 9573 -2130 9607 -2104
rect 9573 -2198 9607 -2176
rect 9573 -2266 9607 -2248
rect 5214 -2334 5249 -2320
rect 5248 -2392 5249 -2334
rect 5214 -2402 5249 -2392
rect 5248 -2464 5249 -2402
rect 5214 -2470 5249 -2464
rect 856 -2538 890 -2536
rect 5248 -2536 5249 -2470
rect 5328 -2338 5362 -2319
rect 5328 -2406 5362 -2404
rect 5328 -2442 5362 -2440
rect 5328 -2527 5362 -2508
rect 5586 -2338 5620 -2319
rect 5586 -2406 5620 -2404
rect 5586 -2442 5620 -2440
rect 5586 -2527 5620 -2508
rect 5780 -2338 5814 -2319
rect 5780 -2406 5814 -2404
rect 5780 -2442 5814 -2440
rect 5780 -2527 5814 -2508
rect 6038 -2338 6072 -2319
rect 6038 -2406 6072 -2404
rect 6038 -2442 6072 -2440
rect 6038 -2527 6072 -2508
rect 6296 -2338 6330 -2319
rect 6296 -2406 6330 -2404
rect 6296 -2442 6330 -2440
rect 6296 -2527 6330 -2508
rect 6554 -2338 6588 -2319
rect 6554 -2406 6588 -2404
rect 6554 -2442 6588 -2440
rect 6554 -2527 6588 -2508
rect 6812 -2338 6846 -2319
rect 6812 -2406 6846 -2404
rect 6812 -2442 6846 -2440
rect 6812 -2527 6846 -2508
rect 7006 -2338 7040 -2319
rect 7006 -2406 7040 -2404
rect 7006 -2442 7040 -2440
rect 7006 -2527 7040 -2508
rect 7264 -2338 7298 -2319
rect 7264 -2406 7298 -2404
rect 7264 -2442 7298 -2440
rect 7264 -2527 7298 -2508
rect 7522 -2338 7556 -2319
rect 7522 -2406 7556 -2404
rect 7522 -2442 7556 -2440
rect 7522 -2527 7556 -2508
rect 7780 -2338 7814 -2319
rect 7780 -2406 7814 -2404
rect 7780 -2442 7814 -2440
rect 7780 -2527 7814 -2508
rect 7974 -2338 8008 -2319
rect 7974 -2406 8008 -2404
rect 7974 -2442 8008 -2440
rect 7974 -2527 8008 -2508
rect 8232 -2338 8266 -2319
rect 8232 -2406 8266 -2404
rect 8232 -2442 8266 -2440
rect 8232 -2527 8266 -2508
rect 8490 -2338 8524 -2319
rect 8490 -2406 8524 -2404
rect 8490 -2442 8524 -2440
rect 8490 -2527 8524 -2508
rect 8748 -2338 8782 -2319
rect 8748 -2406 8782 -2404
rect 8748 -2442 8782 -2440
rect 8748 -2527 8782 -2508
rect 9006 -2338 9040 -2319
rect 9006 -2406 9040 -2404
rect 9006 -2442 9040 -2440
rect 9006 -2527 9040 -2508
rect 9200 -2338 9234 -2319
rect 9200 -2406 9234 -2404
rect 9200 -2442 9234 -2440
rect 9200 -2527 9234 -2508
rect 9458 -2338 9492 -2319
rect 9458 -2406 9492 -2404
rect 9458 -2442 9492 -2440
rect 9458 -2527 9492 -2508
rect 13931 -1998 13966 -1960
rect 13931 -2032 13932 -1998
rect 13931 -2062 13966 -2032
rect 13931 -2104 13932 -2062
rect 13931 -2130 13966 -2104
rect 13931 -2176 13932 -2130
rect 13931 -2198 13966 -2176
rect 13931 -2248 13932 -2198
rect 13931 -2266 13966 -2248
rect 9573 -2334 9607 -2320
rect 9573 -2402 9607 -2392
rect 9573 -2470 9607 -2464
rect 5214 -2538 5249 -2536
rect 856 -2574 890 -2572
rect 1017 -2604 1064 -2570
rect 1100 -2604 1134 -2570
rect 1170 -2604 1217 -2570
rect 1469 -2604 1516 -2570
rect 1552 -2604 1586 -2570
rect 1622 -2604 1669 -2570
rect 1727 -2604 1774 -2570
rect 1810 -2604 1844 -2570
rect 1880 -2604 1927 -2570
rect 1985 -2604 2032 -2570
rect 2068 -2604 2102 -2570
rect 2138 -2604 2185 -2570
rect 2243 -2604 2290 -2570
rect 2326 -2604 2360 -2570
rect 2396 -2604 2443 -2570
rect 2695 -2604 2742 -2570
rect 2778 -2604 2812 -2570
rect 2848 -2604 2895 -2570
rect 2953 -2604 3000 -2570
rect 3036 -2604 3070 -2570
rect 3106 -2604 3153 -2570
rect 3211 -2604 3258 -2570
rect 3294 -2604 3328 -2570
rect 3364 -2604 3411 -2570
rect 3663 -2604 3710 -2570
rect 3746 -2604 3780 -2570
rect 3816 -2604 3863 -2570
rect 3921 -2604 3968 -2570
rect 4004 -2604 4038 -2570
rect 4074 -2604 4121 -2570
rect 4179 -2604 4226 -2570
rect 4262 -2604 4296 -2570
rect 4332 -2604 4379 -2570
rect 4437 -2604 4484 -2570
rect 4520 -2604 4554 -2570
rect 4590 -2604 4637 -2570
rect 4888 -2604 4935 -2570
rect 4971 -2604 5005 -2570
rect 5041 -2604 5088 -2570
rect 5248 -2572 5249 -2538
rect 9688 -2338 9722 -2319
rect 9688 -2406 9722 -2404
rect 9688 -2442 9722 -2440
rect 9688 -2527 9722 -2508
rect 9946 -2338 9980 -2319
rect 9946 -2406 9980 -2404
rect 9946 -2442 9980 -2440
rect 9946 -2527 9980 -2508
rect 10140 -2338 10174 -2319
rect 10140 -2406 10174 -2404
rect 10140 -2442 10174 -2440
rect 10140 -2527 10174 -2508
rect 10398 -2338 10432 -2319
rect 10398 -2406 10432 -2404
rect 10398 -2442 10432 -2440
rect 10398 -2527 10432 -2508
rect 10656 -2338 10690 -2319
rect 10656 -2406 10690 -2404
rect 10656 -2442 10690 -2440
rect 10656 -2527 10690 -2508
rect 10914 -2338 10948 -2319
rect 10914 -2406 10948 -2404
rect 10914 -2442 10948 -2440
rect 10914 -2527 10948 -2508
rect 11172 -2338 11206 -2319
rect 11172 -2406 11206 -2404
rect 11172 -2442 11206 -2440
rect 11172 -2527 11206 -2508
rect 11366 -2338 11400 -2319
rect 11366 -2406 11400 -2404
rect 11366 -2442 11400 -2440
rect 11366 -2527 11400 -2508
rect 11624 -2338 11658 -2319
rect 11624 -2406 11658 -2404
rect 11624 -2442 11658 -2440
rect 11624 -2527 11658 -2508
rect 11882 -2338 11916 -2319
rect 11882 -2406 11916 -2404
rect 11882 -2442 11916 -2440
rect 11882 -2527 11916 -2508
rect 12140 -2338 12174 -2319
rect 12140 -2406 12174 -2404
rect 12140 -2442 12174 -2440
rect 12140 -2527 12174 -2508
rect 12334 -2338 12368 -2319
rect 12334 -2406 12368 -2404
rect 12334 -2442 12368 -2440
rect 12334 -2527 12368 -2508
rect 12592 -2338 12626 -2319
rect 12592 -2406 12626 -2404
rect 12592 -2442 12626 -2440
rect 12592 -2527 12626 -2508
rect 12850 -2338 12884 -2319
rect 12850 -2406 12884 -2404
rect 12850 -2442 12884 -2440
rect 12850 -2527 12884 -2508
rect 13108 -2338 13142 -2319
rect 13108 -2406 13142 -2404
rect 13108 -2442 13142 -2440
rect 13108 -2527 13142 -2508
rect 13366 -2338 13400 -2319
rect 13366 -2406 13400 -2404
rect 13366 -2442 13400 -2440
rect 13366 -2527 13400 -2508
rect 13560 -2338 13594 -2319
rect 13560 -2406 13594 -2404
rect 13560 -2442 13594 -2440
rect 13560 -2527 13594 -2508
rect 13818 -2338 13852 -2319
rect 13818 -2406 13852 -2404
rect 13818 -2442 13852 -2440
rect 13818 -2527 13852 -2508
rect 13931 -2320 13932 -2266
rect 18290 -1998 18324 -1960
rect 18290 -2062 18324 -2032
rect 18290 -2130 18324 -2104
rect 18290 -2198 18324 -2176
rect 18290 -2266 18324 -2248
rect 13931 -2334 13966 -2320
rect 13931 -2392 13932 -2334
rect 13931 -2402 13966 -2392
rect 13931 -2464 13932 -2402
rect 13931 -2470 13966 -2464
rect 9573 -2538 9607 -2536
rect 5214 -2574 5249 -2572
rect 856 -2646 890 -2640
rect 856 -2718 890 -2708
rect 856 -2790 890 -2776
rect 856 -2862 890 -2844
rect 856 -2934 890 -2912
rect 5248 -2640 5249 -2574
rect 5374 -2604 5421 -2570
rect 5457 -2604 5491 -2570
rect 5527 -2604 5574 -2570
rect 5826 -2604 5873 -2570
rect 5909 -2604 5943 -2570
rect 5979 -2604 6026 -2570
rect 6084 -2604 6131 -2570
rect 6167 -2604 6201 -2570
rect 6237 -2604 6284 -2570
rect 6342 -2604 6389 -2570
rect 6425 -2604 6459 -2570
rect 6495 -2604 6542 -2570
rect 6600 -2604 6647 -2570
rect 6683 -2604 6717 -2570
rect 6753 -2604 6800 -2570
rect 7052 -2604 7099 -2570
rect 7135 -2604 7169 -2570
rect 7205 -2604 7252 -2570
rect 7310 -2604 7357 -2570
rect 7393 -2604 7427 -2570
rect 7463 -2604 7510 -2570
rect 7568 -2604 7615 -2570
rect 7651 -2604 7685 -2570
rect 7721 -2604 7768 -2570
rect 8020 -2604 8067 -2570
rect 8103 -2604 8137 -2570
rect 8173 -2604 8220 -2570
rect 8278 -2604 8325 -2570
rect 8361 -2604 8395 -2570
rect 8431 -2604 8478 -2570
rect 8536 -2604 8583 -2570
rect 8619 -2604 8653 -2570
rect 8689 -2604 8736 -2570
rect 8794 -2604 8841 -2570
rect 8877 -2604 8911 -2570
rect 8947 -2604 8994 -2570
rect 9246 -2604 9293 -2570
rect 9329 -2604 9363 -2570
rect 9399 -2604 9446 -2570
rect 13931 -2536 13932 -2470
rect 14046 -2338 14080 -2319
rect 14046 -2406 14080 -2404
rect 14046 -2442 14080 -2440
rect 14046 -2527 14080 -2508
rect 14304 -2338 14338 -2319
rect 14304 -2406 14338 -2404
rect 14304 -2442 14338 -2440
rect 14304 -2527 14338 -2508
rect 14497 -2338 14531 -2319
rect 14497 -2406 14531 -2404
rect 14497 -2442 14531 -2440
rect 14497 -2527 14531 -2508
rect 14755 -2338 14789 -2319
rect 14755 -2406 14789 -2404
rect 14755 -2442 14789 -2440
rect 14755 -2527 14789 -2508
rect 15013 -2338 15047 -2319
rect 15013 -2406 15047 -2404
rect 15013 -2442 15047 -2440
rect 15013 -2527 15047 -2508
rect 15271 -2338 15305 -2319
rect 15271 -2406 15305 -2404
rect 15271 -2442 15305 -2440
rect 15271 -2527 15305 -2508
rect 15529 -2338 15563 -2319
rect 15529 -2406 15563 -2404
rect 15529 -2442 15563 -2440
rect 15529 -2527 15563 -2508
rect 15723 -2338 15757 -2319
rect 15723 -2406 15757 -2404
rect 15723 -2442 15757 -2440
rect 15723 -2527 15757 -2508
rect 15981 -2338 16015 -2319
rect 15981 -2406 16015 -2404
rect 15981 -2442 16015 -2440
rect 15981 -2527 16015 -2508
rect 16239 -2338 16273 -2319
rect 16239 -2406 16273 -2404
rect 16239 -2442 16273 -2440
rect 16239 -2527 16273 -2508
rect 16497 -2338 16531 -2319
rect 16497 -2406 16531 -2404
rect 16497 -2442 16531 -2440
rect 16497 -2527 16531 -2508
rect 16691 -2338 16725 -2319
rect 16691 -2406 16725 -2404
rect 16691 -2442 16725 -2440
rect 16691 -2527 16725 -2508
rect 16949 -2338 16983 -2319
rect 16949 -2406 16983 -2404
rect 16949 -2442 16983 -2440
rect 16949 -2527 16983 -2508
rect 17207 -2338 17241 -2319
rect 17207 -2406 17241 -2404
rect 17207 -2442 17241 -2440
rect 17207 -2527 17241 -2508
rect 17465 -2338 17499 -2319
rect 17465 -2406 17499 -2404
rect 17465 -2442 17499 -2440
rect 17465 -2527 17499 -2508
rect 17723 -2338 17757 -2319
rect 17723 -2406 17757 -2404
rect 17723 -2442 17757 -2440
rect 17723 -2527 17757 -2508
rect 17917 -2338 17951 -2319
rect 17917 -2406 17951 -2404
rect 17917 -2442 17951 -2440
rect 17917 -2527 17951 -2508
rect 18175 -2338 18209 -2319
rect 18175 -2406 18209 -2404
rect 18175 -2442 18209 -2440
rect 18175 -2527 18209 -2508
rect 18290 -2334 18324 -2320
rect 18290 -2402 18324 -2392
rect 18290 -2470 18324 -2464
rect 13931 -2538 13966 -2536
rect 9573 -2574 9607 -2572
rect 5214 -2646 5249 -2640
rect 5248 -2708 5249 -2646
rect 5214 -2718 5249 -2708
rect 5248 -2776 5249 -2718
rect 5214 -2790 5249 -2776
rect 5248 -2844 5249 -2790
rect 5214 -2862 5249 -2844
rect 5248 -2912 5249 -2862
rect 1017 -2967 1064 -2933
rect 1100 -2967 1134 -2933
rect 1170 -2967 1217 -2933
rect 1469 -2967 1516 -2933
rect 1552 -2967 1586 -2933
rect 1622 -2967 1669 -2933
rect 1727 -2967 1774 -2933
rect 1810 -2967 1844 -2933
rect 1880 -2967 1927 -2933
rect 1985 -2967 2032 -2933
rect 2068 -2967 2102 -2933
rect 2138 -2967 2185 -2933
rect 2243 -2967 2290 -2933
rect 2326 -2967 2360 -2933
rect 2396 -2967 2443 -2933
rect 2695 -2967 2742 -2933
rect 2778 -2967 2812 -2933
rect 2848 -2967 2895 -2933
rect 2953 -2967 3000 -2933
rect 3036 -2967 3070 -2933
rect 3106 -2967 3153 -2933
rect 3211 -2967 3258 -2933
rect 3294 -2967 3328 -2933
rect 3364 -2967 3411 -2933
rect 3663 -2967 3710 -2933
rect 3746 -2967 3780 -2933
rect 3816 -2967 3863 -2933
rect 3921 -2967 3968 -2933
rect 4004 -2967 4038 -2933
rect 4074 -2967 4121 -2933
rect 4179 -2967 4226 -2933
rect 4262 -2967 4296 -2933
rect 4332 -2967 4379 -2933
rect 4437 -2967 4484 -2933
rect 4520 -2967 4554 -2933
rect 4590 -2967 4637 -2933
rect 4888 -2967 4935 -2933
rect 4971 -2967 5005 -2933
rect 5041 -2967 5088 -2933
rect 5214 -2934 5249 -2912
rect 9734 -2604 9781 -2570
rect 9817 -2604 9851 -2570
rect 9887 -2604 9934 -2570
rect 10186 -2604 10233 -2570
rect 10269 -2604 10303 -2570
rect 10339 -2604 10386 -2570
rect 10444 -2604 10491 -2570
rect 10527 -2604 10561 -2570
rect 10597 -2604 10644 -2570
rect 10702 -2604 10749 -2570
rect 10785 -2604 10819 -2570
rect 10855 -2604 10902 -2570
rect 10960 -2604 11007 -2570
rect 11043 -2604 11077 -2570
rect 11113 -2604 11160 -2570
rect 11412 -2604 11459 -2570
rect 11495 -2604 11529 -2570
rect 11565 -2604 11612 -2570
rect 11670 -2604 11717 -2570
rect 11753 -2604 11787 -2570
rect 11823 -2604 11870 -2570
rect 11928 -2604 11975 -2570
rect 12011 -2604 12045 -2570
rect 12081 -2604 12128 -2570
rect 12380 -2604 12427 -2570
rect 12463 -2604 12497 -2570
rect 12533 -2604 12580 -2570
rect 12638 -2604 12685 -2570
rect 12721 -2604 12755 -2570
rect 12791 -2604 12838 -2570
rect 12896 -2604 12943 -2570
rect 12979 -2604 13013 -2570
rect 13049 -2604 13096 -2570
rect 13154 -2604 13201 -2570
rect 13237 -2604 13271 -2570
rect 13307 -2604 13354 -2570
rect 13606 -2604 13653 -2570
rect 13689 -2604 13723 -2570
rect 13759 -2604 13806 -2570
rect 13931 -2572 13932 -2538
rect 18290 -2538 18324 -2536
rect 13931 -2574 13966 -2572
rect 9573 -2646 9607 -2640
rect 9573 -2718 9607 -2708
rect 9573 -2790 9607 -2776
rect 9573 -2862 9607 -2844
rect 856 -3006 890 -2980
rect 5248 -2980 5249 -2934
rect 5374 -2967 5421 -2933
rect 5457 -2967 5491 -2933
rect 5527 -2967 5574 -2933
rect 5826 -2967 5873 -2933
rect 5909 -2967 5943 -2933
rect 5979 -2967 6026 -2933
rect 6084 -2967 6131 -2933
rect 6167 -2967 6201 -2933
rect 6237 -2967 6284 -2933
rect 6342 -2967 6389 -2933
rect 6425 -2967 6459 -2933
rect 6495 -2967 6542 -2933
rect 6600 -2967 6647 -2933
rect 6683 -2967 6717 -2933
rect 6753 -2967 6800 -2933
rect 7052 -2967 7099 -2933
rect 7135 -2967 7169 -2933
rect 7205 -2967 7252 -2933
rect 7310 -2967 7357 -2933
rect 7393 -2967 7427 -2933
rect 7463 -2967 7510 -2933
rect 7568 -2967 7615 -2933
rect 7651 -2967 7685 -2933
rect 7721 -2967 7768 -2933
rect 8020 -2967 8067 -2933
rect 8103 -2967 8137 -2933
rect 8173 -2967 8220 -2933
rect 8278 -2967 8325 -2933
rect 8361 -2967 8395 -2933
rect 8431 -2967 8478 -2933
rect 8536 -2967 8583 -2933
rect 8619 -2967 8653 -2933
rect 8689 -2967 8736 -2933
rect 8794 -2967 8841 -2933
rect 8877 -2967 8911 -2933
rect 8947 -2967 8994 -2933
rect 9246 -2967 9293 -2933
rect 9329 -2967 9363 -2933
rect 9399 -2967 9446 -2933
rect 9573 -2934 9607 -2912
rect 13931 -2640 13932 -2574
rect 14092 -2604 14139 -2570
rect 14175 -2604 14209 -2570
rect 14245 -2604 14292 -2570
rect 14543 -2604 14590 -2570
rect 14626 -2604 14660 -2570
rect 14696 -2604 14743 -2570
rect 14801 -2604 14848 -2570
rect 14884 -2604 14918 -2570
rect 14954 -2604 15001 -2570
rect 15059 -2604 15106 -2570
rect 15142 -2604 15176 -2570
rect 15212 -2604 15259 -2570
rect 15317 -2604 15364 -2570
rect 15400 -2604 15434 -2570
rect 15470 -2604 15517 -2570
rect 15769 -2604 15816 -2570
rect 15852 -2604 15886 -2570
rect 15922 -2604 15969 -2570
rect 16027 -2604 16074 -2570
rect 16110 -2604 16144 -2570
rect 16180 -2604 16227 -2570
rect 16285 -2604 16332 -2570
rect 16368 -2604 16402 -2570
rect 16438 -2604 16485 -2570
rect 16737 -2604 16784 -2570
rect 16820 -2604 16854 -2570
rect 16890 -2604 16937 -2570
rect 16995 -2604 17042 -2570
rect 17078 -2604 17112 -2570
rect 17148 -2604 17195 -2570
rect 17253 -2604 17300 -2570
rect 17336 -2604 17370 -2570
rect 17406 -2604 17453 -2570
rect 17511 -2604 17558 -2570
rect 17594 -2604 17628 -2570
rect 17664 -2604 17711 -2570
rect 17963 -2604 18010 -2570
rect 18046 -2604 18080 -2570
rect 18116 -2604 18163 -2570
rect 18290 -2574 18324 -2572
rect 13931 -2646 13966 -2640
rect 13931 -2708 13932 -2646
rect 13931 -2718 13966 -2708
rect 13931 -2776 13932 -2718
rect 13931 -2790 13966 -2776
rect 13931 -2844 13932 -2790
rect 13931 -2862 13966 -2844
rect 13931 -2912 13932 -2862
rect 5214 -3006 5249 -2980
rect 856 -3078 890 -3048
rect 856 -3150 890 -3116
rect 856 -3218 890 -3184
rect 971 -3029 1005 -3010
rect 971 -3097 1005 -3095
rect 971 -3133 1005 -3131
rect 971 -3218 1005 -3199
rect 1229 -3029 1263 -3010
rect 1229 -3097 1263 -3095
rect 1229 -3133 1263 -3131
rect 1229 -3218 1263 -3199
rect 1423 -3029 1457 -3010
rect 1423 -3097 1457 -3095
rect 1423 -3133 1457 -3131
rect 1423 -3218 1457 -3199
rect 1681 -3029 1715 -3010
rect 1681 -3097 1715 -3095
rect 1681 -3133 1715 -3131
rect 1681 -3218 1715 -3199
rect 1939 -3029 1973 -3010
rect 1939 -3097 1973 -3095
rect 1939 -3133 1973 -3131
rect 1939 -3218 1973 -3199
rect 2197 -3029 2231 -3010
rect 2197 -3097 2231 -3095
rect 2197 -3133 2231 -3131
rect 2197 -3218 2231 -3199
rect 2455 -3029 2489 -3010
rect 2455 -3097 2489 -3095
rect 2455 -3133 2489 -3131
rect 2455 -3218 2489 -3199
rect 2649 -3029 2683 -3010
rect 2649 -3097 2683 -3095
rect 2649 -3133 2683 -3131
rect 2649 -3218 2683 -3199
rect 2907 -3029 2941 -3010
rect 2907 -3097 2941 -3095
rect 2907 -3133 2941 -3131
rect 2907 -3218 2941 -3199
rect 3165 -3029 3199 -3010
rect 3165 -3097 3199 -3095
rect 3165 -3133 3199 -3131
rect 3165 -3218 3199 -3199
rect 3423 -3029 3457 -3010
rect 3423 -3097 3457 -3095
rect 3423 -3133 3457 -3131
rect 3423 -3218 3457 -3199
rect 3617 -3029 3651 -3010
rect 3617 -3097 3651 -3095
rect 3617 -3133 3651 -3131
rect 3617 -3218 3651 -3199
rect 3875 -3029 3909 -3010
rect 3875 -3097 3909 -3095
rect 3875 -3133 3909 -3131
rect 3875 -3218 3909 -3199
rect 4133 -3029 4167 -3010
rect 4133 -3097 4167 -3095
rect 4133 -3133 4167 -3131
rect 4133 -3218 4167 -3199
rect 4391 -3029 4425 -3010
rect 4391 -3097 4425 -3095
rect 4391 -3133 4425 -3131
rect 4391 -3218 4425 -3199
rect 4649 -3029 4683 -3010
rect 4649 -3097 4683 -3095
rect 4649 -3133 4683 -3131
rect 4649 -3218 4683 -3199
rect 4842 -3029 4876 -3010
rect 4842 -3097 4876 -3095
rect 4842 -3133 4876 -3131
rect 4842 -3218 4876 -3199
rect 5100 -3029 5134 -3010
rect 5100 -3097 5134 -3095
rect 5100 -3133 5134 -3131
rect 5100 -3218 5134 -3199
rect 5248 -3048 5249 -3006
rect 9734 -2967 9781 -2933
rect 9817 -2967 9851 -2933
rect 9887 -2967 9934 -2933
rect 10186 -2967 10233 -2933
rect 10269 -2967 10303 -2933
rect 10339 -2967 10386 -2933
rect 10444 -2967 10491 -2933
rect 10527 -2967 10561 -2933
rect 10597 -2967 10644 -2933
rect 10702 -2967 10749 -2933
rect 10785 -2967 10819 -2933
rect 10855 -2967 10902 -2933
rect 10960 -2967 11007 -2933
rect 11043 -2967 11077 -2933
rect 11113 -2967 11160 -2933
rect 11412 -2967 11459 -2933
rect 11495 -2967 11529 -2933
rect 11565 -2967 11612 -2933
rect 11670 -2967 11717 -2933
rect 11753 -2967 11787 -2933
rect 11823 -2967 11870 -2933
rect 11928 -2967 11975 -2933
rect 12011 -2967 12045 -2933
rect 12081 -2967 12128 -2933
rect 12380 -2967 12427 -2933
rect 12463 -2967 12497 -2933
rect 12533 -2967 12580 -2933
rect 12638 -2967 12685 -2933
rect 12721 -2967 12755 -2933
rect 12791 -2967 12838 -2933
rect 12896 -2967 12943 -2933
rect 12979 -2967 13013 -2933
rect 13049 -2967 13096 -2933
rect 13154 -2967 13201 -2933
rect 13237 -2967 13271 -2933
rect 13307 -2967 13354 -2933
rect 13606 -2967 13653 -2933
rect 13689 -2967 13723 -2933
rect 13759 -2967 13806 -2933
rect 13931 -2934 13966 -2912
rect 18290 -2646 18324 -2640
rect 18290 -2718 18324 -2708
rect 18290 -2790 18324 -2776
rect 18290 -2862 18324 -2844
rect 9573 -3006 9607 -2980
rect 5214 -3078 5249 -3048
rect 5248 -3116 5249 -3078
rect 5214 -3150 5249 -3116
rect 5248 -3184 5249 -3150
rect 5214 -3218 5249 -3184
rect 5328 -3029 5362 -3010
rect 5328 -3097 5362 -3095
rect 5328 -3133 5362 -3131
rect 5328 -3218 5362 -3199
rect 5586 -3029 5620 -3010
rect 5586 -3097 5620 -3095
rect 5586 -3133 5620 -3131
rect 5586 -3218 5620 -3199
rect 5780 -3029 5814 -3010
rect 5780 -3097 5814 -3095
rect 5780 -3133 5814 -3131
rect 5780 -3218 5814 -3199
rect 6038 -3029 6072 -3010
rect 6038 -3097 6072 -3095
rect 6038 -3133 6072 -3131
rect 6038 -3218 6072 -3199
rect 6296 -3029 6330 -3010
rect 6296 -3097 6330 -3095
rect 6296 -3133 6330 -3131
rect 6296 -3218 6330 -3199
rect 6554 -3029 6588 -3010
rect 6554 -3097 6588 -3095
rect 6554 -3133 6588 -3131
rect 6554 -3218 6588 -3199
rect 6812 -3029 6846 -3010
rect 6812 -3097 6846 -3095
rect 6812 -3133 6846 -3131
rect 6812 -3218 6846 -3199
rect 7006 -3029 7040 -3010
rect 7006 -3097 7040 -3095
rect 7006 -3133 7040 -3131
rect 7006 -3218 7040 -3199
rect 7264 -3029 7298 -3010
rect 7264 -3097 7298 -3095
rect 7264 -3133 7298 -3131
rect 7264 -3218 7298 -3199
rect 7522 -3029 7556 -3010
rect 7522 -3097 7556 -3095
rect 7522 -3133 7556 -3131
rect 7522 -3218 7556 -3199
rect 7780 -3029 7814 -3010
rect 7780 -3097 7814 -3095
rect 7780 -3133 7814 -3131
rect 7780 -3218 7814 -3199
rect 7974 -3029 8008 -3010
rect 7974 -3097 8008 -3095
rect 7974 -3133 8008 -3131
rect 7974 -3218 8008 -3199
rect 8232 -3029 8266 -3010
rect 8232 -3097 8266 -3095
rect 8232 -3133 8266 -3131
rect 8232 -3218 8266 -3199
rect 8490 -3029 8524 -3010
rect 8490 -3097 8524 -3095
rect 8490 -3133 8524 -3131
rect 8490 -3218 8524 -3199
rect 8748 -3029 8782 -3010
rect 8748 -3097 8782 -3095
rect 8748 -3133 8782 -3131
rect 8748 -3218 8782 -3199
rect 9006 -3029 9040 -3010
rect 9006 -3097 9040 -3095
rect 9006 -3133 9040 -3131
rect 9006 -3218 9040 -3199
rect 9200 -3029 9234 -3010
rect 9200 -3097 9234 -3095
rect 9200 -3133 9234 -3131
rect 9200 -3218 9234 -3199
rect 9458 -3029 9492 -3010
rect 9458 -3097 9492 -3095
rect 9458 -3133 9492 -3131
rect 9458 -3218 9492 -3199
rect 13931 -2980 13932 -2934
rect 14092 -2967 14139 -2933
rect 14175 -2967 14209 -2933
rect 14245 -2967 14292 -2933
rect 14543 -2967 14590 -2933
rect 14626 -2967 14660 -2933
rect 14696 -2967 14743 -2933
rect 14801 -2967 14848 -2933
rect 14884 -2967 14918 -2933
rect 14954 -2967 15001 -2933
rect 15059 -2967 15106 -2933
rect 15142 -2967 15176 -2933
rect 15212 -2967 15259 -2933
rect 15317 -2967 15364 -2933
rect 15400 -2967 15434 -2933
rect 15470 -2967 15517 -2933
rect 15769 -2967 15816 -2933
rect 15852 -2967 15886 -2933
rect 15922 -2967 15969 -2933
rect 16027 -2967 16074 -2933
rect 16110 -2967 16144 -2933
rect 16180 -2967 16227 -2933
rect 16285 -2967 16332 -2933
rect 16368 -2967 16402 -2933
rect 16438 -2967 16485 -2933
rect 16737 -2967 16784 -2933
rect 16820 -2967 16854 -2933
rect 16890 -2967 16937 -2933
rect 16995 -2967 17042 -2933
rect 17078 -2967 17112 -2933
rect 17148 -2967 17195 -2933
rect 17253 -2967 17300 -2933
rect 17336 -2967 17370 -2933
rect 17406 -2967 17453 -2933
rect 17511 -2967 17558 -2933
rect 17594 -2967 17628 -2933
rect 17664 -2967 17711 -2933
rect 17963 -2967 18010 -2933
rect 18046 -2967 18080 -2933
rect 18116 -2967 18163 -2933
rect 18290 -2934 18324 -2912
rect 13931 -3006 13966 -2980
rect 9573 -3078 9607 -3048
rect 9573 -3150 9607 -3116
rect 9573 -3218 9607 -3184
rect 9688 -3029 9722 -3010
rect 9688 -3097 9722 -3095
rect 9688 -3133 9722 -3131
rect 9688 -3218 9722 -3199
rect 9946 -3029 9980 -3010
rect 9946 -3097 9980 -3095
rect 9946 -3133 9980 -3131
rect 9946 -3218 9980 -3199
rect 10140 -3029 10174 -3010
rect 10140 -3097 10174 -3095
rect 10140 -3133 10174 -3131
rect 10140 -3218 10174 -3199
rect 10398 -3029 10432 -3010
rect 10398 -3097 10432 -3095
rect 10398 -3133 10432 -3131
rect 10398 -3218 10432 -3199
rect 10656 -3029 10690 -3010
rect 10656 -3097 10690 -3095
rect 10656 -3133 10690 -3131
rect 10656 -3218 10690 -3199
rect 10914 -3029 10948 -3010
rect 10914 -3097 10948 -3095
rect 10914 -3133 10948 -3131
rect 10914 -3218 10948 -3199
rect 11172 -3029 11206 -3010
rect 11172 -3097 11206 -3095
rect 11172 -3133 11206 -3131
rect 11172 -3218 11206 -3199
rect 11366 -3029 11400 -3010
rect 11366 -3097 11400 -3095
rect 11366 -3133 11400 -3131
rect 11366 -3218 11400 -3199
rect 11624 -3029 11658 -3010
rect 11624 -3097 11658 -3095
rect 11624 -3133 11658 -3131
rect 11624 -3218 11658 -3199
rect 11882 -3029 11916 -3010
rect 11882 -3097 11916 -3095
rect 11882 -3133 11916 -3131
rect 11882 -3218 11916 -3199
rect 12140 -3029 12174 -3010
rect 12140 -3097 12174 -3095
rect 12140 -3133 12174 -3131
rect 12140 -3218 12174 -3199
rect 12334 -3029 12368 -3010
rect 12334 -3097 12368 -3095
rect 12334 -3133 12368 -3131
rect 12334 -3218 12368 -3199
rect 12592 -3029 12626 -3010
rect 12592 -3097 12626 -3095
rect 12592 -3133 12626 -3131
rect 12592 -3218 12626 -3199
rect 12850 -3029 12884 -3010
rect 12850 -3097 12884 -3095
rect 12850 -3133 12884 -3131
rect 12850 -3218 12884 -3199
rect 13108 -3029 13142 -3010
rect 13108 -3097 13142 -3095
rect 13108 -3133 13142 -3131
rect 13108 -3218 13142 -3199
rect 13366 -3029 13400 -3010
rect 13366 -3097 13400 -3095
rect 13366 -3133 13400 -3131
rect 13366 -3218 13400 -3199
rect 13560 -3029 13594 -3010
rect 13560 -3097 13594 -3095
rect 13560 -3133 13594 -3131
rect 13560 -3218 13594 -3199
rect 13818 -3029 13852 -3010
rect 13818 -3097 13852 -3095
rect 13818 -3133 13852 -3131
rect 13818 -3218 13852 -3199
rect 13931 -3048 13932 -3006
rect 18290 -3006 18324 -2980
rect 13931 -3078 13966 -3048
rect 13931 -3116 13932 -3078
rect 13931 -3150 13966 -3116
rect 13931 -3184 13932 -3150
rect 13931 -3218 13966 -3184
rect 14046 -3029 14080 -3010
rect 14046 -3097 14080 -3095
rect 14046 -3133 14080 -3131
rect 14046 -3218 14080 -3199
rect 14304 -3029 14338 -3010
rect 14304 -3097 14338 -3095
rect 14304 -3133 14338 -3131
rect 14304 -3218 14338 -3199
rect 14497 -3029 14531 -3010
rect 14497 -3097 14531 -3095
rect 14497 -3133 14531 -3131
rect 14497 -3218 14531 -3199
rect 14755 -3029 14789 -3010
rect 14755 -3097 14789 -3095
rect 14755 -3133 14789 -3131
rect 14755 -3218 14789 -3199
rect 15013 -3029 15047 -3010
rect 15013 -3097 15047 -3095
rect 15013 -3133 15047 -3131
rect 15013 -3218 15047 -3199
rect 15271 -3029 15305 -3010
rect 15271 -3097 15305 -3095
rect 15271 -3133 15305 -3131
rect 15271 -3218 15305 -3199
rect 15529 -3029 15563 -3010
rect 15529 -3097 15563 -3095
rect 15529 -3133 15563 -3131
rect 15529 -3218 15563 -3199
rect 15723 -3029 15757 -3010
rect 15723 -3097 15757 -3095
rect 15723 -3133 15757 -3131
rect 15723 -3218 15757 -3199
rect 15981 -3029 16015 -3010
rect 15981 -3097 16015 -3095
rect 15981 -3133 16015 -3131
rect 15981 -3218 16015 -3199
rect 16239 -3029 16273 -3010
rect 16239 -3097 16273 -3095
rect 16239 -3133 16273 -3131
rect 16239 -3218 16273 -3199
rect 16497 -3029 16531 -3010
rect 16497 -3097 16531 -3095
rect 16497 -3133 16531 -3131
rect 16497 -3218 16531 -3199
rect 16691 -3029 16725 -3010
rect 16691 -3097 16725 -3095
rect 16691 -3133 16725 -3131
rect 16691 -3218 16725 -3199
rect 16949 -3029 16983 -3010
rect 16949 -3097 16983 -3095
rect 16949 -3133 16983 -3131
rect 16949 -3218 16983 -3199
rect 17207 -3029 17241 -3010
rect 17207 -3097 17241 -3095
rect 17207 -3133 17241 -3131
rect 17207 -3218 17241 -3199
rect 17465 -3029 17499 -3010
rect 17465 -3097 17499 -3095
rect 17465 -3133 17499 -3131
rect 17465 -3218 17499 -3199
rect 17723 -3029 17757 -3010
rect 17723 -3097 17757 -3095
rect 17723 -3133 17757 -3131
rect 17723 -3218 17757 -3199
rect 17917 -3029 17951 -3010
rect 17917 -3097 17951 -3095
rect 17917 -3133 17951 -3131
rect 17917 -3218 17951 -3199
rect 18175 -3029 18209 -3010
rect 18175 -3097 18209 -3095
rect 18175 -3133 18209 -3131
rect 18175 -3218 18209 -3199
rect 18290 -3078 18324 -3048
rect 18290 -3150 18324 -3116
rect 18290 -3218 18324 -3184
rect 856 -3286 890 -3256
rect 856 -3354 890 -3328
rect 856 -3422 890 -3400
rect 856 -3490 890 -3472
rect 856 -3558 890 -3544
rect 5248 -3256 5249 -3218
rect 5214 -3286 5249 -3256
rect 5248 -3328 5249 -3286
rect 5214 -3354 5249 -3328
rect 5248 -3400 5249 -3354
rect 5214 -3422 5249 -3400
rect 5248 -3472 5249 -3422
rect 5214 -3490 5249 -3472
rect 5248 -3544 5249 -3490
rect 5214 -3558 5249 -3544
rect 5248 -3592 5249 -3558
rect 9573 -3286 9607 -3256
rect 9573 -3354 9607 -3328
rect 9573 -3422 9607 -3400
rect 9573 -3490 9607 -3472
rect 9573 -3558 9607 -3544
rect 13931 -3256 13932 -3218
rect 13931 -3286 13966 -3256
rect 13931 -3328 13932 -3286
rect 13931 -3354 13966 -3328
rect 13931 -3400 13932 -3354
rect 13931 -3422 13966 -3400
rect 13931 -3472 13932 -3422
rect 13931 -3490 13966 -3472
rect 13931 -3544 13932 -3490
rect 13931 -3558 13966 -3544
rect 13931 -3592 13932 -3558
rect 18290 -3286 18324 -3256
rect 18290 -3354 18324 -3328
rect 18290 -3422 18324 -3400
rect 18290 -3490 18324 -3472
rect 18290 -3558 18324 -3544
rect 890 -3616 977 -3592
rect 856 -3626 977 -3616
rect 1011 -3626 1045 -3592
rect 1079 -3626 1113 -3592
rect 1147 -3626 1181 -3592
rect 1215 -3626 1249 -3592
rect 1283 -3626 1317 -3592
rect 1351 -3626 1385 -3592
rect 1419 -3626 1453 -3592
rect 1487 -3626 1521 -3592
rect 1555 -3626 1589 -3592
rect 1623 -3626 1657 -3592
rect 1691 -3626 1725 -3592
rect 1759 -3626 1793 -3592
rect 1827 -3626 1861 -3592
rect 1895 -3626 1929 -3592
rect 1963 -3626 1997 -3592
rect 2031 -3626 2065 -3592
rect 2099 -3626 2133 -3592
rect 2167 -3626 2201 -3592
rect 2235 -3626 2269 -3592
rect 2303 -3626 2337 -3592
rect 2371 -3626 2405 -3592
rect 2439 -3626 2473 -3592
rect 2507 -3626 2541 -3592
rect 2575 -3626 2609 -3592
rect 2643 -3626 2677 -3592
rect 2711 -3626 2745 -3592
rect 2779 -3626 2813 -3592
rect 2847 -3626 2881 -3592
rect 2915 -3626 2949 -3592
rect 2983 -3626 3017 -3592
rect 3051 -3626 3085 -3592
rect 3119 -3626 3153 -3592
rect 3187 -3626 3221 -3592
rect 3255 -3626 3289 -3592
rect 3323 -3626 3357 -3592
rect 3391 -3626 3425 -3592
rect 3459 -3626 3493 -3592
rect 3527 -3626 3561 -3592
rect 3595 -3626 3629 -3592
rect 3663 -3626 3697 -3592
rect 3731 -3626 3765 -3592
rect 3799 -3626 3833 -3592
rect 3867 -3626 3901 -3592
rect 3935 -3626 3969 -3592
rect 4003 -3626 4037 -3592
rect 4071 -3626 4105 -3592
rect 4139 -3626 4173 -3592
rect 4207 -3626 4241 -3592
rect 4275 -3626 4309 -3592
rect 4343 -3626 4377 -3592
rect 4411 -3626 4445 -3592
rect 4479 -3626 4513 -3592
rect 4547 -3626 4581 -3592
rect 4615 -3626 4649 -3592
rect 4683 -3626 4717 -3592
rect 4751 -3626 4785 -3592
rect 4819 -3626 4853 -3592
rect 4887 -3626 4921 -3592
rect 4955 -3626 4989 -3592
rect 5023 -3626 5057 -3592
rect 5091 -3616 5214 -3592
rect 5248 -3616 5372 -3592
rect 5091 -3626 5372 -3616
rect 5406 -3626 5440 -3592
rect 5474 -3626 5508 -3592
rect 5542 -3626 5576 -3592
rect 5610 -3626 5644 -3592
rect 5678 -3626 5712 -3592
rect 5746 -3626 5780 -3592
rect 5814 -3626 5848 -3592
rect 5882 -3626 5916 -3592
rect 5950 -3626 5984 -3592
rect 6018 -3626 6052 -3592
rect 6086 -3626 6120 -3592
rect 6154 -3626 6188 -3592
rect 6222 -3626 6256 -3592
rect 6290 -3626 6324 -3592
rect 6358 -3626 6392 -3592
rect 6426 -3626 6460 -3592
rect 6494 -3626 6528 -3592
rect 6562 -3626 6596 -3592
rect 6630 -3626 6664 -3592
rect 6698 -3626 6732 -3592
rect 6766 -3626 6800 -3592
rect 6834 -3626 6868 -3592
rect 6902 -3626 6936 -3592
rect 6970 -3626 7004 -3592
rect 7038 -3626 7072 -3592
rect 7106 -3626 7140 -3592
rect 7174 -3626 7208 -3592
rect 7242 -3626 7276 -3592
rect 7310 -3626 7344 -3592
rect 7378 -3626 7412 -3592
rect 7446 -3626 7480 -3592
rect 7514 -3626 7548 -3592
rect 7582 -3626 7616 -3592
rect 7650 -3626 7684 -3592
rect 7718 -3626 7752 -3592
rect 7786 -3626 7820 -3592
rect 7854 -3626 7888 -3592
rect 7922 -3626 7956 -3592
rect 7990 -3626 8024 -3592
rect 8058 -3626 8092 -3592
rect 8126 -3626 8160 -3592
rect 8194 -3626 8228 -3592
rect 8262 -3626 8296 -3592
rect 8330 -3626 8364 -3592
rect 8398 -3626 8432 -3592
rect 8466 -3626 8500 -3592
rect 8534 -3626 8568 -3592
rect 8602 -3626 8636 -3592
rect 8670 -3626 8704 -3592
rect 8738 -3626 8772 -3592
rect 8806 -3626 8840 -3592
rect 8874 -3626 8908 -3592
rect 8942 -3626 8976 -3592
rect 9010 -3626 9044 -3592
rect 9078 -3626 9112 -3592
rect 9146 -3626 9180 -3592
rect 9214 -3626 9248 -3592
rect 9282 -3626 9316 -3592
rect 9350 -3626 9384 -3592
rect 9418 -3626 9452 -3592
rect 9486 -3616 9573 -3592
rect 9607 -3616 9694 -3592
rect 9486 -3626 9694 -3616
rect 9728 -3626 9762 -3592
rect 9796 -3626 9830 -3592
rect 9864 -3626 9898 -3592
rect 9932 -3626 9966 -3592
rect 10000 -3626 10034 -3592
rect 10068 -3626 10102 -3592
rect 10136 -3626 10170 -3592
rect 10204 -3626 10238 -3592
rect 10272 -3626 10306 -3592
rect 10340 -3626 10374 -3592
rect 10408 -3626 10442 -3592
rect 10476 -3626 10510 -3592
rect 10544 -3626 10578 -3592
rect 10612 -3626 10646 -3592
rect 10680 -3626 10714 -3592
rect 10748 -3626 10782 -3592
rect 10816 -3626 10850 -3592
rect 10884 -3626 10918 -3592
rect 10952 -3626 10986 -3592
rect 11020 -3626 11054 -3592
rect 11088 -3626 11122 -3592
rect 11156 -3626 11190 -3592
rect 11224 -3626 11258 -3592
rect 11292 -3626 11326 -3592
rect 11360 -3626 11394 -3592
rect 11428 -3626 11462 -3592
rect 11496 -3626 11530 -3592
rect 11564 -3626 11598 -3592
rect 11632 -3626 11666 -3592
rect 11700 -3626 11734 -3592
rect 11768 -3626 11802 -3592
rect 11836 -3626 11870 -3592
rect 11904 -3626 11938 -3592
rect 11972 -3626 12006 -3592
rect 12040 -3626 12074 -3592
rect 12108 -3626 12142 -3592
rect 12176 -3626 12210 -3592
rect 12244 -3626 12278 -3592
rect 12312 -3626 12346 -3592
rect 12380 -3626 12414 -3592
rect 12448 -3626 12482 -3592
rect 12516 -3626 12550 -3592
rect 12584 -3626 12618 -3592
rect 12652 -3626 12686 -3592
rect 12720 -3626 12754 -3592
rect 12788 -3626 12822 -3592
rect 12856 -3626 12890 -3592
rect 12924 -3626 12958 -3592
rect 12992 -3626 13026 -3592
rect 13060 -3626 13094 -3592
rect 13128 -3626 13162 -3592
rect 13196 -3626 13230 -3592
rect 13264 -3626 13298 -3592
rect 13332 -3626 13366 -3592
rect 13400 -3626 13434 -3592
rect 13468 -3626 13502 -3592
rect 13536 -3626 13570 -3592
rect 13604 -3626 13638 -3592
rect 13672 -3626 13706 -3592
rect 13740 -3626 13774 -3592
rect 13808 -3616 13932 -3592
rect 13966 -3616 14089 -3592
rect 13808 -3626 14089 -3616
rect 14123 -3626 14157 -3592
rect 14191 -3626 14225 -3592
rect 14259 -3626 14293 -3592
rect 14327 -3626 14361 -3592
rect 14395 -3626 14429 -3592
rect 14463 -3626 14497 -3592
rect 14531 -3626 14565 -3592
rect 14599 -3626 14633 -3592
rect 14667 -3626 14701 -3592
rect 14735 -3626 14769 -3592
rect 14803 -3626 14837 -3592
rect 14871 -3626 14905 -3592
rect 14939 -3626 14973 -3592
rect 15007 -3626 15041 -3592
rect 15075 -3626 15109 -3592
rect 15143 -3626 15177 -3592
rect 15211 -3626 15245 -3592
rect 15279 -3626 15313 -3592
rect 15347 -3626 15381 -3592
rect 15415 -3626 15449 -3592
rect 15483 -3626 15517 -3592
rect 15551 -3626 15585 -3592
rect 15619 -3626 15653 -3592
rect 15687 -3626 15721 -3592
rect 15755 -3626 15789 -3592
rect 15823 -3626 15857 -3592
rect 15891 -3626 15925 -3592
rect 15959 -3626 15993 -3592
rect 16027 -3626 16061 -3592
rect 16095 -3626 16129 -3592
rect 16163 -3626 16197 -3592
rect 16231 -3626 16265 -3592
rect 16299 -3626 16333 -3592
rect 16367 -3626 16401 -3592
rect 16435 -3626 16469 -3592
rect 16503 -3626 16537 -3592
rect 16571 -3626 16605 -3592
rect 16639 -3626 16673 -3592
rect 16707 -3626 16741 -3592
rect 16775 -3626 16809 -3592
rect 16843 -3626 16877 -3592
rect 16911 -3626 16945 -3592
rect 16979 -3626 17013 -3592
rect 17047 -3626 17081 -3592
rect 17115 -3626 17149 -3592
rect 17183 -3626 17217 -3592
rect 17251 -3626 17285 -3592
rect 17319 -3626 17353 -3592
rect 17387 -3626 17421 -3592
rect 17455 -3626 17489 -3592
rect 17523 -3626 17557 -3592
rect 17591 -3626 17625 -3592
rect 17659 -3626 17693 -3592
rect 17727 -3626 17761 -3592
rect 17795 -3626 17829 -3592
rect 17863 -3626 17897 -3592
rect 17931 -3626 17965 -3592
rect 17999 -3626 18033 -3592
rect 18067 -3626 18101 -3592
rect 18135 -3626 18169 -3592
rect 18203 -3616 18290 -3592
rect 18203 -3626 18324 -3616
rect 856 -3694 890 -3688
rect 856 -3762 890 -3760
rect 856 -3798 890 -3796
rect 856 -3870 890 -3864
rect 856 -3942 890 -3932
rect 5248 -3688 5249 -3626
rect 5214 -3694 5249 -3688
rect 5248 -3760 5249 -3694
rect 5214 -3762 5249 -3760
rect 5248 -3796 5249 -3762
rect 5214 -3798 5249 -3796
rect 5248 -3864 5249 -3798
rect 5214 -3870 5249 -3864
rect 5248 -3932 5249 -3870
rect 5214 -3942 5249 -3932
rect 5248 -4000 5249 -3942
rect 9573 -3694 9607 -3688
rect 9573 -3762 9607 -3760
rect 9573 -3798 9607 -3796
rect 9573 -3870 9607 -3864
rect 9573 -3942 9607 -3932
rect 13931 -3688 13932 -3626
rect 13931 -3694 13966 -3688
rect 13931 -3760 13932 -3694
rect 13931 -3762 13966 -3760
rect 13931 -3796 13932 -3762
rect 13931 -3798 13966 -3796
rect 13931 -3864 13932 -3798
rect 13931 -3870 13966 -3864
rect 13931 -3932 13932 -3870
rect 13931 -3942 13966 -3932
rect 13931 -4000 13932 -3942
rect 18290 -3694 18324 -3688
rect 18290 -3762 18324 -3760
rect 18290 -3798 18324 -3796
rect 18290 -3870 18324 -3864
rect 18290 -3942 18324 -3932
rect 856 -4014 890 -4000
rect 856 -4086 890 -4068
rect 856 -4158 890 -4136
rect 856 -4230 890 -4192
rect 971 -4019 1005 -4000
rect 971 -4087 1005 -4085
rect 971 -4123 1005 -4121
rect 971 -4208 1005 -4189
rect 1229 -4019 1263 -4000
rect 1229 -4087 1263 -4085
rect 1229 -4123 1263 -4121
rect 1229 -4208 1263 -4189
rect 1423 -4019 1457 -4000
rect 1423 -4087 1457 -4085
rect 1423 -4123 1457 -4121
rect 1423 -4208 1457 -4189
rect 1681 -4019 1715 -4000
rect 1681 -4087 1715 -4085
rect 1681 -4123 1715 -4121
rect 1681 -4208 1715 -4189
rect 1939 -4019 1973 -4000
rect 1939 -4087 1973 -4085
rect 1939 -4123 1973 -4121
rect 1939 -4208 1973 -4189
rect 2197 -4019 2231 -4000
rect 2197 -4087 2231 -4085
rect 2197 -4123 2231 -4121
rect 2197 -4208 2231 -4189
rect 2455 -4019 2489 -4000
rect 2455 -4087 2489 -4085
rect 2455 -4123 2489 -4121
rect 2455 -4208 2489 -4189
rect 2649 -4019 2683 -4000
rect 2649 -4087 2683 -4085
rect 2649 -4123 2683 -4121
rect 2649 -4208 2683 -4189
rect 2907 -4019 2941 -4000
rect 2907 -4087 2941 -4085
rect 2907 -4123 2941 -4121
rect 2907 -4208 2941 -4189
rect 3165 -4019 3199 -4000
rect 3165 -4087 3199 -4085
rect 3165 -4123 3199 -4121
rect 3165 -4208 3199 -4189
rect 3423 -4019 3457 -4000
rect 3423 -4087 3457 -4085
rect 3423 -4123 3457 -4121
rect 3423 -4208 3457 -4189
rect 3617 -4019 3651 -4000
rect 3617 -4087 3651 -4085
rect 3617 -4123 3651 -4121
rect 3617 -4208 3651 -4189
rect 3875 -4019 3909 -4000
rect 3875 -4087 3909 -4085
rect 3875 -4123 3909 -4121
rect 3875 -4208 3909 -4189
rect 4133 -4019 4167 -4000
rect 4133 -4087 4167 -4085
rect 4133 -4123 4167 -4121
rect 4133 -4208 4167 -4189
rect 4391 -4019 4425 -4000
rect 4391 -4087 4425 -4085
rect 4391 -4123 4425 -4121
rect 4391 -4208 4425 -4189
rect 4649 -4019 4683 -4000
rect 4649 -4087 4683 -4085
rect 4649 -4123 4683 -4121
rect 4649 -4208 4683 -4189
rect 4842 -4019 4876 -4000
rect 4842 -4087 4876 -4085
rect 4842 -4123 4876 -4121
rect 4842 -4208 4876 -4189
rect 5100 -4019 5134 -4000
rect 5100 -4087 5134 -4085
rect 5100 -4123 5134 -4121
rect 5100 -4208 5134 -4189
rect 5214 -4014 5249 -4000
rect 5248 -4068 5249 -4014
rect 5214 -4086 5249 -4068
rect 5248 -4136 5249 -4086
rect 5214 -4158 5249 -4136
rect 5248 -4192 5249 -4158
rect 5214 -4230 5249 -4192
rect 5328 -4019 5362 -4000
rect 5328 -4087 5362 -4085
rect 5328 -4123 5362 -4121
rect 5328 -4208 5362 -4189
rect 5586 -4019 5620 -4000
rect 5586 -4087 5620 -4085
rect 5586 -4123 5620 -4121
rect 5586 -4208 5620 -4189
rect 5780 -4019 5814 -4000
rect 5780 -4087 5814 -4085
rect 5780 -4123 5814 -4121
rect 5780 -4208 5814 -4189
rect 6038 -4019 6072 -4000
rect 6038 -4087 6072 -4085
rect 6038 -4123 6072 -4121
rect 6038 -4208 6072 -4189
rect 6296 -4019 6330 -4000
rect 6296 -4087 6330 -4085
rect 6296 -4123 6330 -4121
rect 6296 -4208 6330 -4189
rect 6554 -4019 6588 -4000
rect 6554 -4087 6588 -4085
rect 6554 -4123 6588 -4121
rect 6554 -4208 6588 -4189
rect 6812 -4019 6846 -4000
rect 6812 -4087 6846 -4085
rect 6812 -4123 6846 -4121
rect 6812 -4208 6846 -4189
rect 7006 -4019 7040 -4000
rect 7006 -4087 7040 -4085
rect 7006 -4123 7040 -4121
rect 7006 -4208 7040 -4189
rect 7264 -4019 7298 -4000
rect 7264 -4087 7298 -4085
rect 7264 -4123 7298 -4121
rect 7264 -4208 7298 -4189
rect 7522 -4019 7556 -4000
rect 7522 -4087 7556 -4085
rect 7522 -4123 7556 -4121
rect 7522 -4208 7556 -4189
rect 7780 -4019 7814 -4000
rect 7780 -4087 7814 -4085
rect 7780 -4123 7814 -4121
rect 7780 -4208 7814 -4189
rect 7974 -4019 8008 -4000
rect 7974 -4087 8008 -4085
rect 7974 -4123 8008 -4121
rect 7974 -4208 8008 -4189
rect 8232 -4019 8266 -4000
rect 8232 -4087 8266 -4085
rect 8232 -4123 8266 -4121
rect 8232 -4208 8266 -4189
rect 8490 -4019 8524 -4000
rect 8490 -4087 8524 -4085
rect 8490 -4123 8524 -4121
rect 8490 -4208 8524 -4189
rect 8748 -4019 8782 -4000
rect 8748 -4087 8782 -4085
rect 8748 -4123 8782 -4121
rect 8748 -4208 8782 -4189
rect 9006 -4019 9040 -4000
rect 9006 -4087 9040 -4085
rect 9006 -4123 9040 -4121
rect 9006 -4208 9040 -4189
rect 9200 -4019 9234 -4000
rect 9200 -4087 9234 -4085
rect 9200 -4123 9234 -4121
rect 9200 -4208 9234 -4189
rect 9458 -4019 9492 -4000
rect 9458 -4087 9492 -4085
rect 9458 -4123 9492 -4121
rect 9458 -4208 9492 -4189
rect 9573 -4014 9607 -4000
rect 9573 -4086 9607 -4068
rect 9573 -4158 9607 -4136
rect 856 -4302 890 -4264
rect 1017 -4285 1064 -4251
rect 1100 -4285 1134 -4251
rect 1170 -4285 1217 -4251
rect 1469 -4285 1516 -4251
rect 1552 -4285 1586 -4251
rect 1622 -4285 1669 -4251
rect 1727 -4285 1774 -4251
rect 1810 -4285 1844 -4251
rect 1880 -4285 1927 -4251
rect 1985 -4285 2032 -4251
rect 2068 -4285 2102 -4251
rect 2138 -4285 2185 -4251
rect 2243 -4285 2290 -4251
rect 2326 -4285 2360 -4251
rect 2396 -4285 2443 -4251
rect 2695 -4285 2742 -4251
rect 2778 -4285 2812 -4251
rect 2848 -4285 2895 -4251
rect 2953 -4285 3000 -4251
rect 3036 -4285 3070 -4251
rect 3106 -4285 3153 -4251
rect 3211 -4285 3258 -4251
rect 3294 -4285 3328 -4251
rect 3364 -4285 3411 -4251
rect 3663 -4285 3710 -4251
rect 3746 -4285 3780 -4251
rect 3816 -4285 3863 -4251
rect 3921 -4285 3968 -4251
rect 4004 -4285 4038 -4251
rect 4074 -4285 4121 -4251
rect 4179 -4285 4226 -4251
rect 4262 -4285 4296 -4251
rect 4332 -4285 4379 -4251
rect 4437 -4285 4484 -4251
rect 4520 -4285 4554 -4251
rect 4590 -4285 4637 -4251
rect 4888 -4285 4935 -4251
rect 4971 -4285 5005 -4251
rect 5041 -4285 5088 -4251
rect 5248 -4264 5249 -4230
rect 9573 -4230 9607 -4192
rect 9688 -4019 9722 -4000
rect 9688 -4087 9722 -4085
rect 9688 -4123 9722 -4121
rect 9688 -4208 9722 -4189
rect 9946 -4019 9980 -4000
rect 9946 -4087 9980 -4085
rect 9946 -4123 9980 -4121
rect 9946 -4208 9980 -4189
rect 10140 -4019 10174 -4000
rect 10140 -4087 10174 -4085
rect 10140 -4123 10174 -4121
rect 10140 -4208 10174 -4189
rect 10398 -4019 10432 -4000
rect 10398 -4087 10432 -4085
rect 10398 -4123 10432 -4121
rect 10398 -4208 10432 -4189
rect 10656 -4019 10690 -4000
rect 10656 -4087 10690 -4085
rect 10656 -4123 10690 -4121
rect 10656 -4208 10690 -4189
rect 10914 -4019 10948 -4000
rect 10914 -4087 10948 -4085
rect 10914 -4123 10948 -4121
rect 10914 -4208 10948 -4189
rect 11172 -4019 11206 -4000
rect 11172 -4087 11206 -4085
rect 11172 -4123 11206 -4121
rect 11172 -4208 11206 -4189
rect 11366 -4019 11400 -4000
rect 11366 -4087 11400 -4085
rect 11366 -4123 11400 -4121
rect 11366 -4208 11400 -4189
rect 11624 -4019 11658 -4000
rect 11624 -4087 11658 -4085
rect 11624 -4123 11658 -4121
rect 11624 -4208 11658 -4189
rect 11882 -4019 11916 -4000
rect 11882 -4087 11916 -4085
rect 11882 -4123 11916 -4121
rect 11882 -4208 11916 -4189
rect 12140 -4019 12174 -4000
rect 12140 -4087 12174 -4085
rect 12140 -4123 12174 -4121
rect 12140 -4208 12174 -4189
rect 12334 -4019 12368 -4000
rect 12334 -4087 12368 -4085
rect 12334 -4123 12368 -4121
rect 12334 -4208 12368 -4189
rect 12592 -4019 12626 -4000
rect 12592 -4087 12626 -4085
rect 12592 -4123 12626 -4121
rect 12592 -4208 12626 -4189
rect 12850 -4019 12884 -4000
rect 12850 -4087 12884 -4085
rect 12850 -4123 12884 -4121
rect 12850 -4208 12884 -4189
rect 13108 -4019 13142 -4000
rect 13108 -4087 13142 -4085
rect 13108 -4123 13142 -4121
rect 13108 -4208 13142 -4189
rect 13366 -4019 13400 -4000
rect 13366 -4087 13400 -4085
rect 13366 -4123 13400 -4121
rect 13366 -4208 13400 -4189
rect 13560 -4019 13594 -4000
rect 13560 -4087 13594 -4085
rect 13560 -4123 13594 -4121
rect 13560 -4208 13594 -4189
rect 13818 -4019 13852 -4000
rect 13818 -4087 13852 -4085
rect 13818 -4123 13852 -4121
rect 13818 -4208 13852 -4189
rect 13931 -4014 13966 -4000
rect 13931 -4068 13932 -4014
rect 13931 -4086 13966 -4068
rect 13931 -4136 13932 -4086
rect 13931 -4158 13966 -4136
rect 13931 -4192 13932 -4158
rect 856 -4365 890 -4336
rect 5214 -4302 5249 -4264
rect 5374 -4285 5421 -4251
rect 5457 -4285 5491 -4251
rect 5527 -4285 5574 -4251
rect 5826 -4285 5873 -4251
rect 5909 -4285 5943 -4251
rect 5979 -4285 6026 -4251
rect 6084 -4285 6131 -4251
rect 6167 -4285 6201 -4251
rect 6237 -4285 6284 -4251
rect 6342 -4285 6389 -4251
rect 6425 -4285 6459 -4251
rect 6495 -4285 6542 -4251
rect 6600 -4285 6647 -4251
rect 6683 -4285 6717 -4251
rect 6753 -4285 6800 -4251
rect 7052 -4285 7099 -4251
rect 7135 -4285 7169 -4251
rect 7205 -4285 7252 -4251
rect 7310 -4285 7357 -4251
rect 7393 -4285 7427 -4251
rect 7463 -4285 7510 -4251
rect 7568 -4285 7615 -4251
rect 7651 -4285 7685 -4251
rect 7721 -4285 7768 -4251
rect 8020 -4285 8067 -4251
rect 8103 -4285 8137 -4251
rect 8173 -4285 8220 -4251
rect 8278 -4285 8325 -4251
rect 8361 -4285 8395 -4251
rect 8431 -4285 8478 -4251
rect 8536 -4285 8583 -4251
rect 8619 -4285 8653 -4251
rect 8689 -4285 8736 -4251
rect 8794 -4285 8841 -4251
rect 8877 -4285 8911 -4251
rect 8947 -4285 8994 -4251
rect 9246 -4285 9293 -4251
rect 9329 -4285 9363 -4251
rect 9399 -4285 9446 -4251
rect 13931 -4230 13966 -4192
rect 14046 -4019 14080 -4000
rect 14046 -4087 14080 -4085
rect 14046 -4123 14080 -4121
rect 14046 -4208 14080 -4189
rect 14304 -4019 14338 -4000
rect 14304 -4087 14338 -4085
rect 14304 -4123 14338 -4121
rect 14304 -4208 14338 -4189
rect 14497 -4019 14531 -4000
rect 14497 -4087 14531 -4085
rect 14497 -4123 14531 -4121
rect 14497 -4208 14531 -4189
rect 14755 -4019 14789 -4000
rect 14755 -4087 14789 -4085
rect 14755 -4123 14789 -4121
rect 14755 -4208 14789 -4189
rect 15013 -4019 15047 -4000
rect 15013 -4087 15047 -4085
rect 15013 -4123 15047 -4121
rect 15013 -4208 15047 -4189
rect 15271 -4019 15305 -4000
rect 15271 -4087 15305 -4085
rect 15271 -4123 15305 -4121
rect 15271 -4208 15305 -4189
rect 15529 -4019 15563 -4000
rect 15529 -4087 15563 -4085
rect 15529 -4123 15563 -4121
rect 15529 -4208 15563 -4189
rect 15723 -4019 15757 -4000
rect 15723 -4087 15757 -4085
rect 15723 -4123 15757 -4121
rect 15723 -4208 15757 -4189
rect 15981 -4019 16015 -4000
rect 15981 -4087 16015 -4085
rect 15981 -4123 16015 -4121
rect 15981 -4208 16015 -4189
rect 16239 -4019 16273 -4000
rect 16239 -4087 16273 -4085
rect 16239 -4123 16273 -4121
rect 16239 -4208 16273 -4189
rect 16497 -4019 16531 -4000
rect 16497 -4087 16531 -4085
rect 16497 -4123 16531 -4121
rect 16497 -4208 16531 -4189
rect 16691 -4019 16725 -4000
rect 16691 -4087 16725 -4085
rect 16691 -4123 16725 -4121
rect 16691 -4208 16725 -4189
rect 16949 -4019 16983 -4000
rect 16949 -4087 16983 -4085
rect 16949 -4123 16983 -4121
rect 16949 -4208 16983 -4189
rect 17207 -4019 17241 -4000
rect 17207 -4087 17241 -4085
rect 17207 -4123 17241 -4121
rect 17207 -4208 17241 -4189
rect 17465 -4019 17499 -4000
rect 17465 -4087 17499 -4085
rect 17465 -4123 17499 -4121
rect 17465 -4208 17499 -4189
rect 17723 -4019 17757 -4000
rect 17723 -4087 17757 -4085
rect 17723 -4123 17757 -4121
rect 17723 -4208 17757 -4189
rect 17917 -4019 17951 -4000
rect 17917 -4087 17951 -4085
rect 17917 -4123 17951 -4121
rect 17917 -4208 17951 -4189
rect 18175 -4019 18209 -4000
rect 18175 -4087 18209 -4085
rect 18175 -4123 18209 -4121
rect 18175 -4208 18209 -4189
rect 18290 -4014 18324 -4000
rect 18290 -4086 18324 -4068
rect 18290 -4158 18324 -4136
rect 5248 -4336 5249 -4302
rect 5214 -4365 5249 -4336
rect 9573 -4302 9607 -4264
rect 9734 -4285 9781 -4251
rect 9817 -4285 9851 -4251
rect 9887 -4285 9934 -4251
rect 10186 -4285 10233 -4251
rect 10269 -4285 10303 -4251
rect 10339 -4285 10386 -4251
rect 10444 -4285 10491 -4251
rect 10527 -4285 10561 -4251
rect 10597 -4285 10644 -4251
rect 10702 -4285 10749 -4251
rect 10785 -4285 10819 -4251
rect 10855 -4285 10902 -4251
rect 10960 -4285 11007 -4251
rect 11043 -4285 11077 -4251
rect 11113 -4285 11160 -4251
rect 11412 -4285 11459 -4251
rect 11495 -4285 11529 -4251
rect 11565 -4285 11612 -4251
rect 11670 -4285 11717 -4251
rect 11753 -4285 11787 -4251
rect 11823 -4285 11870 -4251
rect 11928 -4285 11975 -4251
rect 12011 -4285 12045 -4251
rect 12081 -4285 12128 -4251
rect 12380 -4285 12427 -4251
rect 12463 -4285 12497 -4251
rect 12533 -4285 12580 -4251
rect 12638 -4285 12685 -4251
rect 12721 -4285 12755 -4251
rect 12791 -4285 12838 -4251
rect 12896 -4285 12943 -4251
rect 12979 -4285 13013 -4251
rect 13049 -4285 13096 -4251
rect 13154 -4285 13201 -4251
rect 13237 -4285 13271 -4251
rect 13307 -4285 13354 -4251
rect 13606 -4285 13653 -4251
rect 13689 -4285 13723 -4251
rect 13759 -4285 13806 -4251
rect 13931 -4264 13932 -4230
rect 18290 -4230 18324 -4192
rect 9573 -4365 9607 -4336
rect 13931 -4302 13966 -4264
rect 14092 -4285 14139 -4251
rect 14175 -4285 14209 -4251
rect 14245 -4285 14292 -4251
rect 14543 -4285 14590 -4251
rect 14626 -4285 14660 -4251
rect 14696 -4285 14743 -4251
rect 14801 -4285 14848 -4251
rect 14884 -4285 14918 -4251
rect 14954 -4285 15001 -4251
rect 15059 -4285 15106 -4251
rect 15142 -4285 15176 -4251
rect 15212 -4285 15259 -4251
rect 15317 -4285 15364 -4251
rect 15400 -4285 15434 -4251
rect 15470 -4285 15517 -4251
rect 15769 -4285 15816 -4251
rect 15852 -4285 15886 -4251
rect 15922 -4285 15969 -4251
rect 16027 -4285 16074 -4251
rect 16110 -4285 16144 -4251
rect 16180 -4285 16227 -4251
rect 16285 -4285 16332 -4251
rect 16368 -4285 16402 -4251
rect 16438 -4285 16485 -4251
rect 16737 -4285 16784 -4251
rect 16820 -4285 16854 -4251
rect 16890 -4285 16937 -4251
rect 16995 -4285 17042 -4251
rect 17078 -4285 17112 -4251
rect 17148 -4285 17195 -4251
rect 17253 -4285 17300 -4251
rect 17336 -4285 17370 -4251
rect 17406 -4285 17453 -4251
rect 17511 -4285 17558 -4251
rect 17594 -4285 17628 -4251
rect 17664 -4285 17711 -4251
rect 17963 -4285 18010 -4251
rect 18046 -4285 18080 -4251
rect 18116 -4285 18163 -4251
rect 13931 -4336 13932 -4302
rect 13931 -4365 13966 -4336
rect 18290 -4302 18324 -4264
rect 18290 -4365 18324 -4336
rect 856 -4399 930 -4365
rect 964 -4399 977 -4365
rect 1036 -4399 1045 -4365
rect 1108 -4399 1113 -4365
rect 1180 -4399 1181 -4365
rect 1215 -4399 1218 -4365
rect 1283 -4399 1290 -4365
rect 1351 -4399 1362 -4365
rect 1419 -4399 1434 -4365
rect 1487 -4399 1506 -4365
rect 1555 -4399 1578 -4365
rect 1623 -4399 1650 -4365
rect 1691 -4399 1722 -4365
rect 1759 -4399 1793 -4365
rect 1828 -4399 1861 -4365
rect 1900 -4399 1929 -4365
rect 1972 -4399 1997 -4365
rect 2044 -4399 2065 -4365
rect 2116 -4399 2133 -4365
rect 2188 -4399 2201 -4365
rect 2260 -4399 2269 -4365
rect 2332 -4399 2337 -4365
rect 2404 -4399 2405 -4365
rect 2439 -4399 2442 -4365
rect 2507 -4399 2514 -4365
rect 2575 -4399 2586 -4365
rect 2643 -4399 2658 -4365
rect 2711 -4399 2730 -4365
rect 2779 -4399 2802 -4365
rect 2847 -4399 2874 -4365
rect 2915 -4399 2946 -4365
rect 2983 -4399 3017 -4365
rect 3052 -4399 3085 -4365
rect 3124 -4399 3153 -4365
rect 3196 -4399 3221 -4365
rect 3268 -4399 3289 -4365
rect 3340 -4399 3357 -4365
rect 3412 -4399 3425 -4365
rect 3484 -4399 3493 -4365
rect 3556 -4399 3561 -4365
rect 3628 -4399 3629 -4365
rect 3663 -4399 3666 -4365
rect 3731 -4399 3738 -4365
rect 3799 -4399 3810 -4365
rect 3867 -4399 3882 -4365
rect 3935 -4399 3954 -4365
rect 4003 -4399 4026 -4365
rect 4071 -4399 4098 -4365
rect 4139 -4399 4170 -4365
rect 4207 -4399 4241 -4365
rect 4276 -4399 4309 -4365
rect 4348 -4399 4377 -4365
rect 4420 -4399 4445 -4365
rect 4492 -4399 4513 -4365
rect 4564 -4399 4581 -4365
rect 4636 -4399 4649 -4365
rect 4708 -4399 4717 -4365
rect 4780 -4399 4785 -4365
rect 4852 -4399 4853 -4365
rect 4887 -4399 4890 -4365
rect 4955 -4399 4962 -4365
rect 5023 -4399 5034 -4365
rect 5091 -4399 5106 -4365
rect 5140 -4399 5323 -4365
rect 5357 -4399 5372 -4365
rect 5429 -4399 5440 -4365
rect 5501 -4399 5508 -4365
rect 5573 -4399 5576 -4365
rect 5610 -4399 5611 -4365
rect 5678 -4399 5683 -4365
rect 5746 -4399 5755 -4365
rect 5814 -4399 5827 -4365
rect 5882 -4399 5899 -4365
rect 5950 -4399 5971 -4365
rect 6018 -4399 6043 -4365
rect 6086 -4399 6115 -4365
rect 6154 -4399 6187 -4365
rect 6222 -4399 6256 -4365
rect 6293 -4399 6324 -4365
rect 6365 -4399 6392 -4365
rect 6437 -4399 6460 -4365
rect 6509 -4399 6528 -4365
rect 6581 -4399 6596 -4365
rect 6653 -4399 6664 -4365
rect 6725 -4399 6732 -4365
rect 6797 -4399 6800 -4365
rect 6834 -4399 6835 -4365
rect 6902 -4399 6907 -4365
rect 6970 -4399 6979 -4365
rect 7038 -4399 7051 -4365
rect 7106 -4399 7123 -4365
rect 7174 -4399 7195 -4365
rect 7242 -4399 7267 -4365
rect 7310 -4399 7339 -4365
rect 7378 -4399 7411 -4365
rect 7446 -4399 7480 -4365
rect 7517 -4399 7548 -4365
rect 7589 -4399 7616 -4365
rect 7661 -4399 7684 -4365
rect 7733 -4399 7752 -4365
rect 7805 -4399 7820 -4365
rect 7877 -4399 7888 -4365
rect 7949 -4399 7956 -4365
rect 8021 -4399 8024 -4365
rect 8058 -4399 8059 -4365
rect 8126 -4399 8131 -4365
rect 8194 -4399 8203 -4365
rect 8262 -4399 8275 -4365
rect 8330 -4399 8347 -4365
rect 8398 -4399 8419 -4365
rect 8466 -4399 8491 -4365
rect 8534 -4399 8563 -4365
rect 8602 -4399 8635 -4365
rect 8670 -4399 8704 -4365
rect 8741 -4399 8772 -4365
rect 8813 -4399 8840 -4365
rect 8885 -4399 8908 -4365
rect 8957 -4399 8976 -4365
rect 9029 -4399 9044 -4365
rect 9101 -4399 9112 -4365
rect 9173 -4399 9180 -4365
rect 9245 -4399 9248 -4365
rect 9282 -4399 9283 -4365
rect 9350 -4399 9355 -4365
rect 9418 -4399 9427 -4365
rect 9486 -4399 9499 -4365
rect 9533 -4399 9647 -4365
rect 9681 -4399 9694 -4365
rect 9753 -4399 9762 -4365
rect 9825 -4399 9830 -4365
rect 9897 -4399 9898 -4365
rect 9932 -4399 9935 -4365
rect 10000 -4399 10007 -4365
rect 10068 -4399 10079 -4365
rect 10136 -4399 10151 -4365
rect 10204 -4399 10223 -4365
rect 10272 -4399 10295 -4365
rect 10340 -4399 10367 -4365
rect 10408 -4399 10439 -4365
rect 10476 -4399 10510 -4365
rect 10545 -4399 10578 -4365
rect 10617 -4399 10646 -4365
rect 10689 -4399 10714 -4365
rect 10761 -4399 10782 -4365
rect 10833 -4399 10850 -4365
rect 10905 -4399 10918 -4365
rect 10977 -4399 10986 -4365
rect 11049 -4399 11054 -4365
rect 11121 -4399 11122 -4365
rect 11156 -4399 11159 -4365
rect 11224 -4399 11231 -4365
rect 11292 -4399 11303 -4365
rect 11360 -4399 11375 -4365
rect 11428 -4399 11447 -4365
rect 11496 -4399 11519 -4365
rect 11564 -4399 11591 -4365
rect 11632 -4399 11663 -4365
rect 11700 -4399 11734 -4365
rect 11769 -4399 11802 -4365
rect 11841 -4399 11870 -4365
rect 11913 -4399 11938 -4365
rect 11985 -4399 12006 -4365
rect 12057 -4399 12074 -4365
rect 12129 -4399 12142 -4365
rect 12201 -4399 12210 -4365
rect 12273 -4399 12278 -4365
rect 12345 -4399 12346 -4365
rect 12380 -4399 12383 -4365
rect 12448 -4399 12455 -4365
rect 12516 -4399 12527 -4365
rect 12584 -4399 12599 -4365
rect 12652 -4399 12671 -4365
rect 12720 -4399 12743 -4365
rect 12788 -4399 12815 -4365
rect 12856 -4399 12887 -4365
rect 12924 -4399 12958 -4365
rect 12993 -4399 13026 -4365
rect 13065 -4399 13094 -4365
rect 13137 -4399 13162 -4365
rect 13209 -4399 13230 -4365
rect 13281 -4399 13298 -4365
rect 13353 -4399 13366 -4365
rect 13425 -4399 13434 -4365
rect 13497 -4399 13502 -4365
rect 13569 -4399 13570 -4365
rect 13604 -4399 13607 -4365
rect 13672 -4399 13679 -4365
rect 13740 -4399 13751 -4365
rect 13808 -4399 13823 -4365
rect 13857 -4399 14040 -4365
rect 14074 -4399 14089 -4365
rect 14146 -4399 14157 -4365
rect 14218 -4399 14225 -4365
rect 14290 -4399 14293 -4365
rect 14327 -4399 14328 -4365
rect 14395 -4399 14400 -4365
rect 14463 -4399 14472 -4365
rect 14531 -4399 14544 -4365
rect 14599 -4399 14616 -4365
rect 14667 -4399 14688 -4365
rect 14735 -4399 14760 -4365
rect 14803 -4399 14832 -4365
rect 14871 -4399 14904 -4365
rect 14939 -4399 14973 -4365
rect 15010 -4399 15041 -4365
rect 15082 -4399 15109 -4365
rect 15154 -4399 15177 -4365
rect 15226 -4399 15245 -4365
rect 15298 -4399 15313 -4365
rect 15370 -4399 15381 -4365
rect 15442 -4399 15449 -4365
rect 15514 -4399 15517 -4365
rect 15551 -4399 15552 -4365
rect 15619 -4399 15624 -4365
rect 15687 -4399 15696 -4365
rect 15755 -4399 15768 -4365
rect 15823 -4399 15840 -4365
rect 15891 -4399 15912 -4365
rect 15959 -4399 15984 -4365
rect 16027 -4399 16056 -4365
rect 16095 -4399 16128 -4365
rect 16163 -4399 16197 -4365
rect 16234 -4399 16265 -4365
rect 16306 -4399 16333 -4365
rect 16378 -4399 16401 -4365
rect 16450 -4399 16469 -4365
rect 16522 -4399 16537 -4365
rect 16594 -4399 16605 -4365
rect 16666 -4399 16673 -4365
rect 16738 -4399 16741 -4365
rect 16775 -4399 16776 -4365
rect 16843 -4399 16848 -4365
rect 16911 -4399 16920 -4365
rect 16979 -4399 16992 -4365
rect 17047 -4399 17064 -4365
rect 17115 -4399 17136 -4365
rect 17183 -4399 17208 -4365
rect 17251 -4399 17280 -4365
rect 17319 -4399 17352 -4365
rect 17387 -4399 17421 -4365
rect 17458 -4399 17489 -4365
rect 17530 -4399 17557 -4365
rect 17602 -4399 17625 -4365
rect 17674 -4399 17693 -4365
rect 17746 -4399 17761 -4365
rect 17818 -4399 17829 -4365
rect 17890 -4399 17897 -4365
rect 17962 -4399 17965 -4365
rect 17999 -4399 18000 -4365
rect 18067 -4399 18072 -4365
rect 18135 -4399 18144 -4365
rect 18203 -4399 18216 -4365
rect 18250 -4399 18324 -4365
rect 856 -4428 890 -4399
rect 856 -4500 890 -4462
rect 5214 -4428 5249 -4399
rect 5248 -4462 5249 -4428
rect 1017 -4513 1064 -4479
rect 1100 -4513 1134 -4479
rect 1170 -4513 1217 -4479
rect 1469 -4513 1516 -4479
rect 1552 -4513 1586 -4479
rect 1622 -4513 1669 -4479
rect 1727 -4513 1774 -4479
rect 1810 -4513 1844 -4479
rect 1880 -4513 1927 -4479
rect 1985 -4513 2032 -4479
rect 2068 -4513 2102 -4479
rect 2138 -4513 2185 -4479
rect 2243 -4513 2290 -4479
rect 2326 -4513 2360 -4479
rect 2396 -4513 2443 -4479
rect 2695 -4513 2742 -4479
rect 2778 -4513 2812 -4479
rect 2848 -4513 2895 -4479
rect 2953 -4513 3000 -4479
rect 3036 -4513 3070 -4479
rect 3106 -4513 3153 -4479
rect 3211 -4513 3258 -4479
rect 3294 -4513 3328 -4479
rect 3364 -4513 3411 -4479
rect 3663 -4513 3710 -4479
rect 3746 -4513 3780 -4479
rect 3816 -4513 3863 -4479
rect 3921 -4513 3968 -4479
rect 4004 -4513 4038 -4479
rect 4074 -4513 4121 -4479
rect 4179 -4513 4226 -4479
rect 4262 -4513 4296 -4479
rect 4332 -4513 4379 -4479
rect 4437 -4513 4484 -4479
rect 4520 -4513 4554 -4479
rect 4590 -4513 4637 -4479
rect 4888 -4513 4935 -4479
rect 4971 -4513 5005 -4479
rect 5041 -4513 5088 -4479
rect 5214 -4500 5249 -4462
rect 9573 -4428 9607 -4399
rect 856 -4572 890 -4534
rect 5248 -4534 5249 -4500
rect 5374 -4513 5421 -4479
rect 5457 -4513 5491 -4479
rect 5527 -4513 5574 -4479
rect 5826 -4513 5873 -4479
rect 5909 -4513 5943 -4479
rect 5979 -4513 6026 -4479
rect 6084 -4513 6131 -4479
rect 6167 -4513 6201 -4479
rect 6237 -4513 6284 -4479
rect 6342 -4513 6389 -4479
rect 6425 -4513 6459 -4479
rect 6495 -4513 6542 -4479
rect 6600 -4513 6647 -4479
rect 6683 -4513 6717 -4479
rect 6753 -4513 6800 -4479
rect 7052 -4513 7099 -4479
rect 7135 -4513 7169 -4479
rect 7205 -4513 7252 -4479
rect 7310 -4513 7357 -4479
rect 7393 -4513 7427 -4479
rect 7463 -4513 7510 -4479
rect 7568 -4513 7615 -4479
rect 7651 -4513 7685 -4479
rect 7721 -4513 7768 -4479
rect 8020 -4513 8067 -4479
rect 8103 -4513 8137 -4479
rect 8173 -4513 8220 -4479
rect 8278 -4513 8325 -4479
rect 8361 -4513 8395 -4479
rect 8431 -4513 8478 -4479
rect 8536 -4513 8583 -4479
rect 8619 -4513 8653 -4479
rect 8689 -4513 8736 -4479
rect 8794 -4513 8841 -4479
rect 8877 -4513 8911 -4479
rect 8947 -4513 8994 -4479
rect 9246 -4513 9293 -4479
rect 9329 -4513 9363 -4479
rect 9399 -4513 9446 -4479
rect 9573 -4500 9607 -4462
rect 13931 -4428 13966 -4399
rect 13931 -4462 13932 -4428
rect 856 -4628 890 -4606
rect 856 -4696 890 -4678
rect 856 -4764 890 -4750
rect 971 -4575 1005 -4556
rect 971 -4643 1005 -4641
rect 971 -4679 1005 -4677
rect 971 -4764 1005 -4745
rect 1229 -4575 1263 -4556
rect 1229 -4643 1263 -4641
rect 1229 -4679 1263 -4677
rect 1229 -4764 1263 -4745
rect 1423 -4575 1457 -4556
rect 1423 -4643 1457 -4641
rect 1423 -4679 1457 -4677
rect 1423 -4764 1457 -4745
rect 1681 -4575 1715 -4556
rect 1681 -4643 1715 -4641
rect 1681 -4679 1715 -4677
rect 1681 -4764 1715 -4745
rect 1939 -4575 1973 -4556
rect 1939 -4643 1973 -4641
rect 1939 -4679 1973 -4677
rect 1939 -4764 1973 -4745
rect 2197 -4575 2231 -4556
rect 2197 -4643 2231 -4641
rect 2197 -4679 2231 -4677
rect 2197 -4764 2231 -4745
rect 2455 -4575 2489 -4556
rect 2455 -4643 2489 -4641
rect 2455 -4679 2489 -4677
rect 2455 -4764 2489 -4745
rect 2649 -4575 2683 -4556
rect 2649 -4643 2683 -4641
rect 2649 -4679 2683 -4677
rect 2649 -4764 2683 -4745
rect 2907 -4575 2941 -4556
rect 2907 -4643 2941 -4641
rect 2907 -4679 2941 -4677
rect 2907 -4764 2941 -4745
rect 3165 -4575 3199 -4556
rect 3165 -4643 3199 -4641
rect 3165 -4679 3199 -4677
rect 3165 -4764 3199 -4745
rect 3423 -4575 3457 -4556
rect 3423 -4643 3457 -4641
rect 3423 -4679 3457 -4677
rect 3423 -4764 3457 -4745
rect 3617 -4575 3651 -4556
rect 3617 -4643 3651 -4641
rect 3617 -4679 3651 -4677
rect 3617 -4764 3651 -4745
rect 3875 -4575 3909 -4556
rect 3875 -4643 3909 -4641
rect 3875 -4679 3909 -4677
rect 3875 -4764 3909 -4745
rect 4133 -4575 4167 -4556
rect 4133 -4643 4167 -4641
rect 4133 -4679 4167 -4677
rect 4133 -4764 4167 -4745
rect 4391 -4575 4425 -4556
rect 4391 -4643 4425 -4641
rect 4391 -4679 4425 -4677
rect 4391 -4764 4425 -4745
rect 4649 -4575 4683 -4556
rect 4649 -4643 4683 -4641
rect 4649 -4679 4683 -4677
rect 4649 -4764 4683 -4745
rect 4842 -4575 4876 -4556
rect 4842 -4643 4876 -4641
rect 4842 -4679 4876 -4677
rect 4842 -4764 4876 -4745
rect 5100 -4575 5134 -4556
rect 5100 -4643 5134 -4641
rect 5100 -4679 5134 -4677
rect 5100 -4764 5134 -4745
rect 5214 -4572 5249 -4534
rect 9734 -4513 9781 -4479
rect 9817 -4513 9851 -4479
rect 9887 -4513 9934 -4479
rect 10186 -4513 10233 -4479
rect 10269 -4513 10303 -4479
rect 10339 -4513 10386 -4479
rect 10444 -4513 10491 -4479
rect 10527 -4513 10561 -4479
rect 10597 -4513 10644 -4479
rect 10702 -4513 10749 -4479
rect 10785 -4513 10819 -4479
rect 10855 -4513 10902 -4479
rect 10960 -4513 11007 -4479
rect 11043 -4513 11077 -4479
rect 11113 -4513 11160 -4479
rect 11412 -4513 11459 -4479
rect 11495 -4513 11529 -4479
rect 11565 -4513 11612 -4479
rect 11670 -4513 11717 -4479
rect 11753 -4513 11787 -4479
rect 11823 -4513 11870 -4479
rect 11928 -4513 11975 -4479
rect 12011 -4513 12045 -4479
rect 12081 -4513 12128 -4479
rect 12380 -4513 12427 -4479
rect 12463 -4513 12497 -4479
rect 12533 -4513 12580 -4479
rect 12638 -4513 12685 -4479
rect 12721 -4513 12755 -4479
rect 12791 -4513 12838 -4479
rect 12896 -4513 12943 -4479
rect 12979 -4513 13013 -4479
rect 13049 -4513 13096 -4479
rect 13154 -4513 13201 -4479
rect 13237 -4513 13271 -4479
rect 13307 -4513 13354 -4479
rect 13606 -4513 13653 -4479
rect 13689 -4513 13723 -4479
rect 13759 -4513 13806 -4479
rect 13931 -4500 13966 -4462
rect 18290 -4428 18324 -4399
rect 5248 -4606 5249 -4572
rect 5214 -4628 5249 -4606
rect 5248 -4678 5249 -4628
rect 5214 -4696 5249 -4678
rect 5248 -4750 5249 -4696
rect 5214 -4764 5249 -4750
rect 5328 -4575 5362 -4556
rect 5328 -4643 5362 -4641
rect 5328 -4679 5362 -4677
rect 5328 -4764 5362 -4745
rect 5586 -4575 5620 -4556
rect 5586 -4643 5620 -4641
rect 5586 -4679 5620 -4677
rect 5586 -4764 5620 -4745
rect 5780 -4575 5814 -4556
rect 5780 -4643 5814 -4641
rect 5780 -4679 5814 -4677
rect 5780 -4764 5814 -4745
rect 6038 -4575 6072 -4556
rect 6038 -4643 6072 -4641
rect 6038 -4679 6072 -4677
rect 6038 -4764 6072 -4745
rect 6296 -4575 6330 -4556
rect 6296 -4643 6330 -4641
rect 6296 -4679 6330 -4677
rect 6296 -4764 6330 -4745
rect 6554 -4575 6588 -4556
rect 6554 -4643 6588 -4641
rect 6554 -4679 6588 -4677
rect 6554 -4764 6588 -4745
rect 6812 -4575 6846 -4556
rect 6812 -4643 6846 -4641
rect 6812 -4679 6846 -4677
rect 6812 -4764 6846 -4745
rect 7006 -4575 7040 -4556
rect 7006 -4643 7040 -4641
rect 7006 -4679 7040 -4677
rect 7006 -4764 7040 -4745
rect 7264 -4575 7298 -4556
rect 7264 -4643 7298 -4641
rect 7264 -4679 7298 -4677
rect 7264 -4764 7298 -4745
rect 7522 -4575 7556 -4556
rect 7522 -4643 7556 -4641
rect 7522 -4679 7556 -4677
rect 7522 -4764 7556 -4745
rect 7780 -4575 7814 -4556
rect 7780 -4643 7814 -4641
rect 7780 -4679 7814 -4677
rect 7780 -4764 7814 -4745
rect 7974 -4575 8008 -4556
rect 7974 -4643 8008 -4641
rect 7974 -4679 8008 -4677
rect 7974 -4764 8008 -4745
rect 8232 -4575 8266 -4556
rect 8232 -4643 8266 -4641
rect 8232 -4679 8266 -4677
rect 8232 -4764 8266 -4745
rect 8490 -4575 8524 -4556
rect 8490 -4643 8524 -4641
rect 8490 -4679 8524 -4677
rect 8490 -4764 8524 -4745
rect 8748 -4575 8782 -4556
rect 8748 -4643 8782 -4641
rect 8748 -4679 8782 -4677
rect 8748 -4764 8782 -4745
rect 9006 -4575 9040 -4556
rect 9006 -4643 9040 -4641
rect 9006 -4679 9040 -4677
rect 9006 -4764 9040 -4745
rect 9200 -4575 9234 -4556
rect 9200 -4643 9234 -4641
rect 9200 -4679 9234 -4677
rect 9200 -4764 9234 -4745
rect 9458 -4575 9492 -4556
rect 9458 -4643 9492 -4641
rect 9458 -4679 9492 -4677
rect 9458 -4764 9492 -4745
rect 9573 -4572 9607 -4534
rect 13931 -4534 13932 -4500
rect 14092 -4513 14139 -4479
rect 14175 -4513 14209 -4479
rect 14245 -4513 14292 -4479
rect 14543 -4513 14590 -4479
rect 14626 -4513 14660 -4479
rect 14696 -4513 14743 -4479
rect 14801 -4513 14848 -4479
rect 14884 -4513 14918 -4479
rect 14954 -4513 15001 -4479
rect 15059 -4513 15106 -4479
rect 15142 -4513 15176 -4479
rect 15212 -4513 15259 -4479
rect 15317 -4513 15364 -4479
rect 15400 -4513 15434 -4479
rect 15470 -4513 15517 -4479
rect 15769 -4513 15816 -4479
rect 15852 -4513 15886 -4479
rect 15922 -4513 15969 -4479
rect 16027 -4513 16074 -4479
rect 16110 -4513 16144 -4479
rect 16180 -4513 16227 -4479
rect 16285 -4513 16332 -4479
rect 16368 -4513 16402 -4479
rect 16438 -4513 16485 -4479
rect 16737 -4513 16784 -4479
rect 16820 -4513 16854 -4479
rect 16890 -4513 16937 -4479
rect 16995 -4513 17042 -4479
rect 17078 -4513 17112 -4479
rect 17148 -4513 17195 -4479
rect 17253 -4513 17300 -4479
rect 17336 -4513 17370 -4479
rect 17406 -4513 17453 -4479
rect 17511 -4513 17558 -4479
rect 17594 -4513 17628 -4479
rect 17664 -4513 17711 -4479
rect 17963 -4513 18010 -4479
rect 18046 -4513 18080 -4479
rect 18116 -4513 18163 -4479
rect 18290 -4500 18324 -4462
rect 9573 -4628 9607 -4606
rect 9573 -4696 9607 -4678
rect 9573 -4764 9607 -4750
rect 9688 -4575 9722 -4556
rect 9688 -4643 9722 -4641
rect 9688 -4679 9722 -4677
rect 9688 -4764 9722 -4745
rect 9946 -4575 9980 -4556
rect 9946 -4643 9980 -4641
rect 9946 -4679 9980 -4677
rect 9946 -4764 9980 -4745
rect 10140 -4575 10174 -4556
rect 10140 -4643 10174 -4641
rect 10140 -4679 10174 -4677
rect 10140 -4764 10174 -4745
rect 10398 -4575 10432 -4556
rect 10398 -4643 10432 -4641
rect 10398 -4679 10432 -4677
rect 10398 -4764 10432 -4745
rect 10656 -4575 10690 -4556
rect 10656 -4643 10690 -4641
rect 10656 -4679 10690 -4677
rect 10656 -4764 10690 -4745
rect 10914 -4575 10948 -4556
rect 10914 -4643 10948 -4641
rect 10914 -4679 10948 -4677
rect 10914 -4764 10948 -4745
rect 11172 -4575 11206 -4556
rect 11172 -4643 11206 -4641
rect 11172 -4679 11206 -4677
rect 11172 -4764 11206 -4745
rect 11366 -4575 11400 -4556
rect 11366 -4643 11400 -4641
rect 11366 -4679 11400 -4677
rect 11366 -4764 11400 -4745
rect 11624 -4575 11658 -4556
rect 11624 -4643 11658 -4641
rect 11624 -4679 11658 -4677
rect 11624 -4764 11658 -4745
rect 11882 -4575 11916 -4556
rect 11882 -4643 11916 -4641
rect 11882 -4679 11916 -4677
rect 11882 -4764 11916 -4745
rect 12140 -4575 12174 -4556
rect 12140 -4643 12174 -4641
rect 12140 -4679 12174 -4677
rect 12140 -4764 12174 -4745
rect 12334 -4575 12368 -4556
rect 12334 -4643 12368 -4641
rect 12334 -4679 12368 -4677
rect 12334 -4764 12368 -4745
rect 12592 -4575 12626 -4556
rect 12592 -4643 12626 -4641
rect 12592 -4679 12626 -4677
rect 12592 -4764 12626 -4745
rect 12850 -4575 12884 -4556
rect 12850 -4643 12884 -4641
rect 12850 -4679 12884 -4677
rect 12850 -4764 12884 -4745
rect 13108 -4575 13142 -4556
rect 13108 -4643 13142 -4641
rect 13108 -4679 13142 -4677
rect 13108 -4764 13142 -4745
rect 13366 -4575 13400 -4556
rect 13366 -4643 13400 -4641
rect 13366 -4679 13400 -4677
rect 13366 -4764 13400 -4745
rect 13560 -4575 13594 -4556
rect 13560 -4643 13594 -4641
rect 13560 -4679 13594 -4677
rect 13560 -4764 13594 -4745
rect 13818 -4575 13852 -4556
rect 13818 -4643 13852 -4641
rect 13818 -4679 13852 -4677
rect 13818 -4764 13852 -4745
rect 13931 -4572 13966 -4534
rect 13931 -4606 13932 -4572
rect 13931 -4628 13966 -4606
rect 13931 -4678 13932 -4628
rect 13931 -4696 13966 -4678
rect 13931 -4750 13932 -4696
rect 13931 -4764 13966 -4750
rect 14046 -4575 14080 -4556
rect 14046 -4643 14080 -4641
rect 14046 -4679 14080 -4677
rect 14046 -4764 14080 -4745
rect 14304 -4575 14338 -4556
rect 14304 -4643 14338 -4641
rect 14304 -4679 14338 -4677
rect 14304 -4764 14338 -4745
rect 14497 -4575 14531 -4556
rect 14497 -4643 14531 -4641
rect 14497 -4679 14531 -4677
rect 14497 -4764 14531 -4745
rect 14755 -4575 14789 -4556
rect 14755 -4643 14789 -4641
rect 14755 -4679 14789 -4677
rect 14755 -4764 14789 -4745
rect 15013 -4575 15047 -4556
rect 15013 -4643 15047 -4641
rect 15013 -4679 15047 -4677
rect 15013 -4764 15047 -4745
rect 15271 -4575 15305 -4556
rect 15271 -4643 15305 -4641
rect 15271 -4679 15305 -4677
rect 15271 -4764 15305 -4745
rect 15529 -4575 15563 -4556
rect 15529 -4643 15563 -4641
rect 15529 -4679 15563 -4677
rect 15529 -4764 15563 -4745
rect 15723 -4575 15757 -4556
rect 15723 -4643 15757 -4641
rect 15723 -4679 15757 -4677
rect 15723 -4764 15757 -4745
rect 15981 -4575 16015 -4556
rect 15981 -4643 16015 -4641
rect 15981 -4679 16015 -4677
rect 15981 -4764 16015 -4745
rect 16239 -4575 16273 -4556
rect 16239 -4643 16273 -4641
rect 16239 -4679 16273 -4677
rect 16239 -4764 16273 -4745
rect 16497 -4575 16531 -4556
rect 16497 -4643 16531 -4641
rect 16497 -4679 16531 -4677
rect 16497 -4764 16531 -4745
rect 16691 -4575 16725 -4556
rect 16691 -4643 16725 -4641
rect 16691 -4679 16725 -4677
rect 16691 -4764 16725 -4745
rect 16949 -4575 16983 -4556
rect 16949 -4643 16983 -4641
rect 16949 -4679 16983 -4677
rect 16949 -4764 16983 -4745
rect 17207 -4575 17241 -4556
rect 17207 -4643 17241 -4641
rect 17207 -4679 17241 -4677
rect 17207 -4764 17241 -4745
rect 17465 -4575 17499 -4556
rect 17465 -4643 17499 -4641
rect 17465 -4679 17499 -4677
rect 17465 -4764 17499 -4745
rect 17723 -4575 17757 -4556
rect 17723 -4643 17757 -4641
rect 17723 -4679 17757 -4677
rect 17723 -4764 17757 -4745
rect 17917 -4575 17951 -4556
rect 17917 -4643 17951 -4641
rect 17917 -4679 17951 -4677
rect 17917 -4764 17951 -4745
rect 18175 -4575 18209 -4556
rect 18175 -4643 18209 -4641
rect 18175 -4679 18209 -4677
rect 18175 -4764 18209 -4745
rect 18290 -4572 18324 -4534
rect 18290 -4628 18324 -4606
rect 18290 -4696 18324 -4678
rect 18290 -4764 18324 -4750
rect 856 -4832 890 -4822
rect 856 -4900 890 -4894
rect 856 -4968 890 -4966
rect 856 -5004 890 -5002
rect 856 -5076 890 -5070
rect 5248 -4822 5249 -4764
rect 5214 -4832 5249 -4822
rect 5248 -4894 5249 -4832
rect 5214 -4900 5249 -4894
rect 5248 -4966 5249 -4900
rect 5214 -4968 5249 -4966
rect 5248 -5002 5249 -4968
rect 5214 -5004 5249 -5002
rect 5248 -5070 5249 -5004
rect 5214 -5076 5249 -5070
rect 5248 -5138 5249 -5076
rect 9573 -4832 9607 -4822
rect 9573 -4900 9607 -4894
rect 9573 -4968 9607 -4966
rect 9573 -5004 9607 -5002
rect 9573 -5076 9607 -5070
rect 13931 -4822 13932 -4764
rect 13931 -4832 13966 -4822
rect 13931 -4894 13932 -4832
rect 13931 -4900 13966 -4894
rect 13931 -4966 13932 -4900
rect 13931 -4968 13966 -4966
rect 13931 -5002 13932 -4968
rect 13931 -5004 13966 -5002
rect 13931 -5070 13932 -5004
rect 13931 -5076 13966 -5070
rect 13931 -5138 13932 -5076
rect 18290 -4832 18324 -4822
rect 18290 -4900 18324 -4894
rect 18290 -4968 18324 -4966
rect 18290 -5004 18324 -5002
rect 18290 -5076 18324 -5070
rect 856 -5148 977 -5138
rect 890 -5172 977 -5148
rect 1011 -5172 1045 -5138
rect 1079 -5172 1113 -5138
rect 1147 -5172 1181 -5138
rect 1215 -5172 1249 -5138
rect 1283 -5172 1317 -5138
rect 1351 -5172 1385 -5138
rect 1419 -5172 1453 -5138
rect 1487 -5172 1521 -5138
rect 1555 -5172 1589 -5138
rect 1623 -5172 1657 -5138
rect 1691 -5172 1725 -5138
rect 1759 -5172 1793 -5138
rect 1827 -5172 1861 -5138
rect 1895 -5172 1929 -5138
rect 1963 -5172 1997 -5138
rect 2031 -5172 2065 -5138
rect 2099 -5172 2133 -5138
rect 2167 -5172 2201 -5138
rect 2235 -5172 2269 -5138
rect 2303 -5172 2337 -5138
rect 2371 -5172 2405 -5138
rect 2439 -5172 2473 -5138
rect 2507 -5172 2541 -5138
rect 2575 -5172 2609 -5138
rect 2643 -5172 2677 -5138
rect 2711 -5172 2745 -5138
rect 2779 -5172 2813 -5138
rect 2847 -5172 2881 -5138
rect 2915 -5172 2949 -5138
rect 2983 -5172 3017 -5138
rect 3051 -5172 3085 -5138
rect 3119 -5172 3153 -5138
rect 3187 -5172 3221 -5138
rect 3255 -5172 3289 -5138
rect 3323 -5172 3357 -5138
rect 3391 -5172 3425 -5138
rect 3459 -5172 3493 -5138
rect 3527 -5172 3561 -5138
rect 3595 -5172 3629 -5138
rect 3663 -5172 3697 -5138
rect 3731 -5172 3765 -5138
rect 3799 -5172 3833 -5138
rect 3867 -5172 3901 -5138
rect 3935 -5172 3969 -5138
rect 4003 -5172 4037 -5138
rect 4071 -5172 4105 -5138
rect 4139 -5172 4173 -5138
rect 4207 -5172 4241 -5138
rect 4275 -5172 4309 -5138
rect 4343 -5172 4377 -5138
rect 4411 -5172 4445 -5138
rect 4479 -5172 4513 -5138
rect 4547 -5172 4581 -5138
rect 4615 -5172 4649 -5138
rect 4683 -5172 4717 -5138
rect 4751 -5172 4785 -5138
rect 4819 -5172 4853 -5138
rect 4887 -5172 4921 -5138
rect 4955 -5172 4989 -5138
rect 5023 -5172 5057 -5138
rect 5091 -5148 5372 -5138
rect 5091 -5172 5214 -5148
rect 5248 -5172 5372 -5148
rect 5406 -5172 5440 -5138
rect 5474 -5172 5508 -5138
rect 5542 -5172 5576 -5138
rect 5610 -5172 5644 -5138
rect 5678 -5172 5712 -5138
rect 5746 -5172 5780 -5138
rect 5814 -5172 5848 -5138
rect 5882 -5172 5916 -5138
rect 5950 -5172 5984 -5138
rect 6018 -5172 6052 -5138
rect 6086 -5172 6120 -5138
rect 6154 -5172 6188 -5138
rect 6222 -5172 6256 -5138
rect 6290 -5172 6324 -5138
rect 6358 -5172 6392 -5138
rect 6426 -5172 6460 -5138
rect 6494 -5172 6528 -5138
rect 6562 -5172 6596 -5138
rect 6630 -5172 6664 -5138
rect 6698 -5172 6732 -5138
rect 6766 -5172 6800 -5138
rect 6834 -5172 6868 -5138
rect 6902 -5172 6936 -5138
rect 6970 -5172 7004 -5138
rect 7038 -5172 7072 -5138
rect 7106 -5172 7140 -5138
rect 7174 -5172 7208 -5138
rect 7242 -5172 7276 -5138
rect 7310 -5172 7344 -5138
rect 7378 -5172 7412 -5138
rect 7446 -5172 7480 -5138
rect 7514 -5172 7548 -5138
rect 7582 -5172 7616 -5138
rect 7650 -5172 7684 -5138
rect 7718 -5172 7752 -5138
rect 7786 -5172 7820 -5138
rect 7854 -5172 7888 -5138
rect 7922 -5172 7956 -5138
rect 7990 -5172 8024 -5138
rect 8058 -5172 8092 -5138
rect 8126 -5172 8160 -5138
rect 8194 -5172 8228 -5138
rect 8262 -5172 8296 -5138
rect 8330 -5172 8364 -5138
rect 8398 -5172 8432 -5138
rect 8466 -5172 8500 -5138
rect 8534 -5172 8568 -5138
rect 8602 -5172 8636 -5138
rect 8670 -5172 8704 -5138
rect 8738 -5172 8772 -5138
rect 8806 -5172 8840 -5138
rect 8874 -5172 8908 -5138
rect 8942 -5172 8976 -5138
rect 9010 -5172 9044 -5138
rect 9078 -5172 9112 -5138
rect 9146 -5172 9180 -5138
rect 9214 -5172 9248 -5138
rect 9282 -5172 9316 -5138
rect 9350 -5172 9384 -5138
rect 9418 -5172 9452 -5138
rect 9486 -5148 9694 -5138
rect 9486 -5172 9573 -5148
rect 9607 -5172 9694 -5148
rect 9728 -5172 9762 -5138
rect 9796 -5172 9830 -5138
rect 9864 -5172 9898 -5138
rect 9932 -5172 9966 -5138
rect 10000 -5172 10034 -5138
rect 10068 -5172 10102 -5138
rect 10136 -5172 10170 -5138
rect 10204 -5172 10238 -5138
rect 10272 -5172 10306 -5138
rect 10340 -5172 10374 -5138
rect 10408 -5172 10442 -5138
rect 10476 -5172 10510 -5138
rect 10544 -5172 10578 -5138
rect 10612 -5172 10646 -5138
rect 10680 -5172 10714 -5138
rect 10748 -5172 10782 -5138
rect 10816 -5172 10850 -5138
rect 10884 -5172 10918 -5138
rect 10952 -5172 10986 -5138
rect 11020 -5172 11054 -5138
rect 11088 -5172 11122 -5138
rect 11156 -5172 11190 -5138
rect 11224 -5172 11258 -5138
rect 11292 -5172 11326 -5138
rect 11360 -5172 11394 -5138
rect 11428 -5172 11462 -5138
rect 11496 -5172 11530 -5138
rect 11564 -5172 11598 -5138
rect 11632 -5172 11666 -5138
rect 11700 -5172 11734 -5138
rect 11768 -5172 11802 -5138
rect 11836 -5172 11870 -5138
rect 11904 -5172 11938 -5138
rect 11972 -5172 12006 -5138
rect 12040 -5172 12074 -5138
rect 12108 -5172 12142 -5138
rect 12176 -5172 12210 -5138
rect 12244 -5172 12278 -5138
rect 12312 -5172 12346 -5138
rect 12380 -5172 12414 -5138
rect 12448 -5172 12482 -5138
rect 12516 -5172 12550 -5138
rect 12584 -5172 12618 -5138
rect 12652 -5172 12686 -5138
rect 12720 -5172 12754 -5138
rect 12788 -5172 12822 -5138
rect 12856 -5172 12890 -5138
rect 12924 -5172 12958 -5138
rect 12992 -5172 13026 -5138
rect 13060 -5172 13094 -5138
rect 13128 -5172 13162 -5138
rect 13196 -5172 13230 -5138
rect 13264 -5172 13298 -5138
rect 13332 -5172 13366 -5138
rect 13400 -5172 13434 -5138
rect 13468 -5172 13502 -5138
rect 13536 -5172 13570 -5138
rect 13604 -5172 13638 -5138
rect 13672 -5172 13706 -5138
rect 13740 -5172 13774 -5138
rect 13808 -5148 14089 -5138
rect 13808 -5172 13932 -5148
rect 13966 -5172 14089 -5148
rect 14123 -5172 14157 -5138
rect 14191 -5172 14225 -5138
rect 14259 -5172 14293 -5138
rect 14327 -5172 14361 -5138
rect 14395 -5172 14429 -5138
rect 14463 -5172 14497 -5138
rect 14531 -5172 14565 -5138
rect 14599 -5172 14633 -5138
rect 14667 -5172 14701 -5138
rect 14735 -5172 14769 -5138
rect 14803 -5172 14837 -5138
rect 14871 -5172 14905 -5138
rect 14939 -5172 14973 -5138
rect 15007 -5172 15041 -5138
rect 15075 -5172 15109 -5138
rect 15143 -5172 15177 -5138
rect 15211 -5172 15245 -5138
rect 15279 -5172 15313 -5138
rect 15347 -5172 15381 -5138
rect 15415 -5172 15449 -5138
rect 15483 -5172 15517 -5138
rect 15551 -5172 15585 -5138
rect 15619 -5172 15653 -5138
rect 15687 -5172 15721 -5138
rect 15755 -5172 15789 -5138
rect 15823 -5172 15857 -5138
rect 15891 -5172 15925 -5138
rect 15959 -5172 15993 -5138
rect 16027 -5172 16061 -5138
rect 16095 -5172 16129 -5138
rect 16163 -5172 16197 -5138
rect 16231 -5172 16265 -5138
rect 16299 -5172 16333 -5138
rect 16367 -5172 16401 -5138
rect 16435 -5172 16469 -5138
rect 16503 -5172 16537 -5138
rect 16571 -5172 16605 -5138
rect 16639 -5172 16673 -5138
rect 16707 -5172 16741 -5138
rect 16775 -5172 16809 -5138
rect 16843 -5172 16877 -5138
rect 16911 -5172 16945 -5138
rect 16979 -5172 17013 -5138
rect 17047 -5172 17081 -5138
rect 17115 -5172 17149 -5138
rect 17183 -5172 17217 -5138
rect 17251 -5172 17285 -5138
rect 17319 -5172 17353 -5138
rect 17387 -5172 17421 -5138
rect 17455 -5172 17489 -5138
rect 17523 -5172 17557 -5138
rect 17591 -5172 17625 -5138
rect 17659 -5172 17693 -5138
rect 17727 -5172 17761 -5138
rect 17795 -5172 17829 -5138
rect 17863 -5172 17897 -5138
rect 17931 -5172 17965 -5138
rect 17999 -5172 18033 -5138
rect 18067 -5172 18101 -5138
rect 18135 -5172 18169 -5138
rect 18203 -5148 18324 -5138
rect 18203 -5172 18290 -5148
rect 856 -5220 890 -5206
rect 856 -5292 890 -5274
rect 856 -5364 890 -5342
rect 856 -5436 890 -5410
rect 856 -5508 890 -5478
rect 5248 -5206 5249 -5172
rect 5214 -5220 5249 -5206
rect 5248 -5274 5249 -5220
rect 5214 -5292 5249 -5274
rect 5248 -5342 5249 -5292
rect 5214 -5364 5249 -5342
rect 5248 -5410 5249 -5364
rect 5214 -5436 5249 -5410
rect 5248 -5478 5249 -5436
rect 5214 -5508 5249 -5478
rect 5248 -5546 5249 -5508
rect 9573 -5220 9607 -5206
rect 9573 -5292 9607 -5274
rect 9573 -5364 9607 -5342
rect 9573 -5436 9607 -5410
rect 9573 -5508 9607 -5478
rect 13931 -5206 13932 -5172
rect 13931 -5220 13966 -5206
rect 13931 -5274 13932 -5220
rect 13931 -5292 13966 -5274
rect 13931 -5342 13932 -5292
rect 13931 -5364 13966 -5342
rect 13931 -5410 13932 -5364
rect 13931 -5436 13966 -5410
rect 13931 -5478 13932 -5436
rect 13931 -5508 13966 -5478
rect 13931 -5546 13932 -5508
rect 18290 -5220 18324 -5206
rect 18290 -5292 18324 -5274
rect 18290 -5364 18324 -5342
rect 18290 -5436 18324 -5410
rect 18290 -5508 18324 -5478
rect 856 -5580 890 -5546
rect 856 -5648 890 -5614
rect 856 -5716 890 -5686
rect 971 -5565 1005 -5546
rect 971 -5633 1005 -5631
rect 971 -5669 1005 -5667
rect 971 -5754 1005 -5735
rect 1229 -5565 1263 -5546
rect 1229 -5633 1263 -5631
rect 1229 -5669 1263 -5667
rect 1229 -5754 1263 -5735
rect 1423 -5565 1457 -5546
rect 1423 -5633 1457 -5631
rect 1423 -5669 1457 -5667
rect 1423 -5754 1457 -5735
rect 1681 -5565 1715 -5546
rect 1681 -5633 1715 -5631
rect 1681 -5669 1715 -5667
rect 1681 -5754 1715 -5735
rect 1939 -5565 1973 -5546
rect 1939 -5633 1973 -5631
rect 1939 -5669 1973 -5667
rect 1939 -5754 1973 -5735
rect 2197 -5565 2231 -5546
rect 2197 -5633 2231 -5631
rect 2197 -5669 2231 -5667
rect 2197 -5754 2231 -5735
rect 2455 -5565 2489 -5546
rect 2455 -5633 2489 -5631
rect 2455 -5669 2489 -5667
rect 2455 -5754 2489 -5735
rect 2649 -5565 2683 -5546
rect 2649 -5633 2683 -5631
rect 2649 -5669 2683 -5667
rect 2649 -5754 2683 -5735
rect 2907 -5565 2941 -5546
rect 2907 -5633 2941 -5631
rect 2907 -5669 2941 -5667
rect 2907 -5754 2941 -5735
rect 3165 -5565 3199 -5546
rect 3165 -5633 3199 -5631
rect 3165 -5669 3199 -5667
rect 3165 -5754 3199 -5735
rect 3423 -5565 3457 -5546
rect 3423 -5633 3457 -5631
rect 3423 -5669 3457 -5667
rect 3423 -5754 3457 -5735
rect 3617 -5565 3651 -5546
rect 3617 -5633 3651 -5631
rect 3617 -5669 3651 -5667
rect 3617 -5754 3651 -5735
rect 3875 -5565 3909 -5546
rect 3875 -5633 3909 -5631
rect 3875 -5669 3909 -5667
rect 3875 -5754 3909 -5735
rect 4133 -5565 4167 -5546
rect 4133 -5633 4167 -5631
rect 4133 -5669 4167 -5667
rect 4133 -5754 4167 -5735
rect 4391 -5565 4425 -5546
rect 4391 -5633 4425 -5631
rect 4391 -5669 4425 -5667
rect 4391 -5754 4425 -5735
rect 4649 -5565 4683 -5546
rect 4649 -5633 4683 -5631
rect 4649 -5669 4683 -5667
rect 4649 -5754 4683 -5735
rect 4842 -5565 4876 -5546
rect 4842 -5633 4876 -5631
rect 4842 -5669 4876 -5667
rect 4842 -5754 4876 -5735
rect 5100 -5565 5134 -5546
rect 5100 -5633 5134 -5631
rect 5100 -5669 5134 -5667
rect 5100 -5754 5134 -5735
rect 5214 -5580 5249 -5546
rect 5248 -5614 5249 -5580
rect 5214 -5648 5249 -5614
rect 5248 -5686 5249 -5648
rect 5214 -5716 5249 -5686
rect 856 -5784 890 -5758
rect 5248 -5758 5249 -5716
rect 5328 -5565 5362 -5546
rect 5328 -5633 5362 -5631
rect 5328 -5669 5362 -5667
rect 5328 -5754 5362 -5735
rect 5586 -5565 5620 -5546
rect 5586 -5633 5620 -5631
rect 5586 -5669 5620 -5667
rect 5586 -5754 5620 -5735
rect 5780 -5565 5814 -5546
rect 5780 -5633 5814 -5631
rect 5780 -5669 5814 -5667
rect 5780 -5754 5814 -5735
rect 6038 -5565 6072 -5546
rect 6038 -5633 6072 -5631
rect 6038 -5669 6072 -5667
rect 6038 -5754 6072 -5735
rect 6296 -5565 6330 -5546
rect 6296 -5633 6330 -5631
rect 6296 -5669 6330 -5667
rect 6296 -5754 6330 -5735
rect 6554 -5565 6588 -5546
rect 6554 -5633 6588 -5631
rect 6554 -5669 6588 -5667
rect 6554 -5754 6588 -5735
rect 6812 -5565 6846 -5546
rect 6812 -5633 6846 -5631
rect 6812 -5669 6846 -5667
rect 6812 -5754 6846 -5735
rect 7006 -5565 7040 -5546
rect 7006 -5633 7040 -5631
rect 7006 -5669 7040 -5667
rect 7006 -5754 7040 -5735
rect 7264 -5565 7298 -5546
rect 7264 -5633 7298 -5631
rect 7264 -5669 7298 -5667
rect 7264 -5754 7298 -5735
rect 7522 -5565 7556 -5546
rect 7522 -5633 7556 -5631
rect 7522 -5669 7556 -5667
rect 7522 -5754 7556 -5735
rect 7780 -5565 7814 -5546
rect 7780 -5633 7814 -5631
rect 7780 -5669 7814 -5667
rect 7780 -5754 7814 -5735
rect 7974 -5565 8008 -5546
rect 7974 -5633 8008 -5631
rect 7974 -5669 8008 -5667
rect 7974 -5754 8008 -5735
rect 8232 -5565 8266 -5546
rect 8232 -5633 8266 -5631
rect 8232 -5669 8266 -5667
rect 8232 -5754 8266 -5735
rect 8490 -5565 8524 -5546
rect 8490 -5633 8524 -5631
rect 8490 -5669 8524 -5667
rect 8490 -5754 8524 -5735
rect 8748 -5565 8782 -5546
rect 8748 -5633 8782 -5631
rect 8748 -5669 8782 -5667
rect 8748 -5754 8782 -5735
rect 9006 -5565 9040 -5546
rect 9006 -5633 9040 -5631
rect 9006 -5669 9040 -5667
rect 9006 -5754 9040 -5735
rect 9200 -5565 9234 -5546
rect 9200 -5633 9234 -5631
rect 9200 -5669 9234 -5667
rect 9200 -5754 9234 -5735
rect 9458 -5565 9492 -5546
rect 9458 -5633 9492 -5631
rect 9458 -5669 9492 -5667
rect 9458 -5754 9492 -5735
rect 9573 -5580 9607 -5546
rect 9573 -5648 9607 -5614
rect 9573 -5716 9607 -5686
rect 5214 -5784 5249 -5758
rect 856 -5852 890 -5830
rect 1017 -5831 1064 -5797
rect 1100 -5831 1134 -5797
rect 1170 -5831 1217 -5797
rect 1469 -5831 1516 -5797
rect 1552 -5831 1586 -5797
rect 1622 -5831 1669 -5797
rect 1727 -5831 1774 -5797
rect 1810 -5831 1844 -5797
rect 1880 -5831 1927 -5797
rect 1985 -5831 2032 -5797
rect 2068 -5831 2102 -5797
rect 2138 -5831 2185 -5797
rect 2243 -5831 2290 -5797
rect 2326 -5831 2360 -5797
rect 2396 -5831 2443 -5797
rect 2695 -5831 2742 -5797
rect 2778 -5831 2812 -5797
rect 2848 -5831 2895 -5797
rect 2953 -5831 3000 -5797
rect 3036 -5831 3070 -5797
rect 3106 -5831 3153 -5797
rect 3211 -5831 3258 -5797
rect 3294 -5831 3328 -5797
rect 3364 -5831 3411 -5797
rect 3663 -5831 3710 -5797
rect 3746 -5831 3780 -5797
rect 3816 -5831 3863 -5797
rect 3921 -5831 3968 -5797
rect 4004 -5831 4038 -5797
rect 4074 -5831 4121 -5797
rect 4179 -5831 4226 -5797
rect 4262 -5831 4296 -5797
rect 4332 -5831 4379 -5797
rect 4437 -5831 4484 -5797
rect 4520 -5831 4554 -5797
rect 4590 -5831 4637 -5797
rect 4888 -5831 4935 -5797
rect 4971 -5831 5005 -5797
rect 5041 -5831 5088 -5797
rect 5248 -5830 5249 -5784
rect 9688 -5565 9722 -5546
rect 9688 -5633 9722 -5631
rect 9688 -5669 9722 -5667
rect 9688 -5754 9722 -5735
rect 9946 -5565 9980 -5546
rect 9946 -5633 9980 -5631
rect 9946 -5669 9980 -5667
rect 9946 -5754 9980 -5735
rect 10140 -5565 10174 -5546
rect 10140 -5633 10174 -5631
rect 10140 -5669 10174 -5667
rect 10140 -5754 10174 -5735
rect 10398 -5565 10432 -5546
rect 10398 -5633 10432 -5631
rect 10398 -5669 10432 -5667
rect 10398 -5754 10432 -5735
rect 10656 -5565 10690 -5546
rect 10656 -5633 10690 -5631
rect 10656 -5669 10690 -5667
rect 10656 -5754 10690 -5735
rect 10914 -5565 10948 -5546
rect 10914 -5633 10948 -5631
rect 10914 -5669 10948 -5667
rect 10914 -5754 10948 -5735
rect 11172 -5565 11206 -5546
rect 11172 -5633 11206 -5631
rect 11172 -5669 11206 -5667
rect 11172 -5754 11206 -5735
rect 11366 -5565 11400 -5546
rect 11366 -5633 11400 -5631
rect 11366 -5669 11400 -5667
rect 11366 -5754 11400 -5735
rect 11624 -5565 11658 -5546
rect 11624 -5633 11658 -5631
rect 11624 -5669 11658 -5667
rect 11624 -5754 11658 -5735
rect 11882 -5565 11916 -5546
rect 11882 -5633 11916 -5631
rect 11882 -5669 11916 -5667
rect 11882 -5754 11916 -5735
rect 12140 -5565 12174 -5546
rect 12140 -5633 12174 -5631
rect 12140 -5669 12174 -5667
rect 12140 -5754 12174 -5735
rect 12334 -5565 12368 -5546
rect 12334 -5633 12368 -5631
rect 12334 -5669 12368 -5667
rect 12334 -5754 12368 -5735
rect 12592 -5565 12626 -5546
rect 12592 -5633 12626 -5631
rect 12592 -5669 12626 -5667
rect 12592 -5754 12626 -5735
rect 12850 -5565 12884 -5546
rect 12850 -5633 12884 -5631
rect 12850 -5669 12884 -5667
rect 12850 -5754 12884 -5735
rect 13108 -5565 13142 -5546
rect 13108 -5633 13142 -5631
rect 13108 -5669 13142 -5667
rect 13108 -5754 13142 -5735
rect 13366 -5565 13400 -5546
rect 13366 -5633 13400 -5631
rect 13366 -5669 13400 -5667
rect 13366 -5754 13400 -5735
rect 13560 -5565 13594 -5546
rect 13560 -5633 13594 -5631
rect 13560 -5669 13594 -5667
rect 13560 -5754 13594 -5735
rect 13818 -5565 13852 -5546
rect 13818 -5633 13852 -5631
rect 13818 -5669 13852 -5667
rect 13818 -5754 13852 -5735
rect 13931 -5580 13966 -5546
rect 13931 -5614 13932 -5580
rect 13931 -5648 13966 -5614
rect 13931 -5686 13932 -5648
rect 13931 -5716 13966 -5686
rect 9573 -5784 9607 -5758
rect 856 -5920 890 -5902
rect 856 -5988 890 -5974
rect 856 -6056 890 -6046
rect 856 -6124 890 -6118
rect 5214 -5852 5249 -5830
rect 5374 -5831 5421 -5797
rect 5457 -5831 5491 -5797
rect 5527 -5831 5574 -5797
rect 5826 -5831 5873 -5797
rect 5909 -5831 5943 -5797
rect 5979 -5831 6026 -5797
rect 6084 -5831 6131 -5797
rect 6167 -5831 6201 -5797
rect 6237 -5831 6284 -5797
rect 6342 -5831 6389 -5797
rect 6425 -5831 6459 -5797
rect 6495 -5831 6542 -5797
rect 6600 -5831 6647 -5797
rect 6683 -5831 6717 -5797
rect 6753 -5831 6800 -5797
rect 7052 -5831 7099 -5797
rect 7135 -5831 7169 -5797
rect 7205 -5831 7252 -5797
rect 7310 -5831 7357 -5797
rect 7393 -5831 7427 -5797
rect 7463 -5831 7510 -5797
rect 7568 -5831 7615 -5797
rect 7651 -5831 7685 -5797
rect 7721 -5831 7768 -5797
rect 8020 -5831 8067 -5797
rect 8103 -5831 8137 -5797
rect 8173 -5831 8220 -5797
rect 8278 -5831 8325 -5797
rect 8361 -5831 8395 -5797
rect 8431 -5831 8478 -5797
rect 8536 -5831 8583 -5797
rect 8619 -5831 8653 -5797
rect 8689 -5831 8736 -5797
rect 8794 -5831 8841 -5797
rect 8877 -5831 8911 -5797
rect 8947 -5831 8994 -5797
rect 9246 -5831 9293 -5797
rect 9329 -5831 9363 -5797
rect 9399 -5831 9446 -5797
rect 13931 -5758 13932 -5716
rect 14046 -5565 14080 -5546
rect 14046 -5633 14080 -5631
rect 14046 -5669 14080 -5667
rect 14046 -5754 14080 -5735
rect 14304 -5565 14338 -5546
rect 14304 -5633 14338 -5631
rect 14304 -5669 14338 -5667
rect 14304 -5754 14338 -5735
rect 14497 -5565 14531 -5546
rect 14497 -5633 14531 -5631
rect 14497 -5669 14531 -5667
rect 14497 -5754 14531 -5735
rect 14755 -5565 14789 -5546
rect 14755 -5633 14789 -5631
rect 14755 -5669 14789 -5667
rect 14755 -5754 14789 -5735
rect 15013 -5565 15047 -5546
rect 15013 -5633 15047 -5631
rect 15013 -5669 15047 -5667
rect 15013 -5754 15047 -5735
rect 15271 -5565 15305 -5546
rect 15271 -5633 15305 -5631
rect 15271 -5669 15305 -5667
rect 15271 -5754 15305 -5735
rect 15529 -5565 15563 -5546
rect 15529 -5633 15563 -5631
rect 15529 -5669 15563 -5667
rect 15529 -5754 15563 -5735
rect 15723 -5565 15757 -5546
rect 15723 -5633 15757 -5631
rect 15723 -5669 15757 -5667
rect 15723 -5754 15757 -5735
rect 15981 -5565 16015 -5546
rect 15981 -5633 16015 -5631
rect 15981 -5669 16015 -5667
rect 15981 -5754 16015 -5735
rect 16239 -5565 16273 -5546
rect 16239 -5633 16273 -5631
rect 16239 -5669 16273 -5667
rect 16239 -5754 16273 -5735
rect 16497 -5565 16531 -5546
rect 16497 -5633 16531 -5631
rect 16497 -5669 16531 -5667
rect 16497 -5754 16531 -5735
rect 16691 -5565 16725 -5546
rect 16691 -5633 16725 -5631
rect 16691 -5669 16725 -5667
rect 16691 -5754 16725 -5735
rect 16949 -5565 16983 -5546
rect 16949 -5633 16983 -5631
rect 16949 -5669 16983 -5667
rect 16949 -5754 16983 -5735
rect 17207 -5565 17241 -5546
rect 17207 -5633 17241 -5631
rect 17207 -5669 17241 -5667
rect 17207 -5754 17241 -5735
rect 17465 -5565 17499 -5546
rect 17465 -5633 17499 -5631
rect 17465 -5669 17499 -5667
rect 17465 -5754 17499 -5735
rect 17723 -5565 17757 -5546
rect 17723 -5633 17757 -5631
rect 17723 -5669 17757 -5667
rect 17723 -5754 17757 -5735
rect 17917 -5565 17951 -5546
rect 17917 -5633 17951 -5631
rect 17917 -5669 17951 -5667
rect 17917 -5754 17951 -5735
rect 18175 -5565 18209 -5546
rect 18175 -5633 18209 -5631
rect 18175 -5669 18209 -5667
rect 18175 -5754 18209 -5735
rect 18290 -5580 18324 -5546
rect 18290 -5648 18324 -5614
rect 18290 -5716 18324 -5686
rect 13931 -5784 13966 -5758
rect 5248 -5902 5249 -5852
rect 5214 -5920 5249 -5902
rect 5248 -5974 5249 -5920
rect 5214 -5988 5249 -5974
rect 5248 -6046 5249 -5988
rect 5214 -6056 5249 -6046
rect 5248 -6118 5249 -6056
rect 5214 -6124 5249 -6118
rect 856 -6192 890 -6190
rect 1017 -6193 1064 -6159
rect 1100 -6193 1134 -6159
rect 1170 -6193 1217 -6159
rect 1469 -6193 1516 -6159
rect 1552 -6193 1586 -6159
rect 1622 -6193 1669 -6159
rect 1727 -6193 1774 -6159
rect 1810 -6193 1844 -6159
rect 1880 -6193 1927 -6159
rect 1985 -6193 2032 -6159
rect 2068 -6193 2102 -6159
rect 2138 -6193 2185 -6159
rect 2243 -6193 2290 -6159
rect 2326 -6193 2360 -6159
rect 2396 -6193 2443 -6159
rect 2695 -6193 2742 -6159
rect 2778 -6193 2812 -6159
rect 2848 -6193 2895 -6159
rect 2953 -6193 3000 -6159
rect 3036 -6193 3070 -6159
rect 3106 -6193 3153 -6159
rect 3211 -6193 3258 -6159
rect 3294 -6193 3328 -6159
rect 3364 -6193 3411 -6159
rect 3663 -6193 3710 -6159
rect 3746 -6193 3780 -6159
rect 3816 -6193 3863 -6159
rect 3921 -6193 3968 -6159
rect 4004 -6193 4038 -6159
rect 4074 -6193 4121 -6159
rect 4179 -6193 4226 -6159
rect 4262 -6193 4296 -6159
rect 4332 -6193 4379 -6159
rect 4437 -6193 4484 -6159
rect 4520 -6193 4554 -6159
rect 4590 -6193 4637 -6159
rect 4888 -6193 4935 -6159
rect 4971 -6193 5005 -6159
rect 5041 -6193 5088 -6159
rect 5248 -6190 5249 -6124
rect 9573 -5852 9607 -5830
rect 9734 -5831 9781 -5797
rect 9817 -5831 9851 -5797
rect 9887 -5831 9934 -5797
rect 10186 -5831 10233 -5797
rect 10269 -5831 10303 -5797
rect 10339 -5831 10386 -5797
rect 10444 -5831 10491 -5797
rect 10527 -5831 10561 -5797
rect 10597 -5831 10644 -5797
rect 10702 -5831 10749 -5797
rect 10785 -5831 10819 -5797
rect 10855 -5831 10902 -5797
rect 10960 -5831 11007 -5797
rect 11043 -5831 11077 -5797
rect 11113 -5831 11160 -5797
rect 11412 -5831 11459 -5797
rect 11495 -5831 11529 -5797
rect 11565 -5831 11612 -5797
rect 11670 -5831 11717 -5797
rect 11753 -5831 11787 -5797
rect 11823 -5831 11870 -5797
rect 11928 -5831 11975 -5797
rect 12011 -5831 12045 -5797
rect 12081 -5831 12128 -5797
rect 12380 -5831 12427 -5797
rect 12463 -5831 12497 -5797
rect 12533 -5831 12580 -5797
rect 12638 -5831 12685 -5797
rect 12721 -5831 12755 -5797
rect 12791 -5831 12838 -5797
rect 12896 -5831 12943 -5797
rect 12979 -5831 13013 -5797
rect 13049 -5831 13096 -5797
rect 13154 -5831 13201 -5797
rect 13237 -5831 13271 -5797
rect 13307 -5831 13354 -5797
rect 13606 -5831 13653 -5797
rect 13689 -5831 13723 -5797
rect 13759 -5831 13806 -5797
rect 13931 -5830 13932 -5784
rect 18290 -5784 18324 -5758
rect 9573 -5920 9607 -5902
rect 9573 -5988 9607 -5974
rect 9573 -6056 9607 -6046
rect 9573 -6124 9607 -6118
rect 5214 -6192 5249 -6190
rect 856 -6228 890 -6226
rect 5248 -6226 5249 -6192
rect 5374 -6193 5421 -6159
rect 5457 -6193 5491 -6159
rect 5527 -6193 5574 -6159
rect 5826 -6193 5873 -6159
rect 5909 -6193 5943 -6159
rect 5979 -6193 6026 -6159
rect 6084 -6193 6131 -6159
rect 6167 -6193 6201 -6159
rect 6237 -6193 6284 -6159
rect 6342 -6193 6389 -6159
rect 6425 -6193 6459 -6159
rect 6495 -6193 6542 -6159
rect 6600 -6193 6647 -6159
rect 6683 -6193 6717 -6159
rect 6753 -6193 6800 -6159
rect 7052 -6193 7099 -6159
rect 7135 -6193 7169 -6159
rect 7205 -6193 7252 -6159
rect 7310 -6193 7357 -6159
rect 7393 -6193 7427 -6159
rect 7463 -6193 7510 -6159
rect 7568 -6193 7615 -6159
rect 7651 -6193 7685 -6159
rect 7721 -6193 7768 -6159
rect 8020 -6193 8067 -6159
rect 8103 -6193 8137 -6159
rect 8173 -6193 8220 -6159
rect 8278 -6193 8325 -6159
rect 8361 -6193 8395 -6159
rect 8431 -6193 8478 -6159
rect 8536 -6193 8583 -6159
rect 8619 -6193 8653 -6159
rect 8689 -6193 8736 -6159
rect 8794 -6193 8841 -6159
rect 8877 -6193 8911 -6159
rect 8947 -6193 8994 -6159
rect 9246 -6193 9293 -6159
rect 9329 -6193 9363 -6159
rect 9399 -6193 9446 -6159
rect 13931 -5852 13966 -5830
rect 14092 -5831 14139 -5797
rect 14175 -5831 14209 -5797
rect 14245 -5831 14292 -5797
rect 14543 -5831 14590 -5797
rect 14626 -5831 14660 -5797
rect 14696 -5831 14743 -5797
rect 14801 -5831 14848 -5797
rect 14884 -5831 14918 -5797
rect 14954 -5831 15001 -5797
rect 15059 -5831 15106 -5797
rect 15142 -5831 15176 -5797
rect 15212 -5831 15259 -5797
rect 15317 -5831 15364 -5797
rect 15400 -5831 15434 -5797
rect 15470 -5831 15517 -5797
rect 15769 -5831 15816 -5797
rect 15852 -5831 15886 -5797
rect 15922 -5831 15969 -5797
rect 16027 -5831 16074 -5797
rect 16110 -5831 16144 -5797
rect 16180 -5831 16227 -5797
rect 16285 -5831 16332 -5797
rect 16368 -5831 16402 -5797
rect 16438 -5831 16485 -5797
rect 16737 -5831 16784 -5797
rect 16820 -5831 16854 -5797
rect 16890 -5831 16937 -5797
rect 16995 -5831 17042 -5797
rect 17078 -5831 17112 -5797
rect 17148 -5831 17195 -5797
rect 17253 -5831 17300 -5797
rect 17336 -5831 17370 -5797
rect 17406 -5831 17453 -5797
rect 17511 -5831 17558 -5797
rect 17594 -5831 17628 -5797
rect 17664 -5831 17711 -5797
rect 17963 -5831 18010 -5797
rect 18046 -5831 18080 -5797
rect 18116 -5831 18163 -5797
rect 13931 -5902 13932 -5852
rect 13931 -5920 13966 -5902
rect 13931 -5974 13932 -5920
rect 13931 -5988 13966 -5974
rect 13931 -6046 13932 -5988
rect 13931 -6056 13966 -6046
rect 13931 -6118 13932 -6056
rect 13931 -6124 13966 -6118
rect 9573 -6192 9607 -6190
rect 5214 -6228 5249 -6226
rect 856 -6300 890 -6294
rect 856 -6372 890 -6362
rect 856 -6444 890 -6430
rect 971 -6255 1005 -6236
rect 971 -6323 1005 -6321
rect 971 -6359 1005 -6357
rect 971 -6444 1005 -6425
rect 1229 -6255 1263 -6236
rect 1229 -6323 1263 -6321
rect 1229 -6359 1263 -6357
rect 1229 -6444 1263 -6425
rect 1423 -6255 1457 -6236
rect 1423 -6323 1457 -6321
rect 1423 -6359 1457 -6357
rect 1423 -6444 1457 -6425
rect 1681 -6255 1715 -6236
rect 1681 -6323 1715 -6321
rect 1681 -6359 1715 -6357
rect 1681 -6444 1715 -6425
rect 1939 -6255 1973 -6236
rect 1939 -6323 1973 -6321
rect 1939 -6359 1973 -6357
rect 1939 -6444 1973 -6425
rect 2197 -6255 2231 -6236
rect 2197 -6323 2231 -6321
rect 2197 -6359 2231 -6357
rect 2197 -6444 2231 -6425
rect 2455 -6255 2489 -6236
rect 2455 -6323 2489 -6321
rect 2455 -6359 2489 -6357
rect 2455 -6444 2489 -6425
rect 2649 -6255 2683 -6236
rect 2649 -6323 2683 -6321
rect 2649 -6359 2683 -6357
rect 2649 -6444 2683 -6425
rect 2907 -6255 2941 -6236
rect 2907 -6323 2941 -6321
rect 2907 -6359 2941 -6357
rect 2907 -6444 2941 -6425
rect 3165 -6255 3199 -6236
rect 3165 -6323 3199 -6321
rect 3165 -6359 3199 -6357
rect 3165 -6444 3199 -6425
rect 3423 -6255 3457 -6236
rect 3423 -6323 3457 -6321
rect 3423 -6359 3457 -6357
rect 3423 -6444 3457 -6425
rect 3617 -6255 3651 -6236
rect 3617 -6323 3651 -6321
rect 3617 -6359 3651 -6357
rect 3617 -6444 3651 -6425
rect 3875 -6255 3909 -6236
rect 3875 -6323 3909 -6321
rect 3875 -6359 3909 -6357
rect 3875 -6444 3909 -6425
rect 4133 -6255 4167 -6236
rect 4133 -6323 4167 -6321
rect 4133 -6359 4167 -6357
rect 4133 -6444 4167 -6425
rect 4391 -6255 4425 -6236
rect 4391 -6323 4425 -6321
rect 4391 -6359 4425 -6357
rect 4391 -6444 4425 -6425
rect 4649 -6255 4683 -6236
rect 4649 -6323 4683 -6321
rect 4649 -6359 4683 -6357
rect 4649 -6444 4683 -6425
rect 4842 -6255 4876 -6236
rect 4842 -6323 4876 -6321
rect 4842 -6359 4876 -6357
rect 4842 -6444 4876 -6425
rect 5100 -6255 5134 -6236
rect 5100 -6323 5134 -6321
rect 5100 -6359 5134 -6357
rect 5100 -6444 5134 -6425
rect 5248 -6294 5249 -6228
rect 9734 -6193 9781 -6159
rect 9817 -6193 9851 -6159
rect 9887 -6193 9934 -6159
rect 10186 -6193 10233 -6159
rect 10269 -6193 10303 -6159
rect 10339 -6193 10386 -6159
rect 10444 -6193 10491 -6159
rect 10527 -6193 10561 -6159
rect 10597 -6193 10644 -6159
rect 10702 -6193 10749 -6159
rect 10785 -6193 10819 -6159
rect 10855 -6193 10902 -6159
rect 10960 -6193 11007 -6159
rect 11043 -6193 11077 -6159
rect 11113 -6193 11160 -6159
rect 11412 -6193 11459 -6159
rect 11495 -6193 11529 -6159
rect 11565 -6193 11612 -6159
rect 11670 -6193 11717 -6159
rect 11753 -6193 11787 -6159
rect 11823 -6193 11870 -6159
rect 11928 -6193 11975 -6159
rect 12011 -6193 12045 -6159
rect 12081 -6193 12128 -6159
rect 12380 -6193 12427 -6159
rect 12463 -6193 12497 -6159
rect 12533 -6193 12580 -6159
rect 12638 -6193 12685 -6159
rect 12721 -6193 12755 -6159
rect 12791 -6193 12838 -6159
rect 12896 -6193 12943 -6159
rect 12979 -6193 13013 -6159
rect 13049 -6193 13096 -6159
rect 13154 -6193 13201 -6159
rect 13237 -6193 13271 -6159
rect 13307 -6193 13354 -6159
rect 13606 -6193 13653 -6159
rect 13689 -6193 13723 -6159
rect 13759 -6193 13806 -6159
rect 13931 -6190 13932 -6124
rect 18290 -5852 18324 -5830
rect 18290 -5920 18324 -5902
rect 18290 -5988 18324 -5974
rect 18290 -6056 18324 -6046
rect 18290 -6124 18324 -6118
rect 13931 -6192 13966 -6190
rect 9573 -6228 9607 -6226
rect 5214 -6300 5249 -6294
rect 5248 -6362 5249 -6300
rect 5214 -6372 5249 -6362
rect 5248 -6430 5249 -6372
rect 5214 -6444 5249 -6430
rect 5328 -6255 5362 -6236
rect 5328 -6323 5362 -6321
rect 5328 -6359 5362 -6357
rect 5328 -6444 5362 -6425
rect 5586 -6255 5620 -6236
rect 5586 -6323 5620 -6321
rect 5586 -6359 5620 -6357
rect 5586 -6444 5620 -6425
rect 5780 -6255 5814 -6236
rect 5780 -6323 5814 -6321
rect 5780 -6359 5814 -6357
rect 5780 -6444 5814 -6425
rect 6038 -6255 6072 -6236
rect 6038 -6323 6072 -6321
rect 6038 -6359 6072 -6357
rect 6038 -6444 6072 -6425
rect 6296 -6255 6330 -6236
rect 6296 -6323 6330 -6321
rect 6296 -6359 6330 -6357
rect 6296 -6444 6330 -6425
rect 6554 -6255 6588 -6236
rect 6554 -6323 6588 -6321
rect 6554 -6359 6588 -6357
rect 6554 -6444 6588 -6425
rect 6812 -6255 6846 -6236
rect 6812 -6323 6846 -6321
rect 6812 -6359 6846 -6357
rect 6812 -6444 6846 -6425
rect 7006 -6255 7040 -6236
rect 7006 -6323 7040 -6321
rect 7006 -6359 7040 -6357
rect 7006 -6444 7040 -6425
rect 7264 -6255 7298 -6236
rect 7264 -6323 7298 -6321
rect 7264 -6359 7298 -6357
rect 7264 -6444 7298 -6425
rect 7522 -6255 7556 -6236
rect 7522 -6323 7556 -6321
rect 7522 -6359 7556 -6357
rect 7522 -6444 7556 -6425
rect 7780 -6255 7814 -6236
rect 7780 -6323 7814 -6321
rect 7780 -6359 7814 -6357
rect 7780 -6444 7814 -6425
rect 7974 -6255 8008 -6236
rect 7974 -6323 8008 -6321
rect 7974 -6359 8008 -6357
rect 7974 -6444 8008 -6425
rect 8232 -6255 8266 -6236
rect 8232 -6323 8266 -6321
rect 8232 -6359 8266 -6357
rect 8232 -6444 8266 -6425
rect 8490 -6255 8524 -6236
rect 8490 -6323 8524 -6321
rect 8490 -6359 8524 -6357
rect 8490 -6444 8524 -6425
rect 8748 -6255 8782 -6236
rect 8748 -6323 8782 -6321
rect 8748 -6359 8782 -6357
rect 8748 -6444 8782 -6425
rect 9006 -6255 9040 -6236
rect 9006 -6323 9040 -6321
rect 9006 -6359 9040 -6357
rect 9006 -6444 9040 -6425
rect 9200 -6255 9234 -6236
rect 9200 -6323 9234 -6321
rect 9200 -6359 9234 -6357
rect 9200 -6444 9234 -6425
rect 9458 -6255 9492 -6236
rect 9458 -6323 9492 -6321
rect 9458 -6359 9492 -6357
rect 9458 -6444 9492 -6425
rect 13931 -6226 13932 -6192
rect 14092 -6193 14139 -6159
rect 14175 -6193 14209 -6159
rect 14245 -6193 14292 -6159
rect 14543 -6193 14590 -6159
rect 14626 -6193 14660 -6159
rect 14696 -6193 14743 -6159
rect 14801 -6193 14848 -6159
rect 14884 -6193 14918 -6159
rect 14954 -6193 15001 -6159
rect 15059 -6193 15106 -6159
rect 15142 -6193 15176 -6159
rect 15212 -6193 15259 -6159
rect 15317 -6193 15364 -6159
rect 15400 -6193 15434 -6159
rect 15470 -6193 15517 -6159
rect 15769 -6193 15816 -6159
rect 15852 -6193 15886 -6159
rect 15922 -6193 15969 -6159
rect 16027 -6193 16074 -6159
rect 16110 -6193 16144 -6159
rect 16180 -6193 16227 -6159
rect 16285 -6193 16332 -6159
rect 16368 -6193 16402 -6159
rect 16438 -6193 16485 -6159
rect 16737 -6193 16784 -6159
rect 16820 -6193 16854 -6159
rect 16890 -6193 16937 -6159
rect 16995 -6193 17042 -6159
rect 17078 -6193 17112 -6159
rect 17148 -6193 17195 -6159
rect 17253 -6193 17300 -6159
rect 17336 -6193 17370 -6159
rect 17406 -6193 17453 -6159
rect 17511 -6193 17558 -6159
rect 17594 -6193 17628 -6159
rect 17664 -6193 17711 -6159
rect 17963 -6193 18010 -6159
rect 18046 -6193 18080 -6159
rect 18116 -6193 18163 -6159
rect 18290 -6192 18324 -6190
rect 13931 -6228 13966 -6226
rect 9573 -6300 9607 -6294
rect 9573 -6372 9607 -6362
rect 9573 -6444 9607 -6430
rect 9688 -6255 9722 -6236
rect 9688 -6323 9722 -6321
rect 9688 -6359 9722 -6357
rect 9688 -6444 9722 -6425
rect 9946 -6255 9980 -6236
rect 9946 -6323 9980 -6321
rect 9946 -6359 9980 -6357
rect 9946 -6444 9980 -6425
rect 10140 -6255 10174 -6236
rect 10140 -6323 10174 -6321
rect 10140 -6359 10174 -6357
rect 10140 -6444 10174 -6425
rect 10398 -6255 10432 -6236
rect 10398 -6323 10432 -6321
rect 10398 -6359 10432 -6357
rect 10398 -6444 10432 -6425
rect 10656 -6255 10690 -6236
rect 10656 -6323 10690 -6321
rect 10656 -6359 10690 -6357
rect 10656 -6444 10690 -6425
rect 10914 -6255 10948 -6236
rect 10914 -6323 10948 -6321
rect 10914 -6359 10948 -6357
rect 10914 -6444 10948 -6425
rect 11172 -6255 11206 -6236
rect 11172 -6323 11206 -6321
rect 11172 -6359 11206 -6357
rect 11172 -6444 11206 -6425
rect 11366 -6255 11400 -6236
rect 11366 -6323 11400 -6321
rect 11366 -6359 11400 -6357
rect 11366 -6444 11400 -6425
rect 11624 -6255 11658 -6236
rect 11624 -6323 11658 -6321
rect 11624 -6359 11658 -6357
rect 11624 -6444 11658 -6425
rect 11882 -6255 11916 -6236
rect 11882 -6323 11916 -6321
rect 11882 -6359 11916 -6357
rect 11882 -6444 11916 -6425
rect 12140 -6255 12174 -6236
rect 12140 -6323 12174 -6321
rect 12140 -6359 12174 -6357
rect 12140 -6444 12174 -6425
rect 12334 -6255 12368 -6236
rect 12334 -6323 12368 -6321
rect 12334 -6359 12368 -6357
rect 12334 -6444 12368 -6425
rect 12592 -6255 12626 -6236
rect 12592 -6323 12626 -6321
rect 12592 -6359 12626 -6357
rect 12592 -6444 12626 -6425
rect 12850 -6255 12884 -6236
rect 12850 -6323 12884 -6321
rect 12850 -6359 12884 -6357
rect 12850 -6444 12884 -6425
rect 13108 -6255 13142 -6236
rect 13108 -6323 13142 -6321
rect 13108 -6359 13142 -6357
rect 13108 -6444 13142 -6425
rect 13366 -6255 13400 -6236
rect 13366 -6323 13400 -6321
rect 13366 -6359 13400 -6357
rect 13366 -6444 13400 -6425
rect 13560 -6255 13594 -6236
rect 13560 -6323 13594 -6321
rect 13560 -6359 13594 -6357
rect 13560 -6444 13594 -6425
rect 13818 -6255 13852 -6236
rect 13818 -6323 13852 -6321
rect 13818 -6359 13852 -6357
rect 13818 -6444 13852 -6425
rect 13931 -6294 13932 -6228
rect 18290 -6228 18324 -6226
rect 13931 -6300 13966 -6294
rect 13931 -6362 13932 -6300
rect 13931 -6372 13966 -6362
rect 13931 -6430 13932 -6372
rect 13931 -6444 13966 -6430
rect 14046 -6255 14080 -6236
rect 14046 -6323 14080 -6321
rect 14046 -6359 14080 -6357
rect 14046 -6444 14080 -6425
rect 14304 -6255 14338 -6236
rect 14304 -6323 14338 -6321
rect 14304 -6359 14338 -6357
rect 14304 -6444 14338 -6425
rect 14497 -6255 14531 -6236
rect 14497 -6323 14531 -6321
rect 14497 -6359 14531 -6357
rect 14497 -6444 14531 -6425
rect 14755 -6255 14789 -6236
rect 14755 -6323 14789 -6321
rect 14755 -6359 14789 -6357
rect 14755 -6444 14789 -6425
rect 15013 -6255 15047 -6236
rect 15013 -6323 15047 -6321
rect 15013 -6359 15047 -6357
rect 15013 -6444 15047 -6425
rect 15271 -6255 15305 -6236
rect 15271 -6323 15305 -6321
rect 15271 -6359 15305 -6357
rect 15271 -6444 15305 -6425
rect 15529 -6255 15563 -6236
rect 15529 -6323 15563 -6321
rect 15529 -6359 15563 -6357
rect 15529 -6444 15563 -6425
rect 15723 -6255 15757 -6236
rect 15723 -6323 15757 -6321
rect 15723 -6359 15757 -6357
rect 15723 -6444 15757 -6425
rect 15981 -6255 16015 -6236
rect 15981 -6323 16015 -6321
rect 15981 -6359 16015 -6357
rect 15981 -6444 16015 -6425
rect 16239 -6255 16273 -6236
rect 16239 -6323 16273 -6321
rect 16239 -6359 16273 -6357
rect 16239 -6444 16273 -6425
rect 16497 -6255 16531 -6236
rect 16497 -6323 16531 -6321
rect 16497 -6359 16531 -6357
rect 16497 -6444 16531 -6425
rect 16691 -6255 16725 -6236
rect 16691 -6323 16725 -6321
rect 16691 -6359 16725 -6357
rect 16691 -6444 16725 -6425
rect 16949 -6255 16983 -6236
rect 16949 -6323 16983 -6321
rect 16949 -6359 16983 -6357
rect 16949 -6444 16983 -6425
rect 17207 -6255 17241 -6236
rect 17207 -6323 17241 -6321
rect 17207 -6359 17241 -6357
rect 17207 -6444 17241 -6425
rect 17465 -6255 17499 -6236
rect 17465 -6323 17499 -6321
rect 17465 -6359 17499 -6357
rect 17465 -6444 17499 -6425
rect 17723 -6255 17757 -6236
rect 17723 -6323 17757 -6321
rect 17723 -6359 17757 -6357
rect 17723 -6444 17757 -6425
rect 17917 -6255 17951 -6236
rect 17917 -6323 17951 -6321
rect 17917 -6359 17951 -6357
rect 17917 -6444 17951 -6425
rect 18175 -6255 18209 -6236
rect 18175 -6323 18209 -6321
rect 18175 -6359 18209 -6357
rect 18175 -6444 18209 -6425
rect 18290 -6300 18324 -6294
rect 18290 -6372 18324 -6362
rect 18290 -6444 18324 -6430
rect 856 -6516 890 -6498
rect 856 -6588 890 -6566
rect 856 -6660 890 -6634
rect 856 -6732 890 -6702
rect 856 -6804 890 -6766
rect 5248 -6498 5249 -6444
rect 5214 -6516 5249 -6498
rect 5248 -6566 5249 -6516
rect 5214 -6588 5249 -6566
rect 5248 -6634 5249 -6588
rect 5214 -6660 5249 -6634
rect 5248 -6702 5249 -6660
rect 5214 -6732 5249 -6702
rect 5248 -6766 5249 -6732
rect 5214 -6804 5249 -6766
rect 9573 -6516 9607 -6498
rect 9573 -6588 9607 -6566
rect 9573 -6660 9607 -6634
rect 9573 -6732 9607 -6702
rect 9573 -6804 9607 -6766
rect 13931 -6498 13932 -6444
rect 13931 -6516 13966 -6498
rect 13931 -6566 13932 -6516
rect 13931 -6588 13966 -6566
rect 13931 -6634 13932 -6588
rect 13931 -6660 13966 -6634
rect 13931 -6702 13932 -6660
rect 13931 -6732 13966 -6702
rect 13931 -6766 13932 -6732
rect 13931 -6804 13966 -6766
rect 18290 -6516 18324 -6498
rect 18290 -6588 18324 -6566
rect 18290 -6660 18324 -6634
rect 18290 -6732 18324 -6702
rect 18290 -6804 18324 -6766
rect 890 -6838 977 -6804
rect 1011 -6838 1045 -6804
rect 1079 -6838 1113 -6804
rect 1147 -6838 1181 -6804
rect 1215 -6838 1249 -6804
rect 1283 -6838 1317 -6804
rect 1351 -6838 1385 -6804
rect 1419 -6838 1453 -6804
rect 1487 -6838 1521 -6804
rect 1555 -6838 1589 -6804
rect 1623 -6838 1657 -6804
rect 1691 -6838 1725 -6804
rect 1759 -6838 1793 -6804
rect 1827 -6838 1861 -6804
rect 1895 -6838 1929 -6804
rect 1963 -6838 1997 -6804
rect 2031 -6838 2065 -6804
rect 2099 -6838 2133 -6804
rect 2167 -6838 2201 -6804
rect 2235 -6838 2269 -6804
rect 2303 -6838 2337 -6804
rect 2371 -6838 2405 -6804
rect 2439 -6838 2473 -6804
rect 2507 -6838 2541 -6804
rect 2575 -6838 2609 -6804
rect 2643 -6838 2677 -6804
rect 2711 -6838 2745 -6804
rect 2779 -6838 2813 -6804
rect 2847 -6838 2881 -6804
rect 2915 -6838 2949 -6804
rect 2983 -6838 3017 -6804
rect 3051 -6838 3085 -6804
rect 3119 -6838 3153 -6804
rect 3187 -6838 3221 -6804
rect 3255 -6838 3289 -6804
rect 3323 -6838 3357 -6804
rect 3391 -6838 3425 -6804
rect 3459 -6838 3493 -6804
rect 3527 -6838 3561 -6804
rect 3595 -6838 3629 -6804
rect 3663 -6838 3697 -6804
rect 3731 -6838 3765 -6804
rect 3799 -6838 3833 -6804
rect 3867 -6838 3901 -6804
rect 3935 -6838 3969 -6804
rect 4003 -6838 4037 -6804
rect 4071 -6838 4105 -6804
rect 4139 -6838 4173 -6804
rect 4207 -6838 4241 -6804
rect 4275 -6838 4309 -6804
rect 4343 -6838 4377 -6804
rect 4411 -6838 4445 -6804
rect 4479 -6838 4513 -6804
rect 4547 -6838 4581 -6804
rect 4615 -6838 4649 -6804
rect 4683 -6838 4717 -6804
rect 4751 -6838 4785 -6804
rect 4819 -6838 4853 -6804
rect 4887 -6838 4921 -6804
rect 4955 -6838 4989 -6804
rect 5023 -6838 5057 -6804
rect 5091 -6838 5214 -6804
rect 5248 -6838 5372 -6804
rect 5406 -6838 5440 -6804
rect 5474 -6838 5508 -6804
rect 5542 -6838 5576 -6804
rect 5610 -6838 5644 -6804
rect 5678 -6838 5712 -6804
rect 5746 -6838 5780 -6804
rect 5814 -6838 5848 -6804
rect 5882 -6838 5916 -6804
rect 5950 -6838 5984 -6804
rect 6018 -6838 6052 -6804
rect 6086 -6838 6120 -6804
rect 6154 -6838 6188 -6804
rect 6222 -6838 6256 -6804
rect 6290 -6838 6324 -6804
rect 6358 -6838 6392 -6804
rect 6426 -6838 6460 -6804
rect 6494 -6838 6528 -6804
rect 6562 -6838 6596 -6804
rect 6630 -6838 6664 -6804
rect 6698 -6838 6732 -6804
rect 6766 -6838 6800 -6804
rect 6834 -6838 6868 -6804
rect 6902 -6838 6936 -6804
rect 6970 -6838 7004 -6804
rect 7038 -6838 7072 -6804
rect 7106 -6838 7140 -6804
rect 7174 -6838 7208 -6804
rect 7242 -6838 7276 -6804
rect 7310 -6838 7344 -6804
rect 7378 -6838 7412 -6804
rect 7446 -6838 7480 -6804
rect 7514 -6838 7548 -6804
rect 7582 -6838 7616 -6804
rect 7650 -6838 7684 -6804
rect 7718 -6838 7752 -6804
rect 7786 -6838 7820 -6804
rect 7854 -6838 7888 -6804
rect 7922 -6838 7956 -6804
rect 7990 -6838 8024 -6804
rect 8058 -6838 8092 -6804
rect 8126 -6838 8160 -6804
rect 8194 -6838 8228 -6804
rect 8262 -6838 8296 -6804
rect 8330 -6838 8364 -6804
rect 8398 -6838 8432 -6804
rect 8466 -6838 8500 -6804
rect 8534 -6838 8568 -6804
rect 8602 -6838 8636 -6804
rect 8670 -6838 8704 -6804
rect 8738 -6838 8772 -6804
rect 8806 -6838 8840 -6804
rect 8874 -6838 8908 -6804
rect 8942 -6838 8976 -6804
rect 9010 -6838 9044 -6804
rect 9078 -6838 9112 -6804
rect 9146 -6838 9180 -6804
rect 9214 -6838 9248 -6804
rect 9282 -6838 9316 -6804
rect 9350 -6838 9384 -6804
rect 9418 -6838 9452 -6804
rect 9486 -6838 9573 -6804
rect 9607 -6838 9694 -6804
rect 9728 -6838 9762 -6804
rect 9796 -6838 9830 -6804
rect 9864 -6838 9898 -6804
rect 9932 -6838 9966 -6804
rect 10000 -6838 10034 -6804
rect 10068 -6838 10102 -6804
rect 10136 -6838 10170 -6804
rect 10204 -6838 10238 -6804
rect 10272 -6838 10306 -6804
rect 10340 -6838 10374 -6804
rect 10408 -6838 10442 -6804
rect 10476 -6838 10510 -6804
rect 10544 -6838 10578 -6804
rect 10612 -6838 10646 -6804
rect 10680 -6838 10714 -6804
rect 10748 -6838 10782 -6804
rect 10816 -6838 10850 -6804
rect 10884 -6838 10918 -6804
rect 10952 -6838 10986 -6804
rect 11020 -6838 11054 -6804
rect 11088 -6838 11122 -6804
rect 11156 -6838 11190 -6804
rect 11224 -6838 11258 -6804
rect 11292 -6838 11326 -6804
rect 11360 -6838 11394 -6804
rect 11428 -6838 11462 -6804
rect 11496 -6838 11530 -6804
rect 11564 -6838 11598 -6804
rect 11632 -6838 11666 -6804
rect 11700 -6838 11734 -6804
rect 11768 -6838 11802 -6804
rect 11836 -6838 11870 -6804
rect 11904 -6838 11938 -6804
rect 11972 -6838 12006 -6804
rect 12040 -6838 12074 -6804
rect 12108 -6838 12142 -6804
rect 12176 -6838 12210 -6804
rect 12244 -6838 12278 -6804
rect 12312 -6838 12346 -6804
rect 12380 -6838 12414 -6804
rect 12448 -6838 12482 -6804
rect 12516 -6838 12550 -6804
rect 12584 -6838 12618 -6804
rect 12652 -6838 12686 -6804
rect 12720 -6838 12754 -6804
rect 12788 -6838 12822 -6804
rect 12856 -6838 12890 -6804
rect 12924 -6838 12958 -6804
rect 12992 -6838 13026 -6804
rect 13060 -6838 13094 -6804
rect 13128 -6838 13162 -6804
rect 13196 -6838 13230 -6804
rect 13264 -6838 13298 -6804
rect 13332 -6838 13366 -6804
rect 13400 -6838 13434 -6804
rect 13468 -6838 13502 -6804
rect 13536 -6838 13570 -6804
rect 13604 -6838 13638 -6804
rect 13672 -6838 13706 -6804
rect 13740 -6838 13774 -6804
rect 13808 -6838 13932 -6804
rect 13966 -6838 14089 -6804
rect 14123 -6838 14157 -6804
rect 14191 -6838 14225 -6804
rect 14259 -6838 14293 -6804
rect 14327 -6838 14361 -6804
rect 14395 -6838 14429 -6804
rect 14463 -6838 14497 -6804
rect 14531 -6838 14565 -6804
rect 14599 -6838 14633 -6804
rect 14667 -6838 14701 -6804
rect 14735 -6838 14769 -6804
rect 14803 -6838 14837 -6804
rect 14871 -6838 14905 -6804
rect 14939 -6838 14973 -6804
rect 15007 -6838 15041 -6804
rect 15075 -6838 15109 -6804
rect 15143 -6838 15177 -6804
rect 15211 -6838 15245 -6804
rect 15279 -6838 15313 -6804
rect 15347 -6838 15381 -6804
rect 15415 -6838 15449 -6804
rect 15483 -6838 15517 -6804
rect 15551 -6838 15585 -6804
rect 15619 -6838 15653 -6804
rect 15687 -6838 15721 -6804
rect 15755 -6838 15789 -6804
rect 15823 -6838 15857 -6804
rect 15891 -6838 15925 -6804
rect 15959 -6838 15993 -6804
rect 16027 -6838 16061 -6804
rect 16095 -6838 16129 -6804
rect 16163 -6838 16197 -6804
rect 16231 -6838 16265 -6804
rect 16299 -6838 16333 -6804
rect 16367 -6838 16401 -6804
rect 16435 -6838 16469 -6804
rect 16503 -6838 16537 -6804
rect 16571 -6838 16605 -6804
rect 16639 -6838 16673 -6804
rect 16707 -6838 16741 -6804
rect 16775 -6838 16809 -6804
rect 16843 -6838 16877 -6804
rect 16911 -6838 16945 -6804
rect 16979 -6838 17013 -6804
rect 17047 -6838 17081 -6804
rect 17115 -6838 17149 -6804
rect 17183 -6838 17217 -6804
rect 17251 -6838 17285 -6804
rect 17319 -6838 17353 -6804
rect 17387 -6838 17421 -6804
rect 17455 -6838 17489 -6804
rect 17523 -6838 17557 -6804
rect 17591 -6838 17625 -6804
rect 17659 -6838 17693 -6804
rect 17727 -6838 17761 -6804
rect 17795 -6838 17829 -6804
rect 17863 -6838 17897 -6804
rect 17931 -6838 17965 -6804
rect 17999 -6838 18033 -6804
rect 18067 -6838 18101 -6804
rect 18135 -6838 18169 -6804
rect 18203 -6838 18290 -6804
rect 856 -6876 890 -6838
rect 856 -6940 890 -6910
rect 856 -7008 890 -6982
rect 856 -7076 890 -7054
rect 856 -7144 890 -7126
rect 5214 -6876 5249 -6838
rect 5248 -6910 5249 -6876
rect 5214 -6940 5249 -6910
rect 5248 -6982 5249 -6940
rect 5214 -7008 5249 -6982
rect 5248 -7054 5249 -7008
rect 5214 -7076 5249 -7054
rect 5248 -7126 5249 -7076
rect 5214 -7144 5249 -7126
rect 856 -7212 890 -7198
rect 856 -7280 890 -7270
rect 856 -7348 890 -7342
rect 971 -7212 1005 -7193
rect 971 -7280 1005 -7278
rect 971 -7316 1005 -7314
rect 971 -7401 1005 -7382
rect 1229 -7212 1263 -7193
rect 1229 -7280 1263 -7278
rect 1229 -7316 1263 -7314
rect 1229 -7401 1263 -7382
rect 1423 -7212 1457 -7193
rect 1423 -7280 1457 -7278
rect 1423 -7316 1457 -7314
rect 1423 -7401 1457 -7382
rect 1681 -7212 1715 -7193
rect 1681 -7280 1715 -7278
rect 1681 -7316 1715 -7314
rect 1681 -7401 1715 -7382
rect 1939 -7212 1973 -7193
rect 1939 -7280 1973 -7278
rect 1939 -7316 1973 -7314
rect 1939 -7401 1973 -7382
rect 2197 -7212 2231 -7193
rect 2197 -7280 2231 -7278
rect 2197 -7316 2231 -7314
rect 2197 -7401 2231 -7382
rect 2455 -7212 2489 -7193
rect 2455 -7280 2489 -7278
rect 2455 -7316 2489 -7314
rect 2455 -7401 2489 -7382
rect 2649 -7212 2683 -7193
rect 2649 -7280 2683 -7278
rect 2649 -7316 2683 -7314
rect 2649 -7401 2683 -7382
rect 2907 -7212 2941 -7193
rect 2907 -7280 2941 -7278
rect 2907 -7316 2941 -7314
rect 2907 -7401 2941 -7382
rect 3165 -7212 3199 -7193
rect 3165 -7280 3199 -7278
rect 3165 -7316 3199 -7314
rect 3165 -7401 3199 -7382
rect 3423 -7212 3457 -7193
rect 3423 -7280 3457 -7278
rect 3423 -7316 3457 -7314
rect 3423 -7401 3457 -7382
rect 3617 -7212 3651 -7193
rect 3617 -7280 3651 -7278
rect 3617 -7316 3651 -7314
rect 3617 -7401 3651 -7382
rect 3875 -7212 3909 -7193
rect 3875 -7280 3909 -7278
rect 3875 -7316 3909 -7314
rect 3875 -7401 3909 -7382
rect 4133 -7212 4167 -7193
rect 4133 -7280 4167 -7278
rect 4133 -7316 4167 -7314
rect 4133 -7401 4167 -7382
rect 4391 -7212 4425 -7193
rect 4391 -7280 4425 -7278
rect 4391 -7316 4425 -7314
rect 4391 -7401 4425 -7382
rect 4649 -7212 4683 -7193
rect 4649 -7280 4683 -7278
rect 4649 -7316 4683 -7314
rect 4649 -7401 4683 -7382
rect 4842 -7212 4876 -7193
rect 4842 -7280 4876 -7278
rect 4842 -7316 4876 -7314
rect 4842 -7401 4876 -7382
rect 5100 -7212 5134 -7193
rect 5100 -7280 5134 -7278
rect 5100 -7316 5134 -7314
rect 5100 -7401 5134 -7382
rect 5248 -7198 5249 -7144
rect 9573 -6876 9607 -6838
rect 9573 -6940 9607 -6910
rect 9573 -7008 9607 -6982
rect 9573 -7076 9607 -7054
rect 9573 -7144 9607 -7126
rect 5214 -7212 5249 -7198
rect 5248 -7270 5249 -7212
rect 5214 -7280 5249 -7270
rect 5248 -7342 5249 -7280
rect 5214 -7348 5249 -7342
rect 856 -7416 890 -7414
rect 5248 -7414 5249 -7348
rect 5328 -7212 5362 -7193
rect 5328 -7280 5362 -7278
rect 5328 -7316 5362 -7314
rect 5328 -7401 5362 -7382
rect 5586 -7212 5620 -7193
rect 5586 -7280 5620 -7278
rect 5586 -7316 5620 -7314
rect 5586 -7401 5620 -7382
rect 5780 -7212 5814 -7193
rect 5780 -7280 5814 -7278
rect 5780 -7316 5814 -7314
rect 5780 -7401 5814 -7382
rect 6038 -7212 6072 -7193
rect 6038 -7280 6072 -7278
rect 6038 -7316 6072 -7314
rect 6038 -7401 6072 -7382
rect 6296 -7212 6330 -7193
rect 6296 -7280 6330 -7278
rect 6296 -7316 6330 -7314
rect 6296 -7401 6330 -7382
rect 6554 -7212 6588 -7193
rect 6554 -7280 6588 -7278
rect 6554 -7316 6588 -7314
rect 6554 -7401 6588 -7382
rect 6812 -7212 6846 -7193
rect 6812 -7280 6846 -7278
rect 6812 -7316 6846 -7314
rect 6812 -7401 6846 -7382
rect 7006 -7212 7040 -7193
rect 7006 -7280 7040 -7278
rect 7006 -7316 7040 -7314
rect 7006 -7401 7040 -7382
rect 7264 -7212 7298 -7193
rect 7264 -7280 7298 -7278
rect 7264 -7316 7298 -7314
rect 7264 -7401 7298 -7382
rect 7522 -7212 7556 -7193
rect 7522 -7280 7556 -7278
rect 7522 -7316 7556 -7314
rect 7522 -7401 7556 -7382
rect 7780 -7212 7814 -7193
rect 7780 -7280 7814 -7278
rect 7780 -7316 7814 -7314
rect 7780 -7401 7814 -7382
rect 7974 -7212 8008 -7193
rect 7974 -7280 8008 -7278
rect 7974 -7316 8008 -7314
rect 7974 -7401 8008 -7382
rect 8232 -7212 8266 -7193
rect 8232 -7280 8266 -7278
rect 8232 -7316 8266 -7314
rect 8232 -7401 8266 -7382
rect 8490 -7212 8524 -7193
rect 8490 -7280 8524 -7278
rect 8490 -7316 8524 -7314
rect 8490 -7401 8524 -7382
rect 8748 -7212 8782 -7193
rect 8748 -7280 8782 -7278
rect 8748 -7316 8782 -7314
rect 8748 -7401 8782 -7382
rect 9006 -7212 9040 -7193
rect 9006 -7280 9040 -7278
rect 9006 -7316 9040 -7314
rect 9006 -7401 9040 -7382
rect 9200 -7212 9234 -7193
rect 9200 -7280 9234 -7278
rect 9200 -7316 9234 -7314
rect 9200 -7401 9234 -7382
rect 9458 -7212 9492 -7193
rect 9458 -7280 9492 -7278
rect 9458 -7316 9492 -7314
rect 9458 -7401 9492 -7382
rect 13931 -6876 13966 -6838
rect 13931 -6910 13932 -6876
rect 13931 -6940 13966 -6910
rect 13931 -6982 13932 -6940
rect 13931 -7008 13966 -6982
rect 13931 -7054 13932 -7008
rect 13931 -7076 13966 -7054
rect 13931 -7126 13932 -7076
rect 13931 -7144 13966 -7126
rect 9573 -7212 9607 -7198
rect 9573 -7280 9607 -7270
rect 9573 -7348 9607 -7342
rect 5214 -7416 5249 -7414
rect 856 -7452 890 -7450
rect 1017 -7478 1064 -7444
rect 1100 -7478 1134 -7444
rect 1170 -7478 1217 -7444
rect 1469 -7478 1516 -7444
rect 1552 -7478 1586 -7444
rect 1622 -7478 1669 -7444
rect 1727 -7478 1774 -7444
rect 1810 -7478 1844 -7444
rect 1880 -7478 1927 -7444
rect 1985 -7478 2032 -7444
rect 2068 -7478 2102 -7444
rect 2138 -7478 2185 -7444
rect 2243 -7478 2290 -7444
rect 2326 -7478 2360 -7444
rect 2396 -7478 2443 -7444
rect 2695 -7478 2742 -7444
rect 2778 -7478 2812 -7444
rect 2848 -7478 2895 -7444
rect 2953 -7478 3000 -7444
rect 3036 -7478 3070 -7444
rect 3106 -7478 3153 -7444
rect 3211 -7478 3258 -7444
rect 3294 -7478 3328 -7444
rect 3364 -7478 3411 -7444
rect 3663 -7478 3710 -7444
rect 3746 -7478 3780 -7444
rect 3816 -7478 3863 -7444
rect 3921 -7478 3968 -7444
rect 4004 -7478 4038 -7444
rect 4074 -7478 4121 -7444
rect 4179 -7478 4226 -7444
rect 4262 -7478 4296 -7444
rect 4332 -7478 4379 -7444
rect 4437 -7478 4484 -7444
rect 4520 -7478 4554 -7444
rect 4590 -7478 4637 -7444
rect 4888 -7478 4935 -7444
rect 4971 -7478 5005 -7444
rect 5041 -7478 5088 -7444
rect 5248 -7450 5249 -7416
rect 9688 -7212 9722 -7193
rect 9688 -7280 9722 -7278
rect 9688 -7316 9722 -7314
rect 9688 -7401 9722 -7382
rect 9946 -7212 9980 -7193
rect 9946 -7280 9980 -7278
rect 9946 -7316 9980 -7314
rect 9946 -7401 9980 -7382
rect 10140 -7212 10174 -7193
rect 10140 -7280 10174 -7278
rect 10140 -7316 10174 -7314
rect 10140 -7401 10174 -7382
rect 10398 -7212 10432 -7193
rect 10398 -7280 10432 -7278
rect 10398 -7316 10432 -7314
rect 10398 -7401 10432 -7382
rect 10656 -7212 10690 -7193
rect 10656 -7280 10690 -7278
rect 10656 -7316 10690 -7314
rect 10656 -7401 10690 -7382
rect 10914 -7212 10948 -7193
rect 10914 -7280 10948 -7278
rect 10914 -7316 10948 -7314
rect 10914 -7401 10948 -7382
rect 11172 -7212 11206 -7193
rect 11172 -7280 11206 -7278
rect 11172 -7316 11206 -7314
rect 11172 -7401 11206 -7382
rect 11366 -7212 11400 -7193
rect 11366 -7280 11400 -7278
rect 11366 -7316 11400 -7314
rect 11366 -7401 11400 -7382
rect 11624 -7212 11658 -7193
rect 11624 -7280 11658 -7278
rect 11624 -7316 11658 -7314
rect 11624 -7401 11658 -7382
rect 11882 -7212 11916 -7193
rect 11882 -7280 11916 -7278
rect 11882 -7316 11916 -7314
rect 11882 -7401 11916 -7382
rect 12140 -7212 12174 -7193
rect 12140 -7280 12174 -7278
rect 12140 -7316 12174 -7314
rect 12140 -7401 12174 -7382
rect 12334 -7212 12368 -7193
rect 12334 -7280 12368 -7278
rect 12334 -7316 12368 -7314
rect 12334 -7401 12368 -7382
rect 12592 -7212 12626 -7193
rect 12592 -7280 12626 -7278
rect 12592 -7316 12626 -7314
rect 12592 -7401 12626 -7382
rect 12850 -7212 12884 -7193
rect 12850 -7280 12884 -7278
rect 12850 -7316 12884 -7314
rect 12850 -7401 12884 -7382
rect 13108 -7212 13142 -7193
rect 13108 -7280 13142 -7278
rect 13108 -7316 13142 -7314
rect 13108 -7401 13142 -7382
rect 13366 -7212 13400 -7193
rect 13366 -7280 13400 -7278
rect 13366 -7316 13400 -7314
rect 13366 -7401 13400 -7382
rect 13560 -7212 13594 -7193
rect 13560 -7280 13594 -7278
rect 13560 -7316 13594 -7314
rect 13560 -7401 13594 -7382
rect 13818 -7212 13852 -7193
rect 13818 -7280 13852 -7278
rect 13818 -7316 13852 -7314
rect 13818 -7401 13852 -7382
rect 13931 -7198 13932 -7144
rect 18290 -6876 18324 -6838
rect 18290 -6940 18324 -6910
rect 18290 -7008 18324 -6982
rect 18290 -7076 18324 -7054
rect 18290 -7144 18324 -7126
rect 13931 -7212 13966 -7198
rect 13931 -7270 13932 -7212
rect 13931 -7280 13966 -7270
rect 13931 -7342 13932 -7280
rect 13931 -7348 13966 -7342
rect 9573 -7416 9607 -7414
rect 5214 -7452 5249 -7450
rect 856 -7524 890 -7518
rect 856 -7596 890 -7586
rect 856 -7668 890 -7654
rect 856 -7740 890 -7722
rect 856 -7812 890 -7790
rect 5248 -7518 5249 -7452
rect 5374 -7478 5421 -7444
rect 5457 -7478 5491 -7444
rect 5527 -7478 5574 -7444
rect 5826 -7478 5873 -7444
rect 5909 -7478 5943 -7444
rect 5979 -7478 6026 -7444
rect 6084 -7478 6131 -7444
rect 6167 -7478 6201 -7444
rect 6237 -7478 6284 -7444
rect 6342 -7478 6389 -7444
rect 6425 -7478 6459 -7444
rect 6495 -7478 6542 -7444
rect 6600 -7478 6647 -7444
rect 6683 -7478 6717 -7444
rect 6753 -7478 6800 -7444
rect 7052 -7478 7099 -7444
rect 7135 -7478 7169 -7444
rect 7205 -7478 7252 -7444
rect 7310 -7478 7357 -7444
rect 7393 -7478 7427 -7444
rect 7463 -7478 7510 -7444
rect 7568 -7478 7615 -7444
rect 7651 -7478 7685 -7444
rect 7721 -7478 7768 -7444
rect 8020 -7478 8067 -7444
rect 8103 -7478 8137 -7444
rect 8173 -7478 8220 -7444
rect 8278 -7478 8325 -7444
rect 8361 -7478 8395 -7444
rect 8431 -7478 8478 -7444
rect 8536 -7478 8583 -7444
rect 8619 -7478 8653 -7444
rect 8689 -7478 8736 -7444
rect 8794 -7478 8841 -7444
rect 8877 -7478 8911 -7444
rect 8947 -7478 8994 -7444
rect 9246 -7478 9293 -7444
rect 9329 -7478 9363 -7444
rect 9399 -7478 9446 -7444
rect 13931 -7414 13932 -7348
rect 14046 -7212 14080 -7193
rect 14046 -7280 14080 -7278
rect 14046 -7316 14080 -7314
rect 14046 -7401 14080 -7382
rect 14304 -7212 14338 -7193
rect 14304 -7280 14338 -7278
rect 14304 -7316 14338 -7314
rect 14304 -7401 14338 -7382
rect 14497 -7212 14531 -7193
rect 14497 -7280 14531 -7278
rect 14497 -7316 14531 -7314
rect 14497 -7401 14531 -7382
rect 14755 -7212 14789 -7193
rect 14755 -7280 14789 -7278
rect 14755 -7316 14789 -7314
rect 14755 -7401 14789 -7382
rect 15013 -7212 15047 -7193
rect 15013 -7280 15047 -7278
rect 15013 -7316 15047 -7314
rect 15013 -7401 15047 -7382
rect 15271 -7212 15305 -7193
rect 15271 -7280 15305 -7278
rect 15271 -7316 15305 -7314
rect 15271 -7401 15305 -7382
rect 15529 -7212 15563 -7193
rect 15529 -7280 15563 -7278
rect 15529 -7316 15563 -7314
rect 15529 -7401 15563 -7382
rect 15723 -7212 15757 -7193
rect 15723 -7280 15757 -7278
rect 15723 -7316 15757 -7314
rect 15723 -7401 15757 -7382
rect 15981 -7212 16015 -7193
rect 15981 -7280 16015 -7278
rect 15981 -7316 16015 -7314
rect 15981 -7401 16015 -7382
rect 16239 -7212 16273 -7193
rect 16239 -7280 16273 -7278
rect 16239 -7316 16273 -7314
rect 16239 -7401 16273 -7382
rect 16497 -7212 16531 -7193
rect 16497 -7280 16531 -7278
rect 16497 -7316 16531 -7314
rect 16497 -7401 16531 -7382
rect 16691 -7212 16725 -7193
rect 16691 -7280 16725 -7278
rect 16691 -7316 16725 -7314
rect 16691 -7401 16725 -7382
rect 16949 -7212 16983 -7193
rect 16949 -7280 16983 -7278
rect 16949 -7316 16983 -7314
rect 16949 -7401 16983 -7382
rect 17207 -7212 17241 -7193
rect 17207 -7280 17241 -7278
rect 17207 -7316 17241 -7314
rect 17207 -7401 17241 -7382
rect 17465 -7212 17499 -7193
rect 17465 -7280 17499 -7278
rect 17465 -7316 17499 -7314
rect 17465 -7401 17499 -7382
rect 17723 -7212 17757 -7193
rect 17723 -7280 17757 -7278
rect 17723 -7316 17757 -7314
rect 17723 -7401 17757 -7382
rect 17917 -7212 17951 -7193
rect 17917 -7280 17951 -7278
rect 17917 -7316 17951 -7314
rect 17917 -7401 17951 -7382
rect 18175 -7212 18209 -7193
rect 18175 -7280 18209 -7278
rect 18175 -7316 18209 -7314
rect 18175 -7401 18209 -7382
rect 18290 -7212 18324 -7198
rect 18290 -7280 18324 -7270
rect 18290 -7348 18324 -7342
rect 13931 -7416 13966 -7414
rect 9573 -7452 9607 -7450
rect 5214 -7524 5249 -7518
rect 5248 -7586 5249 -7524
rect 5214 -7596 5249 -7586
rect 5248 -7654 5249 -7596
rect 5214 -7668 5249 -7654
rect 5248 -7722 5249 -7668
rect 5214 -7740 5249 -7722
rect 5248 -7790 5249 -7740
rect 1017 -7840 1064 -7806
rect 1100 -7840 1134 -7806
rect 1170 -7840 1217 -7806
rect 1469 -7840 1516 -7806
rect 1552 -7840 1586 -7806
rect 1622 -7840 1669 -7806
rect 1727 -7840 1774 -7806
rect 1810 -7840 1844 -7806
rect 1880 -7840 1927 -7806
rect 1985 -7840 2032 -7806
rect 2068 -7840 2102 -7806
rect 2138 -7840 2185 -7806
rect 2243 -7840 2290 -7806
rect 2326 -7840 2360 -7806
rect 2396 -7840 2443 -7806
rect 2695 -7840 2742 -7806
rect 2778 -7840 2812 -7806
rect 2848 -7840 2895 -7806
rect 2953 -7840 3000 -7806
rect 3036 -7840 3070 -7806
rect 3106 -7840 3153 -7806
rect 3211 -7840 3258 -7806
rect 3294 -7840 3328 -7806
rect 3364 -7840 3411 -7806
rect 3663 -7840 3710 -7806
rect 3746 -7840 3780 -7806
rect 3816 -7840 3863 -7806
rect 3921 -7840 3968 -7806
rect 4004 -7840 4038 -7806
rect 4074 -7840 4121 -7806
rect 4179 -7840 4226 -7806
rect 4262 -7840 4296 -7806
rect 4332 -7840 4379 -7806
rect 4437 -7840 4484 -7806
rect 4520 -7840 4554 -7806
rect 4590 -7840 4637 -7806
rect 4888 -7840 4935 -7806
rect 4971 -7840 5005 -7806
rect 5041 -7840 5088 -7806
rect 5214 -7812 5249 -7790
rect 9734 -7478 9781 -7444
rect 9817 -7478 9851 -7444
rect 9887 -7478 9934 -7444
rect 10186 -7478 10233 -7444
rect 10269 -7478 10303 -7444
rect 10339 -7478 10386 -7444
rect 10444 -7478 10491 -7444
rect 10527 -7478 10561 -7444
rect 10597 -7478 10644 -7444
rect 10702 -7478 10749 -7444
rect 10785 -7478 10819 -7444
rect 10855 -7478 10902 -7444
rect 10960 -7478 11007 -7444
rect 11043 -7478 11077 -7444
rect 11113 -7478 11160 -7444
rect 11412 -7478 11459 -7444
rect 11495 -7478 11529 -7444
rect 11565 -7478 11612 -7444
rect 11670 -7478 11717 -7444
rect 11753 -7478 11787 -7444
rect 11823 -7478 11870 -7444
rect 11928 -7478 11975 -7444
rect 12011 -7478 12045 -7444
rect 12081 -7478 12128 -7444
rect 12380 -7478 12427 -7444
rect 12463 -7478 12497 -7444
rect 12533 -7478 12580 -7444
rect 12638 -7478 12685 -7444
rect 12721 -7478 12755 -7444
rect 12791 -7478 12838 -7444
rect 12896 -7478 12943 -7444
rect 12979 -7478 13013 -7444
rect 13049 -7478 13096 -7444
rect 13154 -7478 13201 -7444
rect 13237 -7478 13271 -7444
rect 13307 -7478 13354 -7444
rect 13606 -7478 13653 -7444
rect 13689 -7478 13723 -7444
rect 13759 -7478 13806 -7444
rect 13931 -7450 13932 -7416
rect 18290 -7416 18324 -7414
rect 13931 -7452 13966 -7450
rect 9573 -7524 9607 -7518
rect 9573 -7596 9607 -7586
rect 9573 -7668 9607 -7654
rect 9573 -7740 9607 -7722
rect 856 -7884 890 -7858
rect 5248 -7858 5249 -7812
rect 5374 -7840 5421 -7806
rect 5457 -7840 5491 -7806
rect 5527 -7840 5574 -7806
rect 5826 -7840 5873 -7806
rect 5909 -7840 5943 -7806
rect 5979 -7840 6026 -7806
rect 6084 -7840 6131 -7806
rect 6167 -7840 6201 -7806
rect 6237 -7840 6284 -7806
rect 6342 -7840 6389 -7806
rect 6425 -7840 6459 -7806
rect 6495 -7840 6542 -7806
rect 6600 -7840 6647 -7806
rect 6683 -7840 6717 -7806
rect 6753 -7840 6800 -7806
rect 7052 -7840 7099 -7806
rect 7135 -7840 7169 -7806
rect 7205 -7840 7252 -7806
rect 7310 -7840 7357 -7806
rect 7393 -7840 7427 -7806
rect 7463 -7840 7510 -7806
rect 7568 -7840 7615 -7806
rect 7651 -7840 7685 -7806
rect 7721 -7840 7768 -7806
rect 8020 -7840 8067 -7806
rect 8103 -7840 8137 -7806
rect 8173 -7840 8220 -7806
rect 8278 -7840 8325 -7806
rect 8361 -7840 8395 -7806
rect 8431 -7840 8478 -7806
rect 8536 -7840 8583 -7806
rect 8619 -7840 8653 -7806
rect 8689 -7840 8736 -7806
rect 8794 -7840 8841 -7806
rect 8877 -7840 8911 -7806
rect 8947 -7840 8994 -7806
rect 9246 -7840 9293 -7806
rect 9329 -7840 9363 -7806
rect 9399 -7840 9446 -7806
rect 9573 -7812 9607 -7790
rect 13931 -7518 13932 -7452
rect 14092 -7478 14139 -7444
rect 14175 -7478 14209 -7444
rect 14245 -7478 14292 -7444
rect 14543 -7478 14590 -7444
rect 14626 -7478 14660 -7444
rect 14696 -7478 14743 -7444
rect 14801 -7478 14848 -7444
rect 14884 -7478 14918 -7444
rect 14954 -7478 15001 -7444
rect 15059 -7478 15106 -7444
rect 15142 -7478 15176 -7444
rect 15212 -7478 15259 -7444
rect 15317 -7478 15364 -7444
rect 15400 -7478 15434 -7444
rect 15470 -7478 15517 -7444
rect 15769 -7478 15816 -7444
rect 15852 -7478 15886 -7444
rect 15922 -7478 15969 -7444
rect 16027 -7478 16074 -7444
rect 16110 -7478 16144 -7444
rect 16180 -7478 16227 -7444
rect 16285 -7478 16332 -7444
rect 16368 -7478 16402 -7444
rect 16438 -7478 16485 -7444
rect 16737 -7478 16784 -7444
rect 16820 -7478 16854 -7444
rect 16890 -7478 16937 -7444
rect 16995 -7478 17042 -7444
rect 17078 -7478 17112 -7444
rect 17148 -7478 17195 -7444
rect 17253 -7478 17300 -7444
rect 17336 -7478 17370 -7444
rect 17406 -7478 17453 -7444
rect 17511 -7478 17558 -7444
rect 17594 -7478 17628 -7444
rect 17664 -7478 17711 -7444
rect 17963 -7478 18010 -7444
rect 18046 -7478 18080 -7444
rect 18116 -7478 18163 -7444
rect 18290 -7452 18324 -7450
rect 13931 -7524 13966 -7518
rect 13931 -7586 13932 -7524
rect 13931 -7596 13966 -7586
rect 13931 -7654 13932 -7596
rect 13931 -7668 13966 -7654
rect 13931 -7722 13932 -7668
rect 13931 -7740 13966 -7722
rect 13931 -7790 13932 -7740
rect 856 -7956 890 -7926
rect 856 -8028 890 -7994
rect 856 -8096 890 -8062
rect 971 -7902 1005 -7883
rect 971 -7970 1005 -7968
rect 971 -8006 1005 -8004
rect 971 -8091 1005 -8072
rect 1229 -7902 1263 -7883
rect 1229 -7970 1263 -7968
rect 1229 -8006 1263 -8004
rect 1229 -8091 1263 -8072
rect 1423 -7902 1457 -7883
rect 1423 -7970 1457 -7968
rect 1423 -8006 1457 -8004
rect 1423 -8091 1457 -8072
rect 1681 -7902 1715 -7883
rect 1681 -7970 1715 -7968
rect 1681 -8006 1715 -8004
rect 1681 -8091 1715 -8072
rect 1939 -7902 1973 -7883
rect 1939 -7970 1973 -7968
rect 1939 -8006 1973 -8004
rect 1939 -8091 1973 -8072
rect 2197 -7902 2231 -7883
rect 2197 -7970 2231 -7968
rect 2197 -8006 2231 -8004
rect 2197 -8091 2231 -8072
rect 2455 -7902 2489 -7883
rect 2455 -7970 2489 -7968
rect 2455 -8006 2489 -8004
rect 2455 -8091 2489 -8072
rect 2649 -7902 2683 -7883
rect 2649 -7970 2683 -7968
rect 2649 -8006 2683 -8004
rect 2649 -8091 2683 -8072
rect 2907 -7902 2941 -7883
rect 2907 -7970 2941 -7968
rect 2907 -8006 2941 -8004
rect 2907 -8091 2941 -8072
rect 3165 -7902 3199 -7883
rect 3165 -7970 3199 -7968
rect 3165 -8006 3199 -8004
rect 3165 -8091 3199 -8072
rect 3423 -7902 3457 -7883
rect 3423 -7970 3457 -7968
rect 3423 -8006 3457 -8004
rect 3423 -8091 3457 -8072
rect 3617 -7902 3651 -7883
rect 3617 -7970 3651 -7968
rect 3617 -8006 3651 -8004
rect 3617 -8091 3651 -8072
rect 3875 -7902 3909 -7883
rect 3875 -7970 3909 -7968
rect 3875 -8006 3909 -8004
rect 3875 -8091 3909 -8072
rect 4133 -7902 4167 -7883
rect 4133 -7970 4167 -7968
rect 4133 -8006 4167 -8004
rect 4133 -8091 4167 -8072
rect 4391 -7902 4425 -7883
rect 4391 -7970 4425 -7968
rect 4391 -8006 4425 -8004
rect 4391 -8091 4425 -8072
rect 4649 -7902 4683 -7883
rect 4649 -7970 4683 -7968
rect 4649 -8006 4683 -8004
rect 4649 -8091 4683 -8072
rect 4842 -7902 4876 -7883
rect 4842 -7970 4876 -7968
rect 4842 -8006 4876 -8004
rect 4842 -8091 4876 -8072
rect 5100 -7902 5134 -7883
rect 5100 -7970 5134 -7968
rect 5100 -8006 5134 -8004
rect 5100 -8091 5134 -8072
rect 5214 -7884 5249 -7858
rect 9734 -7840 9781 -7806
rect 9817 -7840 9851 -7806
rect 9887 -7840 9934 -7806
rect 10186 -7840 10233 -7806
rect 10269 -7840 10303 -7806
rect 10339 -7840 10386 -7806
rect 10444 -7840 10491 -7806
rect 10527 -7840 10561 -7806
rect 10597 -7840 10644 -7806
rect 10702 -7840 10749 -7806
rect 10785 -7840 10819 -7806
rect 10855 -7840 10902 -7806
rect 10960 -7840 11007 -7806
rect 11043 -7840 11077 -7806
rect 11113 -7840 11160 -7806
rect 11412 -7840 11459 -7806
rect 11495 -7840 11529 -7806
rect 11565 -7840 11612 -7806
rect 11670 -7840 11717 -7806
rect 11753 -7840 11787 -7806
rect 11823 -7840 11870 -7806
rect 11928 -7840 11975 -7806
rect 12011 -7840 12045 -7806
rect 12081 -7840 12128 -7806
rect 12380 -7840 12427 -7806
rect 12463 -7840 12497 -7806
rect 12533 -7840 12580 -7806
rect 12638 -7840 12685 -7806
rect 12721 -7840 12755 -7806
rect 12791 -7840 12838 -7806
rect 12896 -7840 12943 -7806
rect 12979 -7840 13013 -7806
rect 13049 -7840 13096 -7806
rect 13154 -7840 13201 -7806
rect 13237 -7840 13271 -7806
rect 13307 -7840 13354 -7806
rect 13606 -7840 13653 -7806
rect 13689 -7840 13723 -7806
rect 13759 -7840 13806 -7806
rect 13931 -7812 13966 -7790
rect 18290 -7524 18324 -7518
rect 18290 -7596 18324 -7586
rect 18290 -7668 18324 -7654
rect 18290 -7740 18324 -7722
rect 5248 -7926 5249 -7884
rect 5214 -7956 5249 -7926
rect 5248 -7994 5249 -7956
rect 5214 -8028 5249 -7994
rect 5248 -8062 5249 -8028
rect 856 -8164 890 -8134
rect 856 -8232 890 -8206
rect 856 -8300 890 -8278
rect 856 -8368 890 -8350
rect 5214 -8096 5249 -8062
rect 5328 -7902 5362 -7883
rect 5328 -7970 5362 -7968
rect 5328 -8006 5362 -8004
rect 5328 -8091 5362 -8072
rect 5586 -7902 5620 -7883
rect 5586 -7970 5620 -7968
rect 5586 -8006 5620 -8004
rect 5586 -8091 5620 -8072
rect 5780 -7902 5814 -7883
rect 5780 -7970 5814 -7968
rect 5780 -8006 5814 -8004
rect 5780 -8091 5814 -8072
rect 6038 -7902 6072 -7883
rect 6038 -7970 6072 -7968
rect 6038 -8006 6072 -8004
rect 6038 -8091 6072 -8072
rect 6296 -7902 6330 -7883
rect 6296 -7970 6330 -7968
rect 6296 -8006 6330 -8004
rect 6296 -8091 6330 -8072
rect 6554 -7902 6588 -7883
rect 6554 -7970 6588 -7968
rect 6554 -8006 6588 -8004
rect 6554 -8091 6588 -8072
rect 6812 -7902 6846 -7883
rect 6812 -7970 6846 -7968
rect 6812 -8006 6846 -8004
rect 6812 -8091 6846 -8072
rect 7006 -7902 7040 -7883
rect 7006 -7970 7040 -7968
rect 7006 -8006 7040 -8004
rect 7006 -8091 7040 -8072
rect 7264 -7902 7298 -7883
rect 7264 -7970 7298 -7968
rect 7264 -8006 7298 -8004
rect 7264 -8091 7298 -8072
rect 7522 -7902 7556 -7883
rect 7522 -7970 7556 -7968
rect 7522 -8006 7556 -8004
rect 7522 -8091 7556 -8072
rect 7780 -7902 7814 -7883
rect 7780 -7970 7814 -7968
rect 7780 -8006 7814 -8004
rect 7780 -8091 7814 -8072
rect 7974 -7902 8008 -7883
rect 7974 -7970 8008 -7968
rect 7974 -8006 8008 -8004
rect 7974 -8091 8008 -8072
rect 8232 -7902 8266 -7883
rect 8232 -7970 8266 -7968
rect 8232 -8006 8266 -8004
rect 8232 -8091 8266 -8072
rect 8490 -7902 8524 -7883
rect 8490 -7970 8524 -7968
rect 8490 -8006 8524 -8004
rect 8490 -8091 8524 -8072
rect 8748 -7902 8782 -7883
rect 8748 -7970 8782 -7968
rect 8748 -8006 8782 -8004
rect 8748 -8091 8782 -8072
rect 9006 -7902 9040 -7883
rect 9006 -7970 9040 -7968
rect 9006 -8006 9040 -8004
rect 9006 -8091 9040 -8072
rect 9200 -7902 9234 -7883
rect 9200 -7970 9234 -7968
rect 9200 -8006 9234 -8004
rect 9200 -8091 9234 -8072
rect 9458 -7902 9492 -7883
rect 9458 -7970 9492 -7968
rect 9458 -8006 9492 -8004
rect 9458 -8091 9492 -8072
rect 9573 -7884 9607 -7858
rect 13931 -7858 13932 -7812
rect 14092 -7840 14139 -7806
rect 14175 -7840 14209 -7806
rect 14245 -7840 14292 -7806
rect 14543 -7840 14590 -7806
rect 14626 -7840 14660 -7806
rect 14696 -7840 14743 -7806
rect 14801 -7840 14848 -7806
rect 14884 -7840 14918 -7806
rect 14954 -7840 15001 -7806
rect 15059 -7840 15106 -7806
rect 15142 -7840 15176 -7806
rect 15212 -7840 15259 -7806
rect 15317 -7840 15364 -7806
rect 15400 -7840 15434 -7806
rect 15470 -7840 15517 -7806
rect 15769 -7840 15816 -7806
rect 15852 -7840 15886 -7806
rect 15922 -7840 15969 -7806
rect 16027 -7840 16074 -7806
rect 16110 -7840 16144 -7806
rect 16180 -7840 16227 -7806
rect 16285 -7840 16332 -7806
rect 16368 -7840 16402 -7806
rect 16438 -7840 16485 -7806
rect 16737 -7840 16784 -7806
rect 16820 -7840 16854 -7806
rect 16890 -7840 16937 -7806
rect 16995 -7840 17042 -7806
rect 17078 -7840 17112 -7806
rect 17148 -7840 17195 -7806
rect 17253 -7840 17300 -7806
rect 17336 -7840 17370 -7806
rect 17406 -7840 17453 -7806
rect 17511 -7840 17558 -7806
rect 17594 -7840 17628 -7806
rect 17664 -7840 17711 -7806
rect 17963 -7840 18010 -7806
rect 18046 -7840 18080 -7806
rect 18116 -7840 18163 -7806
rect 18290 -7812 18324 -7790
rect 9573 -7956 9607 -7926
rect 9573 -8028 9607 -7994
rect 5248 -8134 5249 -8096
rect 5214 -8164 5249 -8134
rect 5248 -8206 5249 -8164
rect 5214 -8232 5249 -8206
rect 5248 -8278 5249 -8232
rect 5214 -8300 5249 -8278
rect 5248 -8350 5249 -8300
rect 5214 -8368 5249 -8350
rect 5248 -8402 5249 -8368
rect 9573 -8096 9607 -8062
rect 9688 -7902 9722 -7883
rect 9688 -7970 9722 -7968
rect 9688 -8006 9722 -8004
rect 9688 -8091 9722 -8072
rect 9946 -7902 9980 -7883
rect 9946 -7970 9980 -7968
rect 9946 -8006 9980 -8004
rect 9946 -8091 9980 -8072
rect 10140 -7902 10174 -7883
rect 10140 -7970 10174 -7968
rect 10140 -8006 10174 -8004
rect 10140 -8091 10174 -8072
rect 10398 -7902 10432 -7883
rect 10398 -7970 10432 -7968
rect 10398 -8006 10432 -8004
rect 10398 -8091 10432 -8072
rect 10656 -7902 10690 -7883
rect 10656 -7970 10690 -7968
rect 10656 -8006 10690 -8004
rect 10656 -8091 10690 -8072
rect 10914 -7902 10948 -7883
rect 10914 -7970 10948 -7968
rect 10914 -8006 10948 -8004
rect 10914 -8091 10948 -8072
rect 11172 -7902 11206 -7883
rect 11172 -7970 11206 -7968
rect 11172 -8006 11206 -8004
rect 11172 -8091 11206 -8072
rect 11366 -7902 11400 -7883
rect 11366 -7970 11400 -7968
rect 11366 -8006 11400 -8004
rect 11366 -8091 11400 -8072
rect 11624 -7902 11658 -7883
rect 11624 -7970 11658 -7968
rect 11624 -8006 11658 -8004
rect 11624 -8091 11658 -8072
rect 11882 -7902 11916 -7883
rect 11882 -7970 11916 -7968
rect 11882 -8006 11916 -8004
rect 11882 -8091 11916 -8072
rect 12140 -7902 12174 -7883
rect 12140 -7970 12174 -7968
rect 12140 -8006 12174 -8004
rect 12140 -8091 12174 -8072
rect 12334 -7902 12368 -7883
rect 12334 -7970 12368 -7968
rect 12334 -8006 12368 -8004
rect 12334 -8091 12368 -8072
rect 12592 -7902 12626 -7883
rect 12592 -7970 12626 -7968
rect 12592 -8006 12626 -8004
rect 12592 -8091 12626 -8072
rect 12850 -7902 12884 -7883
rect 12850 -7970 12884 -7968
rect 12850 -8006 12884 -8004
rect 12850 -8091 12884 -8072
rect 13108 -7902 13142 -7883
rect 13108 -7970 13142 -7968
rect 13108 -8006 13142 -8004
rect 13108 -8091 13142 -8072
rect 13366 -7902 13400 -7883
rect 13366 -7970 13400 -7968
rect 13366 -8006 13400 -8004
rect 13366 -8091 13400 -8072
rect 13560 -7902 13594 -7883
rect 13560 -7970 13594 -7968
rect 13560 -8006 13594 -8004
rect 13560 -8091 13594 -8072
rect 13818 -7902 13852 -7883
rect 13818 -7970 13852 -7968
rect 13818 -8006 13852 -8004
rect 13818 -8091 13852 -8072
rect 13931 -7884 13966 -7858
rect 13931 -7926 13932 -7884
rect 13931 -7956 13966 -7926
rect 13931 -7994 13932 -7956
rect 13931 -8028 13966 -7994
rect 13931 -8062 13932 -8028
rect 9573 -8164 9607 -8134
rect 9573 -8232 9607 -8206
rect 9573 -8300 9607 -8278
rect 9573 -8368 9607 -8350
rect 13931 -8096 13966 -8062
rect 14046 -7902 14080 -7883
rect 14046 -7970 14080 -7968
rect 14046 -8006 14080 -8004
rect 14046 -8091 14080 -8072
rect 14304 -7902 14338 -7883
rect 14304 -7970 14338 -7968
rect 14304 -8006 14338 -8004
rect 14304 -8091 14338 -8072
rect 14497 -7902 14531 -7883
rect 14497 -7970 14531 -7968
rect 14497 -8006 14531 -8004
rect 14497 -8091 14531 -8072
rect 14755 -7902 14789 -7883
rect 14755 -7970 14789 -7968
rect 14755 -8006 14789 -8004
rect 14755 -8091 14789 -8072
rect 15013 -7902 15047 -7883
rect 15013 -7970 15047 -7968
rect 15013 -8006 15047 -8004
rect 15013 -8091 15047 -8072
rect 15271 -7902 15305 -7883
rect 15271 -7970 15305 -7968
rect 15271 -8006 15305 -8004
rect 15271 -8091 15305 -8072
rect 15529 -7902 15563 -7883
rect 15529 -7970 15563 -7968
rect 15529 -8006 15563 -8004
rect 15529 -8091 15563 -8072
rect 15723 -7902 15757 -7883
rect 15723 -7970 15757 -7968
rect 15723 -8006 15757 -8004
rect 15723 -8091 15757 -8072
rect 15981 -7902 16015 -7883
rect 15981 -7970 16015 -7968
rect 15981 -8006 16015 -8004
rect 15981 -8091 16015 -8072
rect 16239 -7902 16273 -7883
rect 16239 -7970 16273 -7968
rect 16239 -8006 16273 -8004
rect 16239 -8091 16273 -8072
rect 16497 -7902 16531 -7883
rect 16497 -7970 16531 -7968
rect 16497 -8006 16531 -8004
rect 16497 -8091 16531 -8072
rect 16691 -7902 16725 -7883
rect 16691 -7970 16725 -7968
rect 16691 -8006 16725 -8004
rect 16691 -8091 16725 -8072
rect 16949 -7902 16983 -7883
rect 16949 -7970 16983 -7968
rect 16949 -8006 16983 -8004
rect 16949 -8091 16983 -8072
rect 17207 -7902 17241 -7883
rect 17207 -7970 17241 -7968
rect 17207 -8006 17241 -8004
rect 17207 -8091 17241 -8072
rect 17465 -7902 17499 -7883
rect 17465 -7970 17499 -7968
rect 17465 -8006 17499 -8004
rect 17465 -8091 17499 -8072
rect 17723 -7902 17757 -7883
rect 17723 -7970 17757 -7968
rect 17723 -8006 17757 -8004
rect 17723 -8091 17757 -8072
rect 17917 -7902 17951 -7883
rect 17917 -7970 17951 -7968
rect 17917 -8006 17951 -8004
rect 17917 -8091 17951 -8072
rect 18175 -7902 18209 -7883
rect 18175 -7970 18209 -7968
rect 18175 -8006 18209 -8004
rect 18175 -8091 18209 -8072
rect 18290 -7884 18324 -7858
rect 18290 -7956 18324 -7926
rect 18290 -8028 18324 -7994
rect 13931 -8134 13932 -8096
rect 13931 -8164 13966 -8134
rect 13931 -8206 13932 -8164
rect 13931 -8232 13966 -8206
rect 13931 -8278 13932 -8232
rect 13931 -8300 13966 -8278
rect 13931 -8350 13932 -8300
rect 13931 -8368 13966 -8350
rect 13931 -8402 13932 -8368
rect 18290 -8096 18324 -8062
rect 18290 -8164 18324 -8134
rect 18290 -8232 18324 -8206
rect 18290 -8300 18324 -8278
rect 18290 -8368 18324 -8350
rect 890 -8422 977 -8402
rect 856 -8436 977 -8422
rect 1011 -8436 1045 -8402
rect 1079 -8436 1113 -8402
rect 1147 -8436 1181 -8402
rect 1215 -8436 1249 -8402
rect 1283 -8436 1317 -8402
rect 1351 -8436 1385 -8402
rect 1419 -8436 1453 -8402
rect 1487 -8436 1521 -8402
rect 1555 -8436 1589 -8402
rect 1623 -8436 1657 -8402
rect 1691 -8436 1725 -8402
rect 1759 -8436 1793 -8402
rect 1827 -8436 1861 -8402
rect 1895 -8436 1929 -8402
rect 1963 -8436 1997 -8402
rect 2031 -8436 2065 -8402
rect 2099 -8436 2133 -8402
rect 2167 -8436 2201 -8402
rect 2235 -8436 2269 -8402
rect 2303 -8436 2337 -8402
rect 2371 -8436 2405 -8402
rect 2439 -8436 2473 -8402
rect 2507 -8436 2541 -8402
rect 2575 -8436 2609 -8402
rect 2643 -8436 2677 -8402
rect 2711 -8436 2745 -8402
rect 2779 -8436 2813 -8402
rect 2847 -8436 2881 -8402
rect 2915 -8436 2949 -8402
rect 2983 -8436 3017 -8402
rect 3051 -8436 3085 -8402
rect 3119 -8436 3153 -8402
rect 3187 -8436 3221 -8402
rect 3255 -8436 3289 -8402
rect 3323 -8436 3357 -8402
rect 3391 -8436 3425 -8402
rect 3459 -8436 3493 -8402
rect 3527 -8436 3561 -8402
rect 3595 -8436 3629 -8402
rect 3663 -8436 3697 -8402
rect 3731 -8436 3765 -8402
rect 3799 -8436 3833 -8402
rect 3867 -8436 3901 -8402
rect 3935 -8436 3969 -8402
rect 4003 -8436 4037 -8402
rect 4071 -8436 4105 -8402
rect 4139 -8436 4173 -8402
rect 4207 -8436 4241 -8402
rect 4275 -8436 4309 -8402
rect 4343 -8436 4377 -8402
rect 4411 -8436 4445 -8402
rect 4479 -8436 4513 -8402
rect 4547 -8436 4581 -8402
rect 4615 -8436 4649 -8402
rect 4683 -8436 4717 -8402
rect 4751 -8436 4785 -8402
rect 4819 -8436 4853 -8402
rect 4887 -8436 4921 -8402
rect 4955 -8436 4989 -8402
rect 5023 -8436 5057 -8402
rect 5091 -8422 5214 -8402
rect 5248 -8422 5372 -8402
rect 5091 -8436 5372 -8422
rect 5406 -8436 5440 -8402
rect 5474 -8436 5508 -8402
rect 5542 -8436 5576 -8402
rect 5610 -8436 5644 -8402
rect 5678 -8436 5712 -8402
rect 5746 -8436 5780 -8402
rect 5814 -8436 5848 -8402
rect 5882 -8436 5916 -8402
rect 5950 -8436 5984 -8402
rect 6018 -8436 6052 -8402
rect 6086 -8436 6120 -8402
rect 6154 -8436 6188 -8402
rect 6222 -8436 6256 -8402
rect 6290 -8436 6324 -8402
rect 6358 -8436 6392 -8402
rect 6426 -8436 6460 -8402
rect 6494 -8436 6528 -8402
rect 6562 -8436 6596 -8402
rect 6630 -8436 6664 -8402
rect 6698 -8436 6732 -8402
rect 6766 -8436 6800 -8402
rect 6834 -8436 6868 -8402
rect 6902 -8436 6936 -8402
rect 6970 -8436 7004 -8402
rect 7038 -8436 7072 -8402
rect 7106 -8436 7140 -8402
rect 7174 -8436 7208 -8402
rect 7242 -8436 7276 -8402
rect 7310 -8436 7344 -8402
rect 7378 -8436 7412 -8402
rect 7446 -8436 7480 -8402
rect 7514 -8436 7548 -8402
rect 7582 -8436 7616 -8402
rect 7650 -8436 7684 -8402
rect 7718 -8436 7752 -8402
rect 7786 -8436 7820 -8402
rect 7854 -8436 7888 -8402
rect 7922 -8436 7956 -8402
rect 7990 -8436 8024 -8402
rect 8058 -8436 8092 -8402
rect 8126 -8436 8160 -8402
rect 8194 -8436 8228 -8402
rect 8262 -8436 8296 -8402
rect 8330 -8436 8364 -8402
rect 8398 -8436 8432 -8402
rect 8466 -8436 8500 -8402
rect 8534 -8436 8568 -8402
rect 8602 -8436 8636 -8402
rect 8670 -8436 8704 -8402
rect 8738 -8436 8772 -8402
rect 8806 -8436 8840 -8402
rect 8874 -8436 8908 -8402
rect 8942 -8436 8976 -8402
rect 9010 -8436 9044 -8402
rect 9078 -8436 9112 -8402
rect 9146 -8436 9180 -8402
rect 9214 -8436 9248 -8402
rect 9282 -8436 9316 -8402
rect 9350 -8436 9384 -8402
rect 9418 -8436 9452 -8402
rect 9486 -8422 9573 -8402
rect 9607 -8422 9694 -8402
rect 9486 -8436 9694 -8422
rect 9728 -8436 9762 -8402
rect 9796 -8436 9830 -8402
rect 9864 -8436 9898 -8402
rect 9932 -8436 9966 -8402
rect 10000 -8436 10034 -8402
rect 10068 -8436 10102 -8402
rect 10136 -8436 10170 -8402
rect 10204 -8436 10238 -8402
rect 10272 -8436 10306 -8402
rect 10340 -8436 10374 -8402
rect 10408 -8436 10442 -8402
rect 10476 -8436 10510 -8402
rect 10544 -8436 10578 -8402
rect 10612 -8436 10646 -8402
rect 10680 -8436 10714 -8402
rect 10748 -8436 10782 -8402
rect 10816 -8436 10850 -8402
rect 10884 -8436 10918 -8402
rect 10952 -8436 10986 -8402
rect 11020 -8436 11054 -8402
rect 11088 -8436 11122 -8402
rect 11156 -8436 11190 -8402
rect 11224 -8436 11258 -8402
rect 11292 -8436 11326 -8402
rect 11360 -8436 11394 -8402
rect 11428 -8436 11462 -8402
rect 11496 -8436 11530 -8402
rect 11564 -8436 11598 -8402
rect 11632 -8436 11666 -8402
rect 11700 -8436 11734 -8402
rect 11768 -8436 11802 -8402
rect 11836 -8436 11870 -8402
rect 11904 -8436 11938 -8402
rect 11972 -8436 12006 -8402
rect 12040 -8436 12074 -8402
rect 12108 -8436 12142 -8402
rect 12176 -8436 12210 -8402
rect 12244 -8436 12278 -8402
rect 12312 -8436 12346 -8402
rect 12380 -8436 12414 -8402
rect 12448 -8436 12482 -8402
rect 12516 -8436 12550 -8402
rect 12584 -8436 12618 -8402
rect 12652 -8436 12686 -8402
rect 12720 -8436 12754 -8402
rect 12788 -8436 12822 -8402
rect 12856 -8436 12890 -8402
rect 12924 -8436 12958 -8402
rect 12992 -8436 13026 -8402
rect 13060 -8436 13094 -8402
rect 13128 -8436 13162 -8402
rect 13196 -8436 13230 -8402
rect 13264 -8436 13298 -8402
rect 13332 -8436 13366 -8402
rect 13400 -8436 13434 -8402
rect 13468 -8436 13502 -8402
rect 13536 -8436 13570 -8402
rect 13604 -8436 13638 -8402
rect 13672 -8436 13706 -8402
rect 13740 -8436 13774 -8402
rect 13808 -8422 13932 -8402
rect 13966 -8422 14089 -8402
rect 13808 -8436 14089 -8422
rect 14123 -8436 14157 -8402
rect 14191 -8436 14225 -8402
rect 14259 -8436 14293 -8402
rect 14327 -8436 14361 -8402
rect 14395 -8436 14429 -8402
rect 14463 -8436 14497 -8402
rect 14531 -8436 14565 -8402
rect 14599 -8436 14633 -8402
rect 14667 -8436 14701 -8402
rect 14735 -8436 14769 -8402
rect 14803 -8436 14837 -8402
rect 14871 -8436 14905 -8402
rect 14939 -8436 14973 -8402
rect 15007 -8436 15041 -8402
rect 15075 -8436 15109 -8402
rect 15143 -8436 15177 -8402
rect 15211 -8436 15245 -8402
rect 15279 -8436 15313 -8402
rect 15347 -8436 15381 -8402
rect 15415 -8436 15449 -8402
rect 15483 -8436 15517 -8402
rect 15551 -8436 15585 -8402
rect 15619 -8436 15653 -8402
rect 15687 -8436 15721 -8402
rect 15755 -8436 15789 -8402
rect 15823 -8436 15857 -8402
rect 15891 -8436 15925 -8402
rect 15959 -8436 15993 -8402
rect 16027 -8436 16061 -8402
rect 16095 -8436 16129 -8402
rect 16163 -8436 16197 -8402
rect 16231 -8436 16265 -8402
rect 16299 -8436 16333 -8402
rect 16367 -8436 16401 -8402
rect 16435 -8436 16469 -8402
rect 16503 -8436 16537 -8402
rect 16571 -8436 16605 -8402
rect 16639 -8436 16673 -8402
rect 16707 -8436 16741 -8402
rect 16775 -8436 16809 -8402
rect 16843 -8436 16877 -8402
rect 16911 -8436 16945 -8402
rect 16979 -8436 17013 -8402
rect 17047 -8436 17081 -8402
rect 17115 -8436 17149 -8402
rect 17183 -8436 17217 -8402
rect 17251 -8436 17285 -8402
rect 17319 -8436 17353 -8402
rect 17387 -8436 17421 -8402
rect 17455 -8436 17489 -8402
rect 17523 -8436 17557 -8402
rect 17591 -8436 17625 -8402
rect 17659 -8436 17693 -8402
rect 17727 -8436 17761 -8402
rect 17795 -8436 17829 -8402
rect 17863 -8436 17897 -8402
rect 17931 -8436 17965 -8402
rect 17999 -8436 18033 -8402
rect 18067 -8436 18101 -8402
rect 18135 -8436 18169 -8402
rect 18203 -8422 18290 -8402
rect 18203 -8436 18324 -8422
rect 856 -8504 890 -8494
rect 856 -8572 890 -8566
rect 856 -8640 890 -8638
rect 856 -8676 890 -8674
rect 856 -8748 890 -8742
rect 856 -8820 890 -8810
rect 5248 -8494 5249 -8436
rect 5214 -8504 5249 -8494
rect 5248 -8566 5249 -8504
rect 5214 -8572 5249 -8566
rect 5248 -8638 5249 -8572
rect 5214 -8640 5249 -8638
rect 5248 -8674 5249 -8640
rect 5214 -8676 5249 -8674
rect 5248 -8742 5249 -8676
rect 5214 -8748 5249 -8742
rect 5248 -8810 5249 -8748
rect 5214 -8820 5249 -8810
rect 856 -8892 890 -8878
rect 856 -8964 890 -8946
rect 856 -9036 890 -9014
rect 971 -8846 1005 -8827
rect 971 -8914 1005 -8912
rect 971 -8950 1005 -8948
rect 971 -9035 1005 -9016
rect 1229 -8846 1263 -8827
rect 1229 -8914 1263 -8912
rect 1229 -8950 1263 -8948
rect 1229 -9035 1263 -9016
rect 1423 -8846 1457 -8827
rect 1423 -8914 1457 -8912
rect 1423 -8950 1457 -8948
rect 1423 -9035 1457 -9016
rect 1681 -8846 1715 -8827
rect 1681 -8914 1715 -8912
rect 1681 -8950 1715 -8948
rect 1681 -9035 1715 -9016
rect 1939 -8846 1973 -8827
rect 1939 -8914 1973 -8912
rect 1939 -8950 1973 -8948
rect 1939 -9035 1973 -9016
rect 2197 -8846 2231 -8827
rect 2197 -8914 2231 -8912
rect 2197 -8950 2231 -8948
rect 2197 -9035 2231 -9016
rect 2455 -8846 2489 -8827
rect 2455 -8914 2489 -8912
rect 2455 -8950 2489 -8948
rect 2455 -9035 2489 -9016
rect 2649 -8846 2683 -8827
rect 2649 -8914 2683 -8912
rect 2649 -8950 2683 -8948
rect 2649 -9035 2683 -9016
rect 2907 -8846 2941 -8827
rect 2907 -8914 2941 -8912
rect 2907 -8950 2941 -8948
rect 2907 -9035 2941 -9016
rect 3165 -8846 3199 -8827
rect 3165 -8914 3199 -8912
rect 3165 -8950 3199 -8948
rect 3165 -9035 3199 -9016
rect 3423 -8846 3457 -8827
rect 3423 -8914 3457 -8912
rect 3423 -8950 3457 -8948
rect 3423 -9035 3457 -9016
rect 3617 -8846 3651 -8827
rect 3617 -8914 3651 -8912
rect 3617 -8950 3651 -8948
rect 3617 -9035 3651 -9016
rect 3875 -8846 3909 -8827
rect 3875 -8914 3909 -8912
rect 3875 -8950 3909 -8948
rect 3875 -9035 3909 -9016
rect 4133 -8846 4167 -8827
rect 4133 -8914 4167 -8912
rect 4133 -8950 4167 -8948
rect 4133 -9035 4167 -9016
rect 4391 -8846 4425 -8827
rect 4391 -8914 4425 -8912
rect 4391 -8950 4425 -8948
rect 4391 -9035 4425 -9016
rect 4649 -8846 4683 -8827
rect 4649 -8914 4683 -8912
rect 4649 -8950 4683 -8948
rect 4649 -9035 4683 -9016
rect 4842 -8846 4876 -8827
rect 4842 -8914 4876 -8912
rect 4842 -8950 4876 -8948
rect 4842 -9035 4876 -9016
rect 5100 -8846 5134 -8827
rect 5100 -8914 5134 -8912
rect 5100 -8950 5134 -8948
rect 5100 -9035 5134 -9016
rect 5248 -8878 5249 -8820
rect 9573 -8504 9607 -8494
rect 9573 -8572 9607 -8566
rect 9573 -8640 9607 -8638
rect 9573 -8676 9607 -8674
rect 9573 -8748 9607 -8742
rect 9573 -8820 9607 -8810
rect 5214 -8892 5249 -8878
rect 5248 -8946 5249 -8892
rect 5214 -8964 5249 -8946
rect 5248 -9014 5249 -8964
rect 856 -9192 890 -9070
rect 5214 -9036 5249 -9014
rect 5328 -8846 5362 -8827
rect 5328 -8914 5362 -8912
rect 5328 -8950 5362 -8948
rect 5328 -9035 5362 -9016
rect 5586 -8846 5620 -8827
rect 5586 -8914 5620 -8912
rect 5586 -8950 5620 -8948
rect 5586 -9035 5620 -9016
rect 5780 -8846 5814 -8827
rect 5780 -8914 5814 -8912
rect 5780 -8950 5814 -8948
rect 5780 -9035 5814 -9016
rect 6038 -8846 6072 -8827
rect 6038 -8914 6072 -8912
rect 6038 -8950 6072 -8948
rect 6038 -9035 6072 -9016
rect 6296 -8846 6330 -8827
rect 6296 -8914 6330 -8912
rect 6296 -8950 6330 -8948
rect 6296 -9035 6330 -9016
rect 6554 -8846 6588 -8827
rect 6554 -8914 6588 -8912
rect 6554 -8950 6588 -8948
rect 6554 -9035 6588 -9016
rect 6812 -8846 6846 -8827
rect 6812 -8914 6846 -8912
rect 6812 -8950 6846 -8948
rect 6812 -9035 6846 -9016
rect 7006 -8846 7040 -8827
rect 7006 -8914 7040 -8912
rect 7006 -8950 7040 -8948
rect 7006 -9035 7040 -9016
rect 7264 -8846 7298 -8827
rect 7264 -8914 7298 -8912
rect 7264 -8950 7298 -8948
rect 7264 -9035 7298 -9016
rect 7522 -8846 7556 -8827
rect 7522 -8914 7556 -8912
rect 7522 -8950 7556 -8948
rect 7522 -9035 7556 -9016
rect 7780 -8846 7814 -8827
rect 7780 -8914 7814 -8912
rect 7780 -8950 7814 -8948
rect 7780 -9035 7814 -9016
rect 7974 -8846 8008 -8827
rect 7974 -8914 8008 -8912
rect 7974 -8950 8008 -8948
rect 7974 -9035 8008 -9016
rect 8232 -8846 8266 -8827
rect 8232 -8914 8266 -8912
rect 8232 -8950 8266 -8948
rect 8232 -9035 8266 -9016
rect 8490 -8846 8524 -8827
rect 8490 -8914 8524 -8912
rect 8490 -8950 8524 -8948
rect 8490 -9035 8524 -9016
rect 8748 -8846 8782 -8827
rect 8748 -8914 8782 -8912
rect 8748 -8950 8782 -8948
rect 8748 -9035 8782 -9016
rect 9006 -8846 9040 -8827
rect 9006 -8914 9040 -8912
rect 9006 -8950 9040 -8948
rect 9006 -9035 9040 -9016
rect 9200 -8846 9234 -8827
rect 9200 -8914 9234 -8912
rect 9200 -8950 9234 -8948
rect 9200 -9035 9234 -9016
rect 9458 -8846 9492 -8827
rect 9458 -8914 9492 -8912
rect 9458 -8950 9492 -8948
rect 9458 -9035 9492 -9016
rect 13931 -8494 13932 -8436
rect 13931 -8504 13966 -8494
rect 13931 -8566 13932 -8504
rect 13931 -8572 13966 -8566
rect 13931 -8638 13932 -8572
rect 13931 -8640 13966 -8638
rect 13931 -8674 13932 -8640
rect 13931 -8676 13966 -8674
rect 13931 -8742 13932 -8676
rect 13931 -8748 13966 -8742
rect 13931 -8810 13932 -8748
rect 13931 -8820 13966 -8810
rect 9573 -8892 9607 -8878
rect 9573 -8964 9607 -8946
rect 5248 -9070 5249 -9036
rect 1017 -9112 1064 -9078
rect 1100 -9112 1134 -9078
rect 1170 -9112 1217 -9078
rect 1469 -9112 1516 -9078
rect 1552 -9112 1586 -9078
rect 1622 -9112 1669 -9078
rect 1727 -9112 1774 -9078
rect 1810 -9112 1844 -9078
rect 1880 -9112 1927 -9078
rect 1985 -9112 2032 -9078
rect 2068 -9112 2102 -9078
rect 2138 -9112 2185 -9078
rect 2243 -9112 2290 -9078
rect 2326 -9112 2360 -9078
rect 2396 -9112 2443 -9078
rect 2695 -9112 2742 -9078
rect 2778 -9112 2812 -9078
rect 2848 -9112 2895 -9078
rect 2953 -9112 3000 -9078
rect 3036 -9112 3070 -9078
rect 3106 -9112 3153 -9078
rect 3211 -9112 3258 -9078
rect 3294 -9112 3328 -9078
rect 3364 -9112 3411 -9078
rect 3663 -9112 3710 -9078
rect 3746 -9112 3780 -9078
rect 3816 -9112 3863 -9078
rect 3921 -9112 3968 -9078
rect 4004 -9112 4038 -9078
rect 4074 -9112 4121 -9078
rect 4179 -9112 4226 -9078
rect 4262 -9112 4296 -9078
rect 4332 -9112 4379 -9078
rect 4437 -9112 4484 -9078
rect 4520 -9112 4554 -9078
rect 4590 -9112 4637 -9078
rect 4888 -9112 4935 -9078
rect 4971 -9112 5005 -9078
rect 5041 -9112 5088 -9078
rect 5214 -9192 5249 -9070
rect 9573 -9036 9607 -9014
rect 9688 -8846 9722 -8827
rect 9688 -8914 9722 -8912
rect 9688 -8950 9722 -8948
rect 9688 -9035 9722 -9016
rect 9946 -8846 9980 -8827
rect 9946 -8914 9980 -8912
rect 9946 -8950 9980 -8948
rect 9946 -9035 9980 -9016
rect 10140 -8846 10174 -8827
rect 10140 -8914 10174 -8912
rect 10140 -8950 10174 -8948
rect 10140 -9035 10174 -9016
rect 10398 -8846 10432 -8827
rect 10398 -8914 10432 -8912
rect 10398 -8950 10432 -8948
rect 10398 -9035 10432 -9016
rect 10656 -8846 10690 -8827
rect 10656 -8914 10690 -8912
rect 10656 -8950 10690 -8948
rect 10656 -9035 10690 -9016
rect 10914 -8846 10948 -8827
rect 10914 -8914 10948 -8912
rect 10914 -8950 10948 -8948
rect 10914 -9035 10948 -9016
rect 11172 -8846 11206 -8827
rect 11172 -8914 11206 -8912
rect 11172 -8950 11206 -8948
rect 11172 -9035 11206 -9016
rect 11366 -8846 11400 -8827
rect 11366 -8914 11400 -8912
rect 11366 -8950 11400 -8948
rect 11366 -9035 11400 -9016
rect 11624 -8846 11658 -8827
rect 11624 -8914 11658 -8912
rect 11624 -8950 11658 -8948
rect 11624 -9035 11658 -9016
rect 11882 -8846 11916 -8827
rect 11882 -8914 11916 -8912
rect 11882 -8950 11916 -8948
rect 11882 -9035 11916 -9016
rect 12140 -8846 12174 -8827
rect 12140 -8914 12174 -8912
rect 12140 -8950 12174 -8948
rect 12140 -9035 12174 -9016
rect 12334 -8846 12368 -8827
rect 12334 -8914 12368 -8912
rect 12334 -8950 12368 -8948
rect 12334 -9035 12368 -9016
rect 12592 -8846 12626 -8827
rect 12592 -8914 12626 -8912
rect 12592 -8950 12626 -8948
rect 12592 -9035 12626 -9016
rect 12850 -8846 12884 -8827
rect 12850 -8914 12884 -8912
rect 12850 -8950 12884 -8948
rect 12850 -9035 12884 -9016
rect 13108 -8846 13142 -8827
rect 13108 -8914 13142 -8912
rect 13108 -8950 13142 -8948
rect 13108 -9035 13142 -9016
rect 13366 -8846 13400 -8827
rect 13366 -8914 13400 -8912
rect 13366 -8950 13400 -8948
rect 13366 -9035 13400 -9016
rect 13560 -8846 13594 -8827
rect 13560 -8914 13594 -8912
rect 13560 -8950 13594 -8948
rect 13560 -9035 13594 -9016
rect 13818 -8846 13852 -8827
rect 13818 -8914 13852 -8912
rect 13818 -8950 13852 -8948
rect 13818 -9035 13852 -9016
rect 13931 -8878 13932 -8820
rect 18290 -8504 18324 -8494
rect 18290 -8572 18324 -8566
rect 18290 -8640 18324 -8638
rect 18290 -8676 18324 -8674
rect 18290 -8748 18324 -8742
rect 18290 -8820 18324 -8810
rect 13931 -8892 13966 -8878
rect 13931 -8946 13932 -8892
rect 13931 -8964 13966 -8946
rect 13931 -9014 13932 -8964
rect 5374 -9112 5421 -9078
rect 5457 -9112 5491 -9078
rect 5527 -9112 5574 -9078
rect 5826 -9112 5873 -9078
rect 5909 -9112 5943 -9078
rect 5979 -9112 6026 -9078
rect 6084 -9112 6131 -9078
rect 6167 -9112 6201 -9078
rect 6237 -9112 6284 -9078
rect 6342 -9112 6389 -9078
rect 6425 -9112 6459 -9078
rect 6495 -9112 6542 -9078
rect 6600 -9112 6647 -9078
rect 6683 -9112 6717 -9078
rect 6753 -9112 6800 -9078
rect 7052 -9112 7099 -9078
rect 7135 -9112 7169 -9078
rect 7205 -9112 7252 -9078
rect 7310 -9112 7357 -9078
rect 7393 -9112 7427 -9078
rect 7463 -9112 7510 -9078
rect 7568 -9112 7615 -9078
rect 7651 -9112 7685 -9078
rect 7721 -9112 7768 -9078
rect 8020 -9112 8067 -9078
rect 8103 -9112 8137 -9078
rect 8173 -9112 8220 -9078
rect 8278 -9112 8325 -9078
rect 8361 -9112 8395 -9078
rect 8431 -9112 8478 -9078
rect 8536 -9112 8583 -9078
rect 8619 -9112 8653 -9078
rect 8689 -9112 8736 -9078
rect 8794 -9112 8841 -9078
rect 8877 -9112 8911 -9078
rect 8947 -9112 8994 -9078
rect 9246 -9112 9293 -9078
rect 9329 -9112 9363 -9078
rect 9399 -9112 9446 -9078
rect 9573 -9192 9607 -9070
rect 13931 -9036 13966 -9014
rect 14046 -8846 14080 -8827
rect 14046 -8914 14080 -8912
rect 14046 -8950 14080 -8948
rect 14046 -9035 14080 -9016
rect 14304 -8846 14338 -8827
rect 14304 -8914 14338 -8912
rect 14304 -8950 14338 -8948
rect 14304 -9035 14338 -9016
rect 14497 -8846 14531 -8827
rect 14497 -8914 14531 -8912
rect 14497 -8950 14531 -8948
rect 14497 -9035 14531 -9016
rect 14755 -8846 14789 -8827
rect 14755 -8914 14789 -8912
rect 14755 -8950 14789 -8948
rect 14755 -9035 14789 -9016
rect 15013 -8846 15047 -8827
rect 15013 -8914 15047 -8912
rect 15013 -8950 15047 -8948
rect 15013 -9035 15047 -9016
rect 15271 -8846 15305 -8827
rect 15271 -8914 15305 -8912
rect 15271 -8950 15305 -8948
rect 15271 -9035 15305 -9016
rect 15529 -8846 15563 -8827
rect 15529 -8914 15563 -8912
rect 15529 -8950 15563 -8948
rect 15529 -9035 15563 -9016
rect 15723 -8846 15757 -8827
rect 15723 -8914 15757 -8912
rect 15723 -8950 15757 -8948
rect 15723 -9035 15757 -9016
rect 15981 -8846 16015 -8827
rect 15981 -8914 16015 -8912
rect 15981 -8950 16015 -8948
rect 15981 -9035 16015 -9016
rect 16239 -8846 16273 -8827
rect 16239 -8914 16273 -8912
rect 16239 -8950 16273 -8948
rect 16239 -9035 16273 -9016
rect 16497 -8846 16531 -8827
rect 16497 -8914 16531 -8912
rect 16497 -8950 16531 -8948
rect 16497 -9035 16531 -9016
rect 16691 -8846 16725 -8827
rect 16691 -8914 16725 -8912
rect 16691 -8950 16725 -8948
rect 16691 -9035 16725 -9016
rect 16949 -8846 16983 -8827
rect 16949 -8914 16983 -8912
rect 16949 -8950 16983 -8948
rect 16949 -9035 16983 -9016
rect 17207 -8846 17241 -8827
rect 17207 -8914 17241 -8912
rect 17207 -8950 17241 -8948
rect 17207 -9035 17241 -9016
rect 17465 -8846 17499 -8827
rect 17465 -8914 17499 -8912
rect 17465 -8950 17499 -8948
rect 17465 -9035 17499 -9016
rect 17723 -8846 17757 -8827
rect 17723 -8914 17757 -8912
rect 17723 -8950 17757 -8948
rect 17723 -9035 17757 -9016
rect 17917 -8846 17951 -8827
rect 17917 -8914 17951 -8912
rect 17917 -8950 17951 -8948
rect 17917 -9035 17951 -9016
rect 18175 -8846 18209 -8827
rect 18175 -8914 18209 -8912
rect 18175 -8950 18209 -8948
rect 18175 -9035 18209 -9016
rect 18290 -8892 18324 -8878
rect 18290 -8964 18324 -8946
rect 13931 -9070 13932 -9036
rect 9734 -9112 9781 -9078
rect 9817 -9112 9851 -9078
rect 9887 -9112 9934 -9078
rect 10186 -9112 10233 -9078
rect 10269 -9112 10303 -9078
rect 10339 -9112 10386 -9078
rect 10444 -9112 10491 -9078
rect 10527 -9112 10561 -9078
rect 10597 -9112 10644 -9078
rect 10702 -9112 10749 -9078
rect 10785 -9112 10819 -9078
rect 10855 -9112 10902 -9078
rect 10960 -9112 11007 -9078
rect 11043 -9112 11077 -9078
rect 11113 -9112 11160 -9078
rect 11412 -9112 11459 -9078
rect 11495 -9112 11529 -9078
rect 11565 -9112 11612 -9078
rect 11670 -9112 11717 -9078
rect 11753 -9112 11787 -9078
rect 11823 -9112 11870 -9078
rect 11928 -9112 11975 -9078
rect 12011 -9112 12045 -9078
rect 12081 -9112 12128 -9078
rect 12380 -9112 12427 -9078
rect 12463 -9112 12497 -9078
rect 12533 -9112 12580 -9078
rect 12638 -9112 12685 -9078
rect 12721 -9112 12755 -9078
rect 12791 -9112 12838 -9078
rect 12896 -9112 12943 -9078
rect 12979 -9112 13013 -9078
rect 13049 -9112 13096 -9078
rect 13154 -9112 13201 -9078
rect 13237 -9112 13271 -9078
rect 13307 -9112 13354 -9078
rect 13606 -9112 13653 -9078
rect 13689 -9112 13723 -9078
rect 13759 -9112 13806 -9078
rect 13931 -9192 13966 -9070
rect 18290 -9036 18324 -9014
rect 14092 -9112 14139 -9078
rect 14175 -9112 14209 -9078
rect 14245 -9112 14292 -9078
rect 14543 -9112 14590 -9078
rect 14626 -9112 14660 -9078
rect 14696 -9112 14743 -9078
rect 14801 -9112 14848 -9078
rect 14884 -9112 14918 -9078
rect 14954 -9112 15001 -9078
rect 15059 -9112 15106 -9078
rect 15142 -9112 15176 -9078
rect 15212 -9112 15259 -9078
rect 15317 -9112 15364 -9078
rect 15400 -9112 15434 -9078
rect 15470 -9112 15517 -9078
rect 15769 -9112 15816 -9078
rect 15852 -9112 15886 -9078
rect 15922 -9112 15969 -9078
rect 16027 -9112 16074 -9078
rect 16110 -9112 16144 -9078
rect 16180 -9112 16227 -9078
rect 16285 -9112 16332 -9078
rect 16368 -9112 16402 -9078
rect 16438 -9112 16485 -9078
rect 16737 -9112 16784 -9078
rect 16820 -9112 16854 -9078
rect 16890 -9112 16937 -9078
rect 16995 -9112 17042 -9078
rect 17078 -9112 17112 -9078
rect 17148 -9112 17195 -9078
rect 17253 -9112 17300 -9078
rect 17336 -9112 17370 -9078
rect 17406 -9112 17453 -9078
rect 17511 -9112 17558 -9078
rect 17594 -9112 17628 -9078
rect 17664 -9112 17711 -9078
rect 17963 -9112 18010 -9078
rect 18046 -9112 18080 -9078
rect 18116 -9112 18163 -9078
rect 18290 -9192 18324 -9070
rect 856 -9226 930 -9192
rect 964 -9226 977 -9192
rect 1036 -9226 1045 -9192
rect 1108 -9226 1113 -9192
rect 1180 -9226 1181 -9192
rect 1215 -9226 1218 -9192
rect 1283 -9226 1290 -9192
rect 1351 -9226 1362 -9192
rect 1419 -9226 1434 -9192
rect 1487 -9226 1506 -9192
rect 1555 -9226 1578 -9192
rect 1623 -9226 1650 -9192
rect 1691 -9226 1722 -9192
rect 1759 -9226 1793 -9192
rect 1828 -9226 1861 -9192
rect 1900 -9226 1929 -9192
rect 1972 -9226 1997 -9192
rect 2044 -9226 2065 -9192
rect 2116 -9226 2133 -9192
rect 2188 -9226 2201 -9192
rect 2260 -9226 2269 -9192
rect 2332 -9226 2337 -9192
rect 2404 -9226 2405 -9192
rect 2439 -9226 2442 -9192
rect 2507 -9226 2514 -9192
rect 2575 -9226 2586 -9192
rect 2643 -9226 2658 -9192
rect 2711 -9226 2730 -9192
rect 2779 -9226 2802 -9192
rect 2847 -9226 2874 -9192
rect 2915 -9226 2946 -9192
rect 2983 -9226 3017 -9192
rect 3052 -9226 3085 -9192
rect 3124 -9226 3153 -9192
rect 3196 -9226 3221 -9192
rect 3268 -9226 3289 -9192
rect 3340 -9226 3357 -9192
rect 3412 -9226 3425 -9192
rect 3484 -9226 3493 -9192
rect 3556 -9226 3561 -9192
rect 3628 -9226 3629 -9192
rect 3663 -9226 3666 -9192
rect 3731 -9226 3738 -9192
rect 3799 -9226 3810 -9192
rect 3867 -9226 3882 -9192
rect 3935 -9226 3954 -9192
rect 4003 -9226 4026 -9192
rect 4071 -9226 4098 -9192
rect 4139 -9226 4170 -9192
rect 4207 -9226 4241 -9192
rect 4276 -9226 4309 -9192
rect 4348 -9226 4377 -9192
rect 4420 -9226 4445 -9192
rect 4492 -9226 4513 -9192
rect 4564 -9226 4581 -9192
rect 4636 -9226 4649 -9192
rect 4708 -9226 4717 -9192
rect 4780 -9226 4785 -9192
rect 4852 -9226 4853 -9192
rect 4887 -9226 4890 -9192
rect 4955 -9226 4962 -9192
rect 5023 -9226 5034 -9192
rect 5091 -9226 5106 -9192
rect 5140 -9226 5323 -9192
rect 5357 -9226 5372 -9192
rect 5429 -9226 5440 -9192
rect 5501 -9226 5508 -9192
rect 5573 -9226 5576 -9192
rect 5610 -9226 5611 -9192
rect 5678 -9226 5683 -9192
rect 5746 -9226 5755 -9192
rect 5814 -9226 5827 -9192
rect 5882 -9226 5899 -9192
rect 5950 -9226 5971 -9192
rect 6018 -9226 6043 -9192
rect 6086 -9226 6115 -9192
rect 6154 -9226 6187 -9192
rect 6222 -9226 6256 -9192
rect 6293 -9226 6324 -9192
rect 6365 -9226 6392 -9192
rect 6437 -9226 6460 -9192
rect 6509 -9226 6528 -9192
rect 6581 -9226 6596 -9192
rect 6653 -9226 6664 -9192
rect 6725 -9226 6732 -9192
rect 6797 -9226 6800 -9192
rect 6834 -9226 6835 -9192
rect 6902 -9226 6907 -9192
rect 6970 -9226 6979 -9192
rect 7038 -9226 7051 -9192
rect 7106 -9226 7123 -9192
rect 7174 -9226 7195 -9192
rect 7242 -9226 7267 -9192
rect 7310 -9226 7339 -9192
rect 7378 -9226 7411 -9192
rect 7446 -9226 7480 -9192
rect 7517 -9226 7548 -9192
rect 7589 -9226 7616 -9192
rect 7661 -9226 7684 -9192
rect 7733 -9226 7752 -9192
rect 7805 -9226 7820 -9192
rect 7877 -9226 7888 -9192
rect 7949 -9226 7956 -9192
rect 8021 -9226 8024 -9192
rect 8058 -9226 8059 -9192
rect 8126 -9226 8131 -9192
rect 8194 -9226 8203 -9192
rect 8262 -9226 8275 -9192
rect 8330 -9226 8347 -9192
rect 8398 -9226 8419 -9192
rect 8466 -9226 8491 -9192
rect 8534 -9226 8563 -9192
rect 8602 -9226 8635 -9192
rect 8670 -9226 8704 -9192
rect 8741 -9226 8772 -9192
rect 8813 -9226 8840 -9192
rect 8885 -9226 8908 -9192
rect 8957 -9226 8976 -9192
rect 9029 -9226 9044 -9192
rect 9101 -9226 9112 -9192
rect 9173 -9226 9180 -9192
rect 9245 -9226 9248 -9192
rect 9282 -9226 9283 -9192
rect 9350 -9226 9355 -9192
rect 9418 -9226 9427 -9192
rect 9486 -9226 9499 -9192
rect 9533 -9226 9647 -9192
rect 9681 -9226 9694 -9192
rect 9753 -9226 9762 -9192
rect 9825 -9226 9830 -9192
rect 9897 -9226 9898 -9192
rect 9932 -9226 9935 -9192
rect 10000 -9226 10007 -9192
rect 10068 -9226 10079 -9192
rect 10136 -9226 10151 -9192
rect 10204 -9226 10223 -9192
rect 10272 -9226 10295 -9192
rect 10340 -9226 10367 -9192
rect 10408 -9226 10439 -9192
rect 10476 -9226 10510 -9192
rect 10545 -9226 10578 -9192
rect 10617 -9226 10646 -9192
rect 10689 -9226 10714 -9192
rect 10761 -9226 10782 -9192
rect 10833 -9226 10850 -9192
rect 10905 -9226 10918 -9192
rect 10977 -9226 10986 -9192
rect 11049 -9226 11054 -9192
rect 11121 -9226 11122 -9192
rect 11156 -9226 11159 -9192
rect 11224 -9226 11231 -9192
rect 11292 -9226 11303 -9192
rect 11360 -9226 11375 -9192
rect 11428 -9226 11447 -9192
rect 11496 -9226 11519 -9192
rect 11564 -9226 11591 -9192
rect 11632 -9226 11663 -9192
rect 11700 -9226 11734 -9192
rect 11769 -9226 11802 -9192
rect 11841 -9226 11870 -9192
rect 11913 -9226 11938 -9192
rect 11985 -9226 12006 -9192
rect 12057 -9226 12074 -9192
rect 12129 -9226 12142 -9192
rect 12201 -9226 12210 -9192
rect 12273 -9226 12278 -9192
rect 12345 -9226 12346 -9192
rect 12380 -9226 12383 -9192
rect 12448 -9226 12455 -9192
rect 12516 -9226 12527 -9192
rect 12584 -9226 12599 -9192
rect 12652 -9226 12671 -9192
rect 12720 -9226 12743 -9192
rect 12788 -9226 12815 -9192
rect 12856 -9226 12887 -9192
rect 12924 -9226 12958 -9192
rect 12993 -9226 13026 -9192
rect 13065 -9226 13094 -9192
rect 13137 -9226 13162 -9192
rect 13209 -9226 13230 -9192
rect 13281 -9226 13298 -9192
rect 13353 -9226 13366 -9192
rect 13425 -9226 13434 -9192
rect 13497 -9226 13502 -9192
rect 13569 -9226 13570 -9192
rect 13604 -9226 13607 -9192
rect 13672 -9226 13679 -9192
rect 13740 -9226 13751 -9192
rect 13808 -9226 13823 -9192
rect 13857 -9226 14040 -9192
rect 14074 -9226 14089 -9192
rect 14146 -9226 14157 -9192
rect 14218 -9226 14225 -9192
rect 14290 -9226 14293 -9192
rect 14327 -9226 14328 -9192
rect 14395 -9226 14400 -9192
rect 14463 -9226 14472 -9192
rect 14531 -9226 14544 -9192
rect 14599 -9226 14616 -9192
rect 14667 -9226 14688 -9192
rect 14735 -9226 14760 -9192
rect 14803 -9226 14832 -9192
rect 14871 -9226 14904 -9192
rect 14939 -9226 14973 -9192
rect 15010 -9226 15041 -9192
rect 15082 -9226 15109 -9192
rect 15154 -9226 15177 -9192
rect 15226 -9226 15245 -9192
rect 15298 -9226 15313 -9192
rect 15370 -9226 15381 -9192
rect 15442 -9226 15449 -9192
rect 15514 -9226 15517 -9192
rect 15551 -9226 15552 -9192
rect 15619 -9226 15624 -9192
rect 15687 -9226 15696 -9192
rect 15755 -9226 15768 -9192
rect 15823 -9226 15840 -9192
rect 15891 -9226 15912 -9192
rect 15959 -9226 15984 -9192
rect 16027 -9226 16056 -9192
rect 16095 -9226 16128 -9192
rect 16163 -9226 16197 -9192
rect 16234 -9226 16265 -9192
rect 16306 -9226 16333 -9192
rect 16378 -9226 16401 -9192
rect 16450 -9226 16469 -9192
rect 16522 -9226 16537 -9192
rect 16594 -9226 16605 -9192
rect 16666 -9226 16673 -9192
rect 16738 -9226 16741 -9192
rect 16775 -9226 16776 -9192
rect 16843 -9226 16848 -9192
rect 16911 -9226 16920 -9192
rect 16979 -9226 16992 -9192
rect 17047 -9226 17064 -9192
rect 17115 -9226 17136 -9192
rect 17183 -9226 17208 -9192
rect 17251 -9226 17280 -9192
rect 17319 -9226 17352 -9192
rect 17387 -9226 17421 -9192
rect 17458 -9226 17489 -9192
rect 17530 -9226 17557 -9192
rect 17602 -9226 17625 -9192
rect 17674 -9226 17693 -9192
rect 17746 -9226 17761 -9192
rect 17818 -9226 17829 -9192
rect 17890 -9226 17897 -9192
rect 17962 -9226 17965 -9192
rect 17999 -9226 18000 -9192
rect 18067 -9226 18072 -9192
rect 18135 -9226 18144 -9192
rect 18203 -9226 18216 -9192
rect 18250 -9226 18324 -9192
<< viali >>
rect 930 429 964 463
rect 1002 429 1011 463
rect 1011 429 1036 463
rect 1074 429 1079 463
rect 1079 429 1108 463
rect 1146 429 1147 463
rect 1147 429 1180 463
rect 1218 429 1249 463
rect 1249 429 1252 463
rect 1290 429 1317 463
rect 1317 429 1324 463
rect 1362 429 1385 463
rect 1385 429 1396 463
rect 1434 429 1453 463
rect 1453 429 1468 463
rect 1506 429 1521 463
rect 1521 429 1540 463
rect 1578 429 1589 463
rect 1589 429 1612 463
rect 1650 429 1657 463
rect 1657 429 1684 463
rect 1722 429 1725 463
rect 1725 429 1756 463
rect 1794 429 1827 463
rect 1827 429 1828 463
rect 1866 429 1895 463
rect 1895 429 1900 463
rect 1938 429 1963 463
rect 1963 429 1972 463
rect 2010 429 2031 463
rect 2031 429 2044 463
rect 2082 429 2099 463
rect 2099 429 2116 463
rect 2154 429 2167 463
rect 2167 429 2188 463
rect 2226 429 2235 463
rect 2235 429 2260 463
rect 2298 429 2303 463
rect 2303 429 2332 463
rect 2370 429 2371 463
rect 2371 429 2404 463
rect 2442 429 2473 463
rect 2473 429 2476 463
rect 2514 429 2541 463
rect 2541 429 2548 463
rect 2586 429 2609 463
rect 2609 429 2620 463
rect 2658 429 2677 463
rect 2677 429 2692 463
rect 2730 429 2745 463
rect 2745 429 2764 463
rect 2802 429 2813 463
rect 2813 429 2836 463
rect 2874 429 2881 463
rect 2881 429 2908 463
rect 2946 429 2949 463
rect 2949 429 2980 463
rect 3018 429 3051 463
rect 3051 429 3052 463
rect 3090 429 3119 463
rect 3119 429 3124 463
rect 3162 429 3187 463
rect 3187 429 3196 463
rect 3234 429 3255 463
rect 3255 429 3268 463
rect 3306 429 3323 463
rect 3323 429 3340 463
rect 3378 429 3391 463
rect 3391 429 3412 463
rect 3450 429 3459 463
rect 3459 429 3484 463
rect 3522 429 3527 463
rect 3527 429 3556 463
rect 3594 429 3595 463
rect 3595 429 3628 463
rect 3666 429 3697 463
rect 3697 429 3700 463
rect 3738 429 3765 463
rect 3765 429 3772 463
rect 3810 429 3833 463
rect 3833 429 3844 463
rect 3882 429 3901 463
rect 3901 429 3916 463
rect 3954 429 3969 463
rect 3969 429 3988 463
rect 4026 429 4037 463
rect 4037 429 4060 463
rect 4098 429 4105 463
rect 4105 429 4132 463
rect 4170 429 4173 463
rect 4173 429 4204 463
rect 4242 429 4275 463
rect 4275 429 4276 463
rect 4314 429 4343 463
rect 4343 429 4348 463
rect 4386 429 4411 463
rect 4411 429 4420 463
rect 4458 429 4479 463
rect 4479 429 4492 463
rect 4530 429 4547 463
rect 4547 429 4564 463
rect 4602 429 4615 463
rect 4615 429 4636 463
rect 4674 429 4683 463
rect 4683 429 4708 463
rect 4746 429 4751 463
rect 4751 429 4780 463
rect 4818 429 4819 463
rect 4819 429 4852 463
rect 4890 429 4921 463
rect 4921 429 4924 463
rect 4962 429 4989 463
rect 4989 429 4996 463
rect 5034 429 5057 463
rect 5057 429 5068 463
rect 5106 429 5140 463
rect 5323 429 5357 463
rect 5395 429 5406 463
rect 5406 429 5429 463
rect 5467 429 5474 463
rect 5474 429 5501 463
rect 5539 429 5542 463
rect 5542 429 5573 463
rect 5611 429 5644 463
rect 5644 429 5645 463
rect 5683 429 5712 463
rect 5712 429 5717 463
rect 5755 429 5780 463
rect 5780 429 5789 463
rect 5827 429 5848 463
rect 5848 429 5861 463
rect 5899 429 5916 463
rect 5916 429 5933 463
rect 5971 429 5984 463
rect 5984 429 6005 463
rect 6043 429 6052 463
rect 6052 429 6077 463
rect 6115 429 6120 463
rect 6120 429 6149 463
rect 6187 429 6188 463
rect 6188 429 6221 463
rect 6259 429 6290 463
rect 6290 429 6293 463
rect 6331 429 6358 463
rect 6358 429 6365 463
rect 6403 429 6426 463
rect 6426 429 6437 463
rect 6475 429 6494 463
rect 6494 429 6509 463
rect 6547 429 6562 463
rect 6562 429 6581 463
rect 6619 429 6630 463
rect 6630 429 6653 463
rect 6691 429 6698 463
rect 6698 429 6725 463
rect 6763 429 6766 463
rect 6766 429 6797 463
rect 6835 429 6868 463
rect 6868 429 6869 463
rect 6907 429 6936 463
rect 6936 429 6941 463
rect 6979 429 7004 463
rect 7004 429 7013 463
rect 7051 429 7072 463
rect 7072 429 7085 463
rect 7123 429 7140 463
rect 7140 429 7157 463
rect 7195 429 7208 463
rect 7208 429 7229 463
rect 7267 429 7276 463
rect 7276 429 7301 463
rect 7339 429 7344 463
rect 7344 429 7373 463
rect 7411 429 7412 463
rect 7412 429 7445 463
rect 7483 429 7514 463
rect 7514 429 7517 463
rect 7555 429 7582 463
rect 7582 429 7589 463
rect 7627 429 7650 463
rect 7650 429 7661 463
rect 7699 429 7718 463
rect 7718 429 7733 463
rect 7771 429 7786 463
rect 7786 429 7805 463
rect 7843 429 7854 463
rect 7854 429 7877 463
rect 7915 429 7922 463
rect 7922 429 7949 463
rect 7987 429 7990 463
rect 7990 429 8021 463
rect 8059 429 8092 463
rect 8092 429 8093 463
rect 8131 429 8160 463
rect 8160 429 8165 463
rect 8203 429 8228 463
rect 8228 429 8237 463
rect 8275 429 8296 463
rect 8296 429 8309 463
rect 8347 429 8364 463
rect 8364 429 8381 463
rect 8419 429 8432 463
rect 8432 429 8453 463
rect 8491 429 8500 463
rect 8500 429 8525 463
rect 8563 429 8568 463
rect 8568 429 8597 463
rect 8635 429 8636 463
rect 8636 429 8669 463
rect 8707 429 8738 463
rect 8738 429 8741 463
rect 8779 429 8806 463
rect 8806 429 8813 463
rect 8851 429 8874 463
rect 8874 429 8885 463
rect 8923 429 8942 463
rect 8942 429 8957 463
rect 8995 429 9010 463
rect 9010 429 9029 463
rect 9067 429 9078 463
rect 9078 429 9101 463
rect 9139 429 9146 463
rect 9146 429 9173 463
rect 9211 429 9214 463
rect 9214 429 9245 463
rect 9283 429 9316 463
rect 9316 429 9317 463
rect 9355 429 9384 463
rect 9384 429 9389 463
rect 9427 429 9452 463
rect 9452 429 9461 463
rect 9499 429 9533 463
rect 9647 429 9681 463
rect 9719 429 9728 463
rect 9728 429 9753 463
rect 9791 429 9796 463
rect 9796 429 9825 463
rect 9863 429 9864 463
rect 9864 429 9897 463
rect 9935 429 9966 463
rect 9966 429 9969 463
rect 10007 429 10034 463
rect 10034 429 10041 463
rect 10079 429 10102 463
rect 10102 429 10113 463
rect 10151 429 10170 463
rect 10170 429 10185 463
rect 10223 429 10238 463
rect 10238 429 10257 463
rect 10295 429 10306 463
rect 10306 429 10329 463
rect 10367 429 10374 463
rect 10374 429 10401 463
rect 10439 429 10442 463
rect 10442 429 10473 463
rect 10511 429 10544 463
rect 10544 429 10545 463
rect 10583 429 10612 463
rect 10612 429 10617 463
rect 10655 429 10680 463
rect 10680 429 10689 463
rect 10727 429 10748 463
rect 10748 429 10761 463
rect 10799 429 10816 463
rect 10816 429 10833 463
rect 10871 429 10884 463
rect 10884 429 10905 463
rect 10943 429 10952 463
rect 10952 429 10977 463
rect 11015 429 11020 463
rect 11020 429 11049 463
rect 11087 429 11088 463
rect 11088 429 11121 463
rect 11159 429 11190 463
rect 11190 429 11193 463
rect 11231 429 11258 463
rect 11258 429 11265 463
rect 11303 429 11326 463
rect 11326 429 11337 463
rect 11375 429 11394 463
rect 11394 429 11409 463
rect 11447 429 11462 463
rect 11462 429 11481 463
rect 11519 429 11530 463
rect 11530 429 11553 463
rect 11591 429 11598 463
rect 11598 429 11625 463
rect 11663 429 11666 463
rect 11666 429 11697 463
rect 11735 429 11768 463
rect 11768 429 11769 463
rect 11807 429 11836 463
rect 11836 429 11841 463
rect 11879 429 11904 463
rect 11904 429 11913 463
rect 11951 429 11972 463
rect 11972 429 11985 463
rect 12023 429 12040 463
rect 12040 429 12057 463
rect 12095 429 12108 463
rect 12108 429 12129 463
rect 12167 429 12176 463
rect 12176 429 12201 463
rect 12239 429 12244 463
rect 12244 429 12273 463
rect 12311 429 12312 463
rect 12312 429 12345 463
rect 12383 429 12414 463
rect 12414 429 12417 463
rect 12455 429 12482 463
rect 12482 429 12489 463
rect 12527 429 12550 463
rect 12550 429 12561 463
rect 12599 429 12618 463
rect 12618 429 12633 463
rect 12671 429 12686 463
rect 12686 429 12705 463
rect 12743 429 12754 463
rect 12754 429 12777 463
rect 12815 429 12822 463
rect 12822 429 12849 463
rect 12887 429 12890 463
rect 12890 429 12921 463
rect 12959 429 12992 463
rect 12992 429 12993 463
rect 13031 429 13060 463
rect 13060 429 13065 463
rect 13103 429 13128 463
rect 13128 429 13137 463
rect 13175 429 13196 463
rect 13196 429 13209 463
rect 13247 429 13264 463
rect 13264 429 13281 463
rect 13319 429 13332 463
rect 13332 429 13353 463
rect 13391 429 13400 463
rect 13400 429 13425 463
rect 13463 429 13468 463
rect 13468 429 13497 463
rect 13535 429 13536 463
rect 13536 429 13569 463
rect 13607 429 13638 463
rect 13638 429 13641 463
rect 13679 429 13706 463
rect 13706 429 13713 463
rect 13751 429 13774 463
rect 13774 429 13785 463
rect 13823 429 13857 463
rect 14040 429 14074 463
rect 14112 429 14123 463
rect 14123 429 14146 463
rect 14184 429 14191 463
rect 14191 429 14218 463
rect 14256 429 14259 463
rect 14259 429 14290 463
rect 14328 429 14361 463
rect 14361 429 14362 463
rect 14400 429 14429 463
rect 14429 429 14434 463
rect 14472 429 14497 463
rect 14497 429 14506 463
rect 14544 429 14565 463
rect 14565 429 14578 463
rect 14616 429 14633 463
rect 14633 429 14650 463
rect 14688 429 14701 463
rect 14701 429 14722 463
rect 14760 429 14769 463
rect 14769 429 14794 463
rect 14832 429 14837 463
rect 14837 429 14866 463
rect 14904 429 14905 463
rect 14905 429 14938 463
rect 14976 429 15007 463
rect 15007 429 15010 463
rect 15048 429 15075 463
rect 15075 429 15082 463
rect 15120 429 15143 463
rect 15143 429 15154 463
rect 15192 429 15211 463
rect 15211 429 15226 463
rect 15264 429 15279 463
rect 15279 429 15298 463
rect 15336 429 15347 463
rect 15347 429 15370 463
rect 15408 429 15415 463
rect 15415 429 15442 463
rect 15480 429 15483 463
rect 15483 429 15514 463
rect 15552 429 15585 463
rect 15585 429 15586 463
rect 15624 429 15653 463
rect 15653 429 15658 463
rect 15696 429 15721 463
rect 15721 429 15730 463
rect 15768 429 15789 463
rect 15789 429 15802 463
rect 15840 429 15857 463
rect 15857 429 15874 463
rect 15912 429 15925 463
rect 15925 429 15946 463
rect 15984 429 15993 463
rect 15993 429 16018 463
rect 16056 429 16061 463
rect 16061 429 16090 463
rect 16128 429 16129 463
rect 16129 429 16162 463
rect 16200 429 16231 463
rect 16231 429 16234 463
rect 16272 429 16299 463
rect 16299 429 16306 463
rect 16344 429 16367 463
rect 16367 429 16378 463
rect 16416 429 16435 463
rect 16435 429 16450 463
rect 16488 429 16503 463
rect 16503 429 16522 463
rect 16560 429 16571 463
rect 16571 429 16594 463
rect 16632 429 16639 463
rect 16639 429 16666 463
rect 16704 429 16707 463
rect 16707 429 16738 463
rect 16776 429 16809 463
rect 16809 429 16810 463
rect 16848 429 16877 463
rect 16877 429 16882 463
rect 16920 429 16945 463
rect 16945 429 16954 463
rect 16992 429 17013 463
rect 17013 429 17026 463
rect 17064 429 17081 463
rect 17081 429 17098 463
rect 17136 429 17149 463
rect 17149 429 17170 463
rect 17208 429 17217 463
rect 17217 429 17242 463
rect 17280 429 17285 463
rect 17285 429 17314 463
rect 17352 429 17353 463
rect 17353 429 17386 463
rect 17424 429 17455 463
rect 17455 429 17458 463
rect 17496 429 17523 463
rect 17523 429 17530 463
rect 17568 429 17591 463
rect 17591 429 17602 463
rect 17640 429 17659 463
rect 17659 429 17674 463
rect 17712 429 17727 463
rect 17727 429 17746 463
rect 17784 429 17795 463
rect 17795 429 17818 463
rect 17856 429 17863 463
rect 17863 429 17890 463
rect 17928 429 17931 463
rect 17931 429 17962 463
rect 18000 429 18033 463
rect 18033 429 18034 463
rect 18072 429 18101 463
rect 18101 429 18106 463
rect 18144 429 18169 463
rect 18169 429 18178 463
rect 18216 429 18250 463
rect 1064 315 1066 349
rect 1066 315 1098 349
rect 1136 315 1168 349
rect 1168 315 1170 349
rect 1516 315 1518 349
rect 1518 315 1550 349
rect 1588 315 1620 349
rect 1620 315 1622 349
rect 1774 315 1776 349
rect 1776 315 1808 349
rect 1846 315 1878 349
rect 1878 315 1880 349
rect 2032 315 2034 349
rect 2034 315 2066 349
rect 2104 315 2136 349
rect 2136 315 2138 349
rect 2290 315 2292 349
rect 2292 315 2324 349
rect 2362 315 2394 349
rect 2394 315 2396 349
rect 2742 315 2744 349
rect 2744 315 2776 349
rect 2814 315 2846 349
rect 2846 315 2848 349
rect 3000 315 3002 349
rect 3002 315 3034 349
rect 3072 315 3104 349
rect 3104 315 3106 349
rect 3258 315 3260 349
rect 3260 315 3292 349
rect 3330 315 3362 349
rect 3362 315 3364 349
rect 3710 315 3712 349
rect 3712 315 3744 349
rect 3782 315 3814 349
rect 3814 315 3816 349
rect 3968 315 3970 349
rect 3970 315 4002 349
rect 4040 315 4072 349
rect 4072 315 4074 349
rect 4226 315 4228 349
rect 4228 315 4260 349
rect 4298 315 4330 349
rect 4330 315 4332 349
rect 4484 315 4486 349
rect 4486 315 4518 349
rect 4556 315 4588 349
rect 4588 315 4590 349
rect 4935 315 4937 349
rect 4937 315 4969 349
rect 5007 315 5039 349
rect 5039 315 5041 349
rect 856 272 890 306
rect 5421 315 5423 349
rect 5423 315 5455 349
rect 5493 315 5525 349
rect 5525 315 5527 349
rect 5873 315 5875 349
rect 5875 315 5907 349
rect 5945 315 5977 349
rect 5977 315 5979 349
rect 6131 315 6133 349
rect 6133 315 6165 349
rect 6203 315 6235 349
rect 6235 315 6237 349
rect 6389 315 6391 349
rect 6391 315 6423 349
rect 6461 315 6493 349
rect 6493 315 6495 349
rect 6647 315 6649 349
rect 6649 315 6681 349
rect 6719 315 6751 349
rect 6751 315 6753 349
rect 7099 315 7101 349
rect 7101 315 7133 349
rect 7171 315 7203 349
rect 7203 315 7205 349
rect 7357 315 7359 349
rect 7359 315 7391 349
rect 7429 315 7461 349
rect 7461 315 7463 349
rect 7615 315 7617 349
rect 7617 315 7649 349
rect 7687 315 7719 349
rect 7719 315 7721 349
rect 8067 315 8069 349
rect 8069 315 8101 349
rect 8139 315 8171 349
rect 8171 315 8173 349
rect 8325 315 8327 349
rect 8327 315 8359 349
rect 8397 315 8429 349
rect 8429 315 8431 349
rect 8583 315 8585 349
rect 8585 315 8617 349
rect 8655 315 8687 349
rect 8687 315 8689 349
rect 8841 315 8843 349
rect 8843 315 8875 349
rect 8913 315 8945 349
rect 8945 315 8947 349
rect 9293 315 9295 349
rect 9295 315 9327 349
rect 9365 315 9397 349
rect 9397 315 9399 349
rect 5214 272 5248 306
rect 9781 315 9783 349
rect 9783 315 9815 349
rect 9853 315 9885 349
rect 9885 315 9887 349
rect 10233 315 10235 349
rect 10235 315 10267 349
rect 10305 315 10337 349
rect 10337 315 10339 349
rect 10491 315 10493 349
rect 10493 315 10525 349
rect 10563 315 10595 349
rect 10595 315 10597 349
rect 10749 315 10751 349
rect 10751 315 10783 349
rect 10821 315 10853 349
rect 10853 315 10855 349
rect 11007 315 11009 349
rect 11009 315 11041 349
rect 11079 315 11111 349
rect 11111 315 11113 349
rect 11459 315 11461 349
rect 11461 315 11493 349
rect 11531 315 11563 349
rect 11563 315 11565 349
rect 11717 315 11719 349
rect 11719 315 11751 349
rect 11789 315 11821 349
rect 11821 315 11823 349
rect 11975 315 11977 349
rect 11977 315 12009 349
rect 12047 315 12079 349
rect 12079 315 12081 349
rect 12427 315 12429 349
rect 12429 315 12461 349
rect 12499 315 12531 349
rect 12531 315 12533 349
rect 12685 315 12687 349
rect 12687 315 12719 349
rect 12757 315 12789 349
rect 12789 315 12791 349
rect 12943 315 12945 349
rect 12945 315 12977 349
rect 13015 315 13047 349
rect 13047 315 13049 349
rect 13201 315 13203 349
rect 13203 315 13235 349
rect 13273 315 13305 349
rect 13305 315 13307 349
rect 13653 315 13655 349
rect 13655 315 13687 349
rect 13725 315 13757 349
rect 13757 315 13759 349
rect 9573 272 9607 306
rect 14139 315 14141 349
rect 14141 315 14173 349
rect 14211 315 14243 349
rect 14243 315 14245 349
rect 14590 315 14592 349
rect 14592 315 14624 349
rect 14662 315 14694 349
rect 14694 315 14696 349
rect 14848 315 14850 349
rect 14850 315 14882 349
rect 14920 315 14952 349
rect 14952 315 14954 349
rect 15106 315 15108 349
rect 15108 315 15140 349
rect 15178 315 15210 349
rect 15210 315 15212 349
rect 15364 315 15366 349
rect 15366 315 15398 349
rect 15436 315 15468 349
rect 15468 315 15470 349
rect 15816 315 15818 349
rect 15818 315 15850 349
rect 15888 315 15920 349
rect 15920 315 15922 349
rect 16074 315 16076 349
rect 16076 315 16108 349
rect 16146 315 16178 349
rect 16178 315 16180 349
rect 16332 315 16334 349
rect 16334 315 16366 349
rect 16404 315 16436 349
rect 16436 315 16438 349
rect 16784 315 16786 349
rect 16786 315 16818 349
rect 16856 315 16888 349
rect 16888 315 16890 349
rect 17042 315 17044 349
rect 17044 315 17076 349
rect 17114 315 17146 349
rect 17146 315 17148 349
rect 17300 315 17302 349
rect 17302 315 17334 349
rect 17372 315 17404 349
rect 17404 315 17406 349
rect 17558 315 17560 349
rect 17560 315 17592 349
rect 17630 315 17662 349
rect 17662 315 17664 349
rect 18010 315 18012 349
rect 18012 315 18044 349
rect 18082 315 18114 349
rect 18114 315 18116 349
rect 13932 272 13966 306
rect 18290 272 18324 306
rect 856 216 890 234
rect 856 200 890 216
rect 856 148 890 162
rect 856 128 890 148
rect 856 80 890 90
rect 856 56 890 80
rect 971 219 1005 221
rect 971 187 1005 219
rect 971 117 1005 149
rect 971 115 1005 117
rect 1229 219 1263 221
rect 1229 187 1263 219
rect 1229 117 1263 149
rect 1229 115 1263 117
rect 1423 219 1457 221
rect 1423 187 1457 219
rect 1423 117 1457 149
rect 1423 115 1457 117
rect 1681 219 1715 221
rect 1681 187 1715 219
rect 1681 117 1715 149
rect 1681 115 1715 117
rect 1939 219 1973 221
rect 1939 187 1973 219
rect 1939 117 1973 149
rect 1939 115 1973 117
rect 2197 219 2231 221
rect 2197 187 2231 219
rect 2197 117 2231 149
rect 2197 115 2231 117
rect 2455 219 2489 221
rect 2455 187 2489 219
rect 2455 117 2489 149
rect 2455 115 2489 117
rect 2649 219 2683 221
rect 2649 187 2683 219
rect 2649 117 2683 149
rect 2649 115 2683 117
rect 2907 219 2941 221
rect 2907 187 2941 219
rect 2907 117 2941 149
rect 2907 115 2941 117
rect 3165 219 3199 221
rect 3165 187 3199 219
rect 3165 117 3199 149
rect 3165 115 3199 117
rect 3423 219 3457 221
rect 3423 187 3457 219
rect 3423 117 3457 149
rect 3423 115 3457 117
rect 3617 219 3651 221
rect 3617 187 3651 219
rect 3617 117 3651 149
rect 3617 115 3651 117
rect 3875 219 3909 221
rect 3875 187 3909 219
rect 3875 117 3909 149
rect 3875 115 3909 117
rect 4133 219 4167 221
rect 4133 187 4167 219
rect 4133 117 4167 149
rect 4133 115 4167 117
rect 4391 219 4425 221
rect 4391 187 4425 219
rect 4391 117 4425 149
rect 4391 115 4425 117
rect 4649 219 4683 221
rect 4649 187 4683 219
rect 4649 117 4683 149
rect 4649 115 4683 117
rect 4842 219 4876 221
rect 4842 187 4876 219
rect 4842 117 4876 149
rect 4842 115 4876 117
rect 5100 219 5134 221
rect 5100 187 5134 219
rect 5100 117 5134 149
rect 5100 115 5134 117
rect 5214 216 5248 234
rect 5214 200 5248 216
rect 5214 148 5248 162
rect 5214 128 5248 148
rect 5214 80 5248 90
rect 856 12 890 18
rect 856 -16 890 12
rect 856 -56 890 -54
rect 856 -88 890 -56
rect 856 -158 890 -126
rect 856 -160 890 -158
rect 856 -226 890 -198
rect 856 -232 890 -226
rect 856 -294 890 -270
rect 856 -304 890 -294
rect 5214 56 5248 80
rect 5328 219 5362 221
rect 5328 187 5362 219
rect 5328 117 5362 149
rect 5328 115 5362 117
rect 5586 219 5620 221
rect 5586 187 5620 219
rect 5586 117 5620 149
rect 5586 115 5620 117
rect 5780 219 5814 221
rect 5780 187 5814 219
rect 5780 117 5814 149
rect 5780 115 5814 117
rect 6038 219 6072 221
rect 6038 187 6072 219
rect 6038 117 6072 149
rect 6038 115 6072 117
rect 6296 219 6330 221
rect 6296 187 6330 219
rect 6296 117 6330 149
rect 6296 115 6330 117
rect 6554 219 6588 221
rect 6554 187 6588 219
rect 6554 117 6588 149
rect 6554 115 6588 117
rect 6812 219 6846 221
rect 6812 187 6846 219
rect 6812 117 6846 149
rect 6812 115 6846 117
rect 7006 219 7040 221
rect 7006 187 7040 219
rect 7006 117 7040 149
rect 7006 115 7040 117
rect 7264 219 7298 221
rect 7264 187 7298 219
rect 7264 117 7298 149
rect 7264 115 7298 117
rect 7522 219 7556 221
rect 7522 187 7556 219
rect 7522 117 7556 149
rect 7522 115 7556 117
rect 7780 219 7814 221
rect 7780 187 7814 219
rect 7780 117 7814 149
rect 7780 115 7814 117
rect 7974 219 8008 221
rect 7974 187 8008 219
rect 7974 117 8008 149
rect 7974 115 8008 117
rect 8232 219 8266 221
rect 8232 187 8266 219
rect 8232 117 8266 149
rect 8232 115 8266 117
rect 8490 219 8524 221
rect 8490 187 8524 219
rect 8490 117 8524 149
rect 8490 115 8524 117
rect 8748 219 8782 221
rect 8748 187 8782 219
rect 8748 117 8782 149
rect 8748 115 8782 117
rect 9006 219 9040 221
rect 9006 187 9040 219
rect 9006 117 9040 149
rect 9006 115 9040 117
rect 9200 219 9234 221
rect 9200 187 9234 219
rect 9200 117 9234 149
rect 9200 115 9234 117
rect 9458 219 9492 221
rect 9458 187 9492 219
rect 9458 117 9492 149
rect 9458 115 9492 117
rect 9573 216 9607 234
rect 9573 200 9607 216
rect 9573 148 9607 162
rect 9573 128 9607 148
rect 9573 80 9607 90
rect 5214 12 5248 18
rect 5214 -16 5248 12
rect 5214 -56 5248 -54
rect 5214 -88 5248 -56
rect 5214 -158 5248 -126
rect 5214 -160 5248 -158
rect 5214 -226 5248 -198
rect 5214 -232 5248 -226
rect 5214 -294 5248 -270
rect 5214 -304 5248 -294
rect 9573 56 9607 80
rect 9688 219 9722 221
rect 9688 187 9722 219
rect 9688 117 9722 149
rect 9688 115 9722 117
rect 9946 219 9980 221
rect 9946 187 9980 219
rect 9946 117 9980 149
rect 9946 115 9980 117
rect 10140 219 10174 221
rect 10140 187 10174 219
rect 10140 117 10174 149
rect 10140 115 10174 117
rect 10398 219 10432 221
rect 10398 187 10432 219
rect 10398 117 10432 149
rect 10398 115 10432 117
rect 10656 219 10690 221
rect 10656 187 10690 219
rect 10656 117 10690 149
rect 10656 115 10690 117
rect 10914 219 10948 221
rect 10914 187 10948 219
rect 10914 117 10948 149
rect 10914 115 10948 117
rect 11172 219 11206 221
rect 11172 187 11206 219
rect 11172 117 11206 149
rect 11172 115 11206 117
rect 11366 219 11400 221
rect 11366 187 11400 219
rect 11366 117 11400 149
rect 11366 115 11400 117
rect 11624 219 11658 221
rect 11624 187 11658 219
rect 11624 117 11658 149
rect 11624 115 11658 117
rect 11882 219 11916 221
rect 11882 187 11916 219
rect 11882 117 11916 149
rect 11882 115 11916 117
rect 12140 219 12174 221
rect 12140 187 12174 219
rect 12140 117 12174 149
rect 12140 115 12174 117
rect 12334 219 12368 221
rect 12334 187 12368 219
rect 12334 117 12368 149
rect 12334 115 12368 117
rect 12592 219 12626 221
rect 12592 187 12626 219
rect 12592 117 12626 149
rect 12592 115 12626 117
rect 12850 219 12884 221
rect 12850 187 12884 219
rect 12850 117 12884 149
rect 12850 115 12884 117
rect 13108 219 13142 221
rect 13108 187 13142 219
rect 13108 117 13142 149
rect 13108 115 13142 117
rect 13366 219 13400 221
rect 13366 187 13400 219
rect 13366 117 13400 149
rect 13366 115 13400 117
rect 13560 219 13594 221
rect 13560 187 13594 219
rect 13560 117 13594 149
rect 13560 115 13594 117
rect 13818 219 13852 221
rect 13818 187 13852 219
rect 13818 117 13852 149
rect 13818 115 13852 117
rect 13932 216 13966 234
rect 13932 200 13966 216
rect 13932 148 13966 162
rect 13932 128 13966 148
rect 9573 12 9607 18
rect 9573 -16 9607 12
rect 9573 -56 9607 -54
rect 9573 -88 9607 -56
rect 9573 -158 9607 -126
rect 9573 -160 9607 -158
rect 9573 -226 9607 -198
rect 9573 -232 9607 -226
rect 9573 -294 9607 -270
rect 9573 -304 9607 -294
rect 13932 80 13966 90
rect 13932 56 13966 80
rect 14046 219 14080 221
rect 14046 187 14080 219
rect 14046 117 14080 149
rect 14046 115 14080 117
rect 14304 219 14338 221
rect 14304 187 14338 219
rect 14304 117 14338 149
rect 14304 115 14338 117
rect 14497 219 14531 221
rect 14497 187 14531 219
rect 14497 117 14531 149
rect 14497 115 14531 117
rect 14755 219 14789 221
rect 14755 187 14789 219
rect 14755 117 14789 149
rect 14755 115 14789 117
rect 15013 219 15047 221
rect 15013 187 15047 219
rect 15013 117 15047 149
rect 15013 115 15047 117
rect 15271 219 15305 221
rect 15271 187 15305 219
rect 15271 117 15305 149
rect 15271 115 15305 117
rect 15529 219 15563 221
rect 15529 187 15563 219
rect 15529 117 15563 149
rect 15529 115 15563 117
rect 15723 219 15757 221
rect 15723 187 15757 219
rect 15723 117 15757 149
rect 15723 115 15757 117
rect 15981 219 16015 221
rect 15981 187 16015 219
rect 15981 117 16015 149
rect 15981 115 16015 117
rect 16239 219 16273 221
rect 16239 187 16273 219
rect 16239 117 16273 149
rect 16239 115 16273 117
rect 16497 219 16531 221
rect 16497 187 16531 219
rect 16497 117 16531 149
rect 16497 115 16531 117
rect 16691 219 16725 221
rect 16691 187 16725 219
rect 16691 117 16725 149
rect 16691 115 16725 117
rect 16949 219 16983 221
rect 16949 187 16983 219
rect 16949 117 16983 149
rect 16949 115 16983 117
rect 17207 219 17241 221
rect 17207 187 17241 219
rect 17207 117 17241 149
rect 17207 115 17241 117
rect 17465 219 17499 221
rect 17465 187 17499 219
rect 17465 117 17499 149
rect 17465 115 17499 117
rect 17723 219 17757 221
rect 17723 187 17757 219
rect 17723 117 17757 149
rect 17723 115 17757 117
rect 17917 219 17951 221
rect 17917 187 17951 219
rect 17917 117 17951 149
rect 17917 115 17951 117
rect 18175 219 18209 221
rect 18175 187 18209 219
rect 18175 117 18209 149
rect 18175 115 18209 117
rect 18290 216 18324 234
rect 18290 200 18324 216
rect 18290 148 18324 162
rect 18290 128 18324 148
rect 18290 80 18324 90
rect 13932 12 13966 18
rect 13932 -16 13966 12
rect 13932 -56 13966 -54
rect 13932 -88 13966 -56
rect 13932 -158 13966 -126
rect 13932 -160 13966 -158
rect 13932 -226 13966 -198
rect 13932 -232 13966 -226
rect 13932 -294 13966 -270
rect 13932 -304 13966 -294
rect 18290 56 18324 80
rect 18290 12 18324 18
rect 18290 -16 18324 12
rect 18290 -56 18324 -54
rect 18290 -88 18324 -56
rect 18290 -158 18324 -126
rect 18290 -160 18324 -158
rect 18290 -226 18324 -198
rect 18290 -232 18324 -226
rect 18290 -294 18324 -270
rect 18290 -304 18324 -294
rect 856 -362 890 -342
rect 5214 -362 5248 -342
rect 9573 -362 9607 -342
rect 13932 -362 13966 -342
rect 18290 -362 18324 -342
rect 856 -376 890 -362
rect 856 -430 890 -414
rect 856 -448 890 -430
rect 856 -498 890 -486
rect 856 -520 890 -498
rect 856 -566 890 -558
rect 856 -592 890 -566
rect 856 -634 890 -630
rect 856 -664 890 -634
rect 5214 -376 5248 -362
rect 5214 -430 5248 -414
rect 5214 -448 5248 -430
rect 5214 -498 5248 -486
rect 5214 -520 5248 -498
rect 5214 -566 5248 -558
rect 5214 -592 5248 -566
rect 5214 -634 5248 -630
rect 5214 -664 5248 -634
rect 856 -736 890 -702
rect 856 -804 890 -774
rect 856 -808 890 -804
rect 856 -872 890 -846
rect 856 -880 890 -872
rect 971 -725 1005 -723
rect 971 -757 1005 -725
rect 971 -827 1005 -795
rect 971 -829 1005 -827
rect 1229 -725 1263 -723
rect 1229 -757 1263 -725
rect 1229 -827 1263 -795
rect 1229 -829 1263 -827
rect 1423 -725 1457 -723
rect 1423 -757 1457 -725
rect 1423 -827 1457 -795
rect 1423 -829 1457 -827
rect 1681 -725 1715 -723
rect 1681 -757 1715 -725
rect 1681 -827 1715 -795
rect 1681 -829 1715 -827
rect 1939 -725 1973 -723
rect 1939 -757 1973 -725
rect 1939 -827 1973 -795
rect 1939 -829 1973 -827
rect 2197 -725 2231 -723
rect 2197 -757 2231 -725
rect 2197 -827 2231 -795
rect 2197 -829 2231 -827
rect 2455 -725 2489 -723
rect 2455 -757 2489 -725
rect 2455 -827 2489 -795
rect 2455 -829 2489 -827
rect 2649 -725 2683 -723
rect 2649 -757 2683 -725
rect 2649 -827 2683 -795
rect 2649 -829 2683 -827
rect 2907 -725 2941 -723
rect 2907 -757 2941 -725
rect 2907 -827 2941 -795
rect 2907 -829 2941 -827
rect 3165 -725 3199 -723
rect 3165 -757 3199 -725
rect 3165 -827 3199 -795
rect 3165 -829 3199 -827
rect 3423 -725 3457 -723
rect 3423 -757 3457 -725
rect 3423 -827 3457 -795
rect 3423 -829 3457 -827
rect 3617 -725 3651 -723
rect 3617 -757 3651 -725
rect 3617 -827 3651 -795
rect 3617 -829 3651 -827
rect 3875 -725 3909 -723
rect 3875 -757 3909 -725
rect 3875 -827 3909 -795
rect 3875 -829 3909 -827
rect 4133 -725 4167 -723
rect 4133 -757 4167 -725
rect 4133 -827 4167 -795
rect 4133 -829 4167 -827
rect 4391 -725 4425 -723
rect 4391 -757 4425 -725
rect 4391 -827 4425 -795
rect 4391 -829 4425 -827
rect 4649 -725 4683 -723
rect 4649 -757 4683 -725
rect 4649 -827 4683 -795
rect 4649 -829 4683 -827
rect 4842 -725 4876 -723
rect 4842 -757 4876 -725
rect 4842 -827 4876 -795
rect 4842 -829 4876 -827
rect 5100 -725 5134 -723
rect 5100 -757 5134 -725
rect 5100 -827 5134 -795
rect 5100 -829 5134 -827
rect 9573 -376 9607 -362
rect 9573 -430 9607 -414
rect 9573 -448 9607 -430
rect 9573 -498 9607 -486
rect 9573 -520 9607 -498
rect 9573 -566 9607 -558
rect 9573 -592 9607 -566
rect 9573 -634 9607 -630
rect 9573 -664 9607 -634
rect 5214 -736 5248 -702
rect 5214 -804 5248 -774
rect 5214 -808 5248 -804
rect 5214 -872 5248 -846
rect 5214 -880 5248 -872
rect 5328 -725 5362 -723
rect 5328 -757 5362 -725
rect 5328 -827 5362 -795
rect 5328 -829 5362 -827
rect 5586 -725 5620 -723
rect 5586 -757 5620 -725
rect 5586 -827 5620 -795
rect 5586 -829 5620 -827
rect 5780 -725 5814 -723
rect 5780 -757 5814 -725
rect 5780 -827 5814 -795
rect 5780 -829 5814 -827
rect 6038 -725 6072 -723
rect 6038 -757 6072 -725
rect 6038 -827 6072 -795
rect 6038 -829 6072 -827
rect 6296 -725 6330 -723
rect 6296 -757 6330 -725
rect 6296 -827 6330 -795
rect 6296 -829 6330 -827
rect 6554 -725 6588 -723
rect 6554 -757 6588 -725
rect 6554 -827 6588 -795
rect 6554 -829 6588 -827
rect 6812 -725 6846 -723
rect 6812 -757 6846 -725
rect 6812 -827 6846 -795
rect 6812 -829 6846 -827
rect 7006 -725 7040 -723
rect 7006 -757 7040 -725
rect 7006 -827 7040 -795
rect 7006 -829 7040 -827
rect 7264 -725 7298 -723
rect 7264 -757 7298 -725
rect 7264 -827 7298 -795
rect 7264 -829 7298 -827
rect 7522 -725 7556 -723
rect 7522 -757 7556 -725
rect 7522 -827 7556 -795
rect 7522 -829 7556 -827
rect 7780 -725 7814 -723
rect 7780 -757 7814 -725
rect 7780 -827 7814 -795
rect 7780 -829 7814 -827
rect 7974 -725 8008 -723
rect 7974 -757 8008 -725
rect 7974 -827 8008 -795
rect 7974 -829 8008 -827
rect 8232 -725 8266 -723
rect 8232 -757 8266 -725
rect 8232 -827 8266 -795
rect 8232 -829 8266 -827
rect 8490 -725 8524 -723
rect 8490 -757 8524 -725
rect 8490 -827 8524 -795
rect 8490 -829 8524 -827
rect 8748 -725 8782 -723
rect 8748 -757 8782 -725
rect 8748 -827 8782 -795
rect 8748 -829 8782 -827
rect 9006 -725 9040 -723
rect 9006 -757 9040 -725
rect 9006 -827 9040 -795
rect 9006 -829 9040 -827
rect 9200 -725 9234 -723
rect 9200 -757 9234 -725
rect 9200 -827 9234 -795
rect 9200 -829 9234 -827
rect 9458 -725 9492 -723
rect 9458 -757 9492 -725
rect 9458 -827 9492 -795
rect 9458 -829 9492 -827
rect 13932 -376 13966 -362
rect 13932 -430 13966 -414
rect 13932 -448 13966 -430
rect 13932 -498 13966 -486
rect 13932 -520 13966 -498
rect 13932 -566 13966 -558
rect 13932 -592 13966 -566
rect 13932 -634 13966 -630
rect 13932 -664 13966 -634
rect 9573 -736 9607 -702
rect 9573 -804 9607 -774
rect 9573 -808 9607 -804
rect 9573 -872 9607 -846
rect 9573 -880 9607 -872
rect 9688 -725 9722 -723
rect 9688 -757 9722 -725
rect 9688 -827 9722 -795
rect 9688 -829 9722 -827
rect 9946 -725 9980 -723
rect 9946 -757 9980 -725
rect 9946 -827 9980 -795
rect 9946 -829 9980 -827
rect 10140 -725 10174 -723
rect 10140 -757 10174 -725
rect 10140 -827 10174 -795
rect 10140 -829 10174 -827
rect 10398 -725 10432 -723
rect 10398 -757 10432 -725
rect 10398 -827 10432 -795
rect 10398 -829 10432 -827
rect 10656 -725 10690 -723
rect 10656 -757 10690 -725
rect 10656 -827 10690 -795
rect 10656 -829 10690 -827
rect 10914 -725 10948 -723
rect 10914 -757 10948 -725
rect 10914 -827 10948 -795
rect 10914 -829 10948 -827
rect 11172 -725 11206 -723
rect 11172 -757 11206 -725
rect 11172 -827 11206 -795
rect 11172 -829 11206 -827
rect 11366 -725 11400 -723
rect 11366 -757 11400 -725
rect 11366 -827 11400 -795
rect 11366 -829 11400 -827
rect 11624 -725 11658 -723
rect 11624 -757 11658 -725
rect 11624 -827 11658 -795
rect 11624 -829 11658 -827
rect 11882 -725 11916 -723
rect 11882 -757 11916 -725
rect 11882 -827 11916 -795
rect 11882 -829 11916 -827
rect 12140 -725 12174 -723
rect 12140 -757 12174 -725
rect 12140 -827 12174 -795
rect 12140 -829 12174 -827
rect 12334 -725 12368 -723
rect 12334 -757 12368 -725
rect 12334 -827 12368 -795
rect 12334 -829 12368 -827
rect 12592 -725 12626 -723
rect 12592 -757 12626 -725
rect 12592 -827 12626 -795
rect 12592 -829 12626 -827
rect 12850 -725 12884 -723
rect 12850 -757 12884 -725
rect 12850 -827 12884 -795
rect 12850 -829 12884 -827
rect 13108 -725 13142 -723
rect 13108 -757 13142 -725
rect 13108 -827 13142 -795
rect 13108 -829 13142 -827
rect 13366 -725 13400 -723
rect 13366 -757 13400 -725
rect 13366 -827 13400 -795
rect 13366 -829 13400 -827
rect 13560 -725 13594 -723
rect 13560 -757 13594 -725
rect 13560 -827 13594 -795
rect 13560 -829 13594 -827
rect 13818 -725 13852 -723
rect 13818 -757 13852 -725
rect 13818 -827 13852 -795
rect 13818 -829 13852 -827
rect 18290 -376 18324 -362
rect 18290 -430 18324 -414
rect 18290 -448 18324 -430
rect 18290 -498 18324 -486
rect 18290 -520 18324 -498
rect 18290 -566 18324 -558
rect 18290 -592 18324 -566
rect 18290 -634 18324 -630
rect 18290 -664 18324 -634
rect 13932 -736 13966 -702
rect 13932 -804 13966 -774
rect 13932 -808 13966 -804
rect 13932 -872 13966 -846
rect 13932 -880 13966 -872
rect 14046 -725 14080 -723
rect 14046 -757 14080 -725
rect 14046 -827 14080 -795
rect 14046 -829 14080 -827
rect 14304 -725 14338 -723
rect 14304 -757 14338 -725
rect 14304 -827 14338 -795
rect 14304 -829 14338 -827
rect 14497 -725 14531 -723
rect 14497 -757 14531 -725
rect 14497 -827 14531 -795
rect 14497 -829 14531 -827
rect 14755 -725 14789 -723
rect 14755 -757 14789 -725
rect 14755 -827 14789 -795
rect 14755 -829 14789 -827
rect 15013 -725 15047 -723
rect 15013 -757 15047 -725
rect 15013 -827 15047 -795
rect 15013 -829 15047 -827
rect 15271 -725 15305 -723
rect 15271 -757 15305 -725
rect 15271 -827 15305 -795
rect 15271 -829 15305 -827
rect 15529 -725 15563 -723
rect 15529 -757 15563 -725
rect 15529 -827 15563 -795
rect 15529 -829 15563 -827
rect 15723 -725 15757 -723
rect 15723 -757 15757 -725
rect 15723 -827 15757 -795
rect 15723 -829 15757 -827
rect 15981 -725 16015 -723
rect 15981 -757 16015 -725
rect 15981 -827 16015 -795
rect 15981 -829 16015 -827
rect 16239 -725 16273 -723
rect 16239 -757 16273 -725
rect 16239 -827 16273 -795
rect 16239 -829 16273 -827
rect 16497 -725 16531 -723
rect 16497 -757 16531 -725
rect 16497 -827 16531 -795
rect 16497 -829 16531 -827
rect 16691 -725 16725 -723
rect 16691 -757 16725 -725
rect 16691 -827 16725 -795
rect 16691 -829 16725 -827
rect 16949 -725 16983 -723
rect 16949 -757 16983 -725
rect 16949 -827 16983 -795
rect 16949 -829 16983 -827
rect 17207 -725 17241 -723
rect 17207 -757 17241 -725
rect 17207 -827 17241 -795
rect 17207 -829 17241 -827
rect 17465 -725 17499 -723
rect 17465 -757 17499 -725
rect 17465 -827 17499 -795
rect 17465 -829 17499 -827
rect 17723 -725 17757 -723
rect 17723 -757 17757 -725
rect 17723 -827 17757 -795
rect 17723 -829 17757 -827
rect 17917 -725 17951 -723
rect 17917 -757 17951 -725
rect 17917 -827 17951 -795
rect 17917 -829 17951 -827
rect 18175 -725 18209 -723
rect 18175 -757 18209 -725
rect 18175 -827 18209 -795
rect 18175 -829 18209 -827
rect 18290 -736 18324 -702
rect 18290 -804 18324 -774
rect 18290 -808 18324 -804
rect 18290 -872 18324 -846
rect 18290 -880 18324 -872
rect 856 -940 890 -918
rect 856 -952 890 -940
rect 1064 -957 1066 -923
rect 1066 -957 1098 -923
rect 1136 -957 1168 -923
rect 1168 -957 1170 -923
rect 1516 -957 1518 -923
rect 1518 -957 1550 -923
rect 1588 -957 1620 -923
rect 1620 -957 1622 -923
rect 1774 -957 1776 -923
rect 1776 -957 1808 -923
rect 1846 -957 1878 -923
rect 1878 -957 1880 -923
rect 2032 -957 2034 -923
rect 2034 -957 2066 -923
rect 2104 -957 2136 -923
rect 2136 -957 2138 -923
rect 2290 -957 2292 -923
rect 2292 -957 2324 -923
rect 2362 -957 2394 -923
rect 2394 -957 2396 -923
rect 2742 -957 2744 -923
rect 2744 -957 2776 -923
rect 2814 -957 2846 -923
rect 2846 -957 2848 -923
rect 3000 -957 3002 -923
rect 3002 -957 3034 -923
rect 3072 -957 3104 -923
rect 3104 -957 3106 -923
rect 3258 -957 3260 -923
rect 3260 -957 3292 -923
rect 3330 -957 3362 -923
rect 3362 -957 3364 -923
rect 3710 -957 3712 -923
rect 3712 -957 3744 -923
rect 3782 -957 3814 -923
rect 3814 -957 3816 -923
rect 3968 -957 3970 -923
rect 3970 -957 4002 -923
rect 4040 -957 4072 -923
rect 4072 -957 4074 -923
rect 4226 -957 4228 -923
rect 4228 -957 4260 -923
rect 4298 -957 4330 -923
rect 4330 -957 4332 -923
rect 4484 -957 4486 -923
rect 4486 -957 4518 -923
rect 4556 -957 4588 -923
rect 4588 -957 4590 -923
rect 4935 -957 4937 -923
rect 4937 -957 4969 -923
rect 5007 -957 5039 -923
rect 5039 -957 5041 -923
rect 5214 -940 5248 -918
rect 5214 -952 5248 -940
rect 856 -1008 890 -990
rect 856 -1024 890 -1008
rect 856 -1076 890 -1062
rect 856 -1096 890 -1076
rect 856 -1144 890 -1134
rect 856 -1168 890 -1144
rect 856 -1212 890 -1206
rect 856 -1240 890 -1212
rect 856 -1280 890 -1278
rect 856 -1312 890 -1280
rect 5421 -957 5423 -923
rect 5423 -957 5455 -923
rect 5493 -957 5525 -923
rect 5525 -957 5527 -923
rect 5873 -957 5875 -923
rect 5875 -957 5907 -923
rect 5945 -957 5977 -923
rect 5977 -957 5979 -923
rect 6131 -957 6133 -923
rect 6133 -957 6165 -923
rect 6203 -957 6235 -923
rect 6235 -957 6237 -923
rect 6389 -957 6391 -923
rect 6391 -957 6423 -923
rect 6461 -957 6493 -923
rect 6493 -957 6495 -923
rect 6647 -957 6649 -923
rect 6649 -957 6681 -923
rect 6719 -957 6751 -923
rect 6751 -957 6753 -923
rect 7099 -957 7101 -923
rect 7101 -957 7133 -923
rect 7171 -957 7203 -923
rect 7203 -957 7205 -923
rect 7357 -957 7359 -923
rect 7359 -957 7391 -923
rect 7429 -957 7461 -923
rect 7461 -957 7463 -923
rect 7615 -957 7617 -923
rect 7617 -957 7649 -923
rect 7687 -957 7719 -923
rect 7719 -957 7721 -923
rect 8067 -957 8069 -923
rect 8069 -957 8101 -923
rect 8139 -957 8171 -923
rect 8171 -957 8173 -923
rect 8325 -957 8327 -923
rect 8327 -957 8359 -923
rect 8397 -957 8429 -923
rect 8429 -957 8431 -923
rect 8583 -957 8585 -923
rect 8585 -957 8617 -923
rect 8655 -957 8687 -923
rect 8687 -957 8689 -923
rect 8841 -957 8843 -923
rect 8843 -957 8875 -923
rect 8913 -957 8945 -923
rect 8945 -957 8947 -923
rect 9293 -957 9295 -923
rect 9295 -957 9327 -923
rect 9365 -957 9397 -923
rect 9397 -957 9399 -923
rect 9573 -940 9607 -918
rect 9573 -952 9607 -940
rect 5214 -1008 5248 -990
rect 5214 -1024 5248 -1008
rect 5214 -1076 5248 -1062
rect 5214 -1096 5248 -1076
rect 5214 -1144 5248 -1134
rect 5214 -1168 5248 -1144
rect 5214 -1212 5248 -1206
rect 5214 -1240 5248 -1212
rect 5214 -1280 5248 -1278
rect 1064 -1320 1066 -1286
rect 1066 -1320 1098 -1286
rect 1136 -1320 1168 -1286
rect 1168 -1320 1170 -1286
rect 1516 -1320 1518 -1286
rect 1518 -1320 1550 -1286
rect 1588 -1320 1620 -1286
rect 1620 -1320 1622 -1286
rect 1774 -1320 1776 -1286
rect 1776 -1320 1808 -1286
rect 1846 -1320 1878 -1286
rect 1878 -1320 1880 -1286
rect 2032 -1320 2034 -1286
rect 2034 -1320 2066 -1286
rect 2104 -1320 2136 -1286
rect 2136 -1320 2138 -1286
rect 2290 -1320 2292 -1286
rect 2292 -1320 2324 -1286
rect 2362 -1320 2394 -1286
rect 2394 -1320 2396 -1286
rect 2742 -1320 2744 -1286
rect 2744 -1320 2776 -1286
rect 2814 -1320 2846 -1286
rect 2846 -1320 2848 -1286
rect 3000 -1320 3002 -1286
rect 3002 -1320 3034 -1286
rect 3072 -1320 3104 -1286
rect 3104 -1320 3106 -1286
rect 3258 -1320 3260 -1286
rect 3260 -1320 3292 -1286
rect 3330 -1320 3362 -1286
rect 3362 -1320 3364 -1286
rect 3710 -1320 3712 -1286
rect 3712 -1320 3744 -1286
rect 3782 -1320 3814 -1286
rect 3814 -1320 3816 -1286
rect 3968 -1320 3970 -1286
rect 3970 -1320 4002 -1286
rect 4040 -1320 4072 -1286
rect 4072 -1320 4074 -1286
rect 4226 -1320 4228 -1286
rect 4228 -1320 4260 -1286
rect 4298 -1320 4330 -1286
rect 4330 -1320 4332 -1286
rect 4484 -1320 4486 -1286
rect 4486 -1320 4518 -1286
rect 4556 -1320 4588 -1286
rect 4588 -1320 4590 -1286
rect 4935 -1320 4937 -1286
rect 4937 -1320 4969 -1286
rect 5007 -1320 5039 -1286
rect 5039 -1320 5041 -1286
rect 5214 -1312 5248 -1280
rect 9781 -957 9783 -923
rect 9783 -957 9815 -923
rect 9853 -957 9885 -923
rect 9885 -957 9887 -923
rect 10233 -957 10235 -923
rect 10235 -957 10267 -923
rect 10305 -957 10337 -923
rect 10337 -957 10339 -923
rect 10491 -957 10493 -923
rect 10493 -957 10525 -923
rect 10563 -957 10595 -923
rect 10595 -957 10597 -923
rect 10749 -957 10751 -923
rect 10751 -957 10783 -923
rect 10821 -957 10853 -923
rect 10853 -957 10855 -923
rect 11007 -957 11009 -923
rect 11009 -957 11041 -923
rect 11079 -957 11111 -923
rect 11111 -957 11113 -923
rect 11459 -957 11461 -923
rect 11461 -957 11493 -923
rect 11531 -957 11563 -923
rect 11563 -957 11565 -923
rect 11717 -957 11719 -923
rect 11719 -957 11751 -923
rect 11789 -957 11821 -923
rect 11821 -957 11823 -923
rect 11975 -957 11977 -923
rect 11977 -957 12009 -923
rect 12047 -957 12079 -923
rect 12079 -957 12081 -923
rect 12427 -957 12429 -923
rect 12429 -957 12461 -923
rect 12499 -957 12531 -923
rect 12531 -957 12533 -923
rect 12685 -957 12687 -923
rect 12687 -957 12719 -923
rect 12757 -957 12789 -923
rect 12789 -957 12791 -923
rect 12943 -957 12945 -923
rect 12945 -957 12977 -923
rect 13015 -957 13047 -923
rect 13047 -957 13049 -923
rect 13201 -957 13203 -923
rect 13203 -957 13235 -923
rect 13273 -957 13305 -923
rect 13305 -957 13307 -923
rect 13653 -957 13655 -923
rect 13655 -957 13687 -923
rect 13725 -957 13757 -923
rect 13757 -957 13759 -923
rect 13932 -940 13966 -918
rect 13932 -952 13966 -940
rect 9573 -1008 9607 -990
rect 9573 -1024 9607 -1008
rect 9573 -1076 9607 -1062
rect 9573 -1096 9607 -1076
rect 9573 -1144 9607 -1134
rect 9573 -1168 9607 -1144
rect 9573 -1212 9607 -1206
rect 9573 -1240 9607 -1212
rect 9573 -1280 9607 -1278
rect 856 -1382 890 -1350
rect 5421 -1320 5423 -1286
rect 5423 -1320 5455 -1286
rect 5493 -1320 5525 -1286
rect 5525 -1320 5527 -1286
rect 5873 -1320 5875 -1286
rect 5875 -1320 5907 -1286
rect 5945 -1320 5977 -1286
rect 5977 -1320 5979 -1286
rect 6131 -1320 6133 -1286
rect 6133 -1320 6165 -1286
rect 6203 -1320 6235 -1286
rect 6235 -1320 6237 -1286
rect 6389 -1320 6391 -1286
rect 6391 -1320 6423 -1286
rect 6461 -1320 6493 -1286
rect 6493 -1320 6495 -1286
rect 6647 -1320 6649 -1286
rect 6649 -1320 6681 -1286
rect 6719 -1320 6751 -1286
rect 6751 -1320 6753 -1286
rect 7099 -1320 7101 -1286
rect 7101 -1320 7133 -1286
rect 7171 -1320 7203 -1286
rect 7203 -1320 7205 -1286
rect 7357 -1320 7359 -1286
rect 7359 -1320 7391 -1286
rect 7429 -1320 7461 -1286
rect 7461 -1320 7463 -1286
rect 7615 -1320 7617 -1286
rect 7617 -1320 7649 -1286
rect 7687 -1320 7719 -1286
rect 7719 -1320 7721 -1286
rect 8067 -1320 8069 -1286
rect 8069 -1320 8101 -1286
rect 8139 -1320 8171 -1286
rect 8171 -1320 8173 -1286
rect 8325 -1320 8327 -1286
rect 8327 -1320 8359 -1286
rect 8397 -1320 8429 -1286
rect 8429 -1320 8431 -1286
rect 8583 -1320 8585 -1286
rect 8585 -1320 8617 -1286
rect 8655 -1320 8687 -1286
rect 8687 -1320 8689 -1286
rect 8841 -1320 8843 -1286
rect 8843 -1320 8875 -1286
rect 8913 -1320 8945 -1286
rect 8945 -1320 8947 -1286
rect 9293 -1320 9295 -1286
rect 9295 -1320 9327 -1286
rect 9365 -1320 9397 -1286
rect 9397 -1320 9399 -1286
rect 9573 -1312 9607 -1280
rect 14139 -957 14141 -923
rect 14141 -957 14173 -923
rect 14211 -957 14243 -923
rect 14243 -957 14245 -923
rect 14590 -957 14592 -923
rect 14592 -957 14624 -923
rect 14662 -957 14694 -923
rect 14694 -957 14696 -923
rect 14848 -957 14850 -923
rect 14850 -957 14882 -923
rect 14920 -957 14952 -923
rect 14952 -957 14954 -923
rect 15106 -957 15108 -923
rect 15108 -957 15140 -923
rect 15178 -957 15210 -923
rect 15210 -957 15212 -923
rect 15364 -957 15366 -923
rect 15366 -957 15398 -923
rect 15436 -957 15468 -923
rect 15468 -957 15470 -923
rect 15816 -957 15818 -923
rect 15818 -957 15850 -923
rect 15888 -957 15920 -923
rect 15920 -957 15922 -923
rect 16074 -957 16076 -923
rect 16076 -957 16108 -923
rect 16146 -957 16178 -923
rect 16178 -957 16180 -923
rect 16332 -957 16334 -923
rect 16334 -957 16366 -923
rect 16404 -957 16436 -923
rect 16436 -957 16438 -923
rect 16784 -957 16786 -923
rect 16786 -957 16818 -923
rect 16856 -957 16888 -923
rect 16888 -957 16890 -923
rect 17042 -957 17044 -923
rect 17044 -957 17076 -923
rect 17114 -957 17146 -923
rect 17146 -957 17148 -923
rect 17300 -957 17302 -923
rect 17302 -957 17334 -923
rect 17372 -957 17404 -923
rect 17404 -957 17406 -923
rect 17558 -957 17560 -923
rect 17560 -957 17592 -923
rect 17630 -957 17662 -923
rect 17662 -957 17664 -923
rect 18010 -957 18012 -923
rect 18012 -957 18044 -923
rect 18082 -957 18114 -923
rect 18114 -957 18116 -923
rect 18290 -940 18324 -918
rect 18290 -952 18324 -940
rect 13932 -1008 13966 -990
rect 13932 -1024 13966 -1008
rect 13932 -1076 13966 -1062
rect 13932 -1096 13966 -1076
rect 13932 -1144 13966 -1134
rect 13932 -1168 13966 -1144
rect 13932 -1212 13966 -1206
rect 13932 -1240 13966 -1212
rect 856 -1384 890 -1382
rect 856 -1450 890 -1422
rect 856 -1456 890 -1450
rect 856 -1518 890 -1494
rect 856 -1528 890 -1518
rect 856 -1586 890 -1566
rect 971 -1416 1005 -1414
rect 971 -1448 1005 -1416
rect 971 -1518 1005 -1486
rect 971 -1520 1005 -1518
rect 1229 -1416 1263 -1414
rect 1229 -1448 1263 -1416
rect 1229 -1518 1263 -1486
rect 1229 -1520 1263 -1518
rect 1423 -1416 1457 -1414
rect 1423 -1448 1457 -1416
rect 1423 -1518 1457 -1486
rect 1423 -1520 1457 -1518
rect 1681 -1416 1715 -1414
rect 1681 -1448 1715 -1416
rect 1681 -1518 1715 -1486
rect 1681 -1520 1715 -1518
rect 1939 -1416 1973 -1414
rect 1939 -1448 1973 -1416
rect 1939 -1518 1973 -1486
rect 1939 -1520 1973 -1518
rect 2197 -1416 2231 -1414
rect 2197 -1448 2231 -1416
rect 2197 -1518 2231 -1486
rect 2197 -1520 2231 -1518
rect 2455 -1416 2489 -1414
rect 2455 -1448 2489 -1416
rect 2455 -1518 2489 -1486
rect 2455 -1520 2489 -1518
rect 2649 -1416 2683 -1414
rect 2649 -1448 2683 -1416
rect 2649 -1518 2683 -1486
rect 2649 -1520 2683 -1518
rect 2907 -1416 2941 -1414
rect 2907 -1448 2941 -1416
rect 2907 -1518 2941 -1486
rect 2907 -1520 2941 -1518
rect 3165 -1416 3199 -1414
rect 3165 -1448 3199 -1416
rect 3165 -1518 3199 -1486
rect 3165 -1520 3199 -1518
rect 3423 -1416 3457 -1414
rect 3423 -1448 3457 -1416
rect 3423 -1518 3457 -1486
rect 3423 -1520 3457 -1518
rect 3617 -1416 3651 -1414
rect 3617 -1448 3651 -1416
rect 3617 -1518 3651 -1486
rect 3617 -1520 3651 -1518
rect 3875 -1416 3909 -1414
rect 3875 -1448 3909 -1416
rect 3875 -1518 3909 -1486
rect 3875 -1520 3909 -1518
rect 4133 -1416 4167 -1414
rect 4133 -1448 4167 -1416
rect 4133 -1518 4167 -1486
rect 4133 -1520 4167 -1518
rect 4391 -1416 4425 -1414
rect 4391 -1448 4425 -1416
rect 4391 -1518 4425 -1486
rect 4391 -1520 4425 -1518
rect 4649 -1416 4683 -1414
rect 4649 -1448 4683 -1416
rect 4649 -1518 4683 -1486
rect 4649 -1520 4683 -1518
rect 4842 -1416 4876 -1414
rect 4842 -1448 4876 -1416
rect 4842 -1518 4876 -1486
rect 4842 -1520 4876 -1518
rect 5100 -1416 5134 -1414
rect 5100 -1448 5134 -1416
rect 5100 -1518 5134 -1486
rect 5100 -1520 5134 -1518
rect 5214 -1382 5248 -1350
rect 5214 -1384 5248 -1382
rect 9781 -1320 9783 -1286
rect 9783 -1320 9815 -1286
rect 9853 -1320 9885 -1286
rect 9885 -1320 9887 -1286
rect 10233 -1320 10235 -1286
rect 10235 -1320 10267 -1286
rect 10305 -1320 10337 -1286
rect 10337 -1320 10339 -1286
rect 10491 -1320 10493 -1286
rect 10493 -1320 10525 -1286
rect 10563 -1320 10595 -1286
rect 10595 -1320 10597 -1286
rect 10749 -1320 10751 -1286
rect 10751 -1320 10783 -1286
rect 10821 -1320 10853 -1286
rect 10853 -1320 10855 -1286
rect 11007 -1320 11009 -1286
rect 11009 -1320 11041 -1286
rect 11079 -1320 11111 -1286
rect 11111 -1320 11113 -1286
rect 11459 -1320 11461 -1286
rect 11461 -1320 11493 -1286
rect 11531 -1320 11563 -1286
rect 11563 -1320 11565 -1286
rect 11717 -1320 11719 -1286
rect 11719 -1320 11751 -1286
rect 11789 -1320 11821 -1286
rect 11821 -1320 11823 -1286
rect 11975 -1320 11977 -1286
rect 11977 -1320 12009 -1286
rect 12047 -1320 12079 -1286
rect 12079 -1320 12081 -1286
rect 12427 -1320 12429 -1286
rect 12429 -1320 12461 -1286
rect 12499 -1320 12531 -1286
rect 12531 -1320 12533 -1286
rect 12685 -1320 12687 -1286
rect 12687 -1320 12719 -1286
rect 12757 -1320 12789 -1286
rect 12789 -1320 12791 -1286
rect 12943 -1320 12945 -1286
rect 12945 -1320 12977 -1286
rect 13015 -1320 13047 -1286
rect 13047 -1320 13049 -1286
rect 13201 -1320 13203 -1286
rect 13203 -1320 13235 -1286
rect 13273 -1320 13305 -1286
rect 13305 -1320 13307 -1286
rect 13653 -1320 13655 -1286
rect 13655 -1320 13687 -1286
rect 13725 -1320 13757 -1286
rect 13757 -1320 13759 -1286
rect 13932 -1280 13966 -1278
rect 13932 -1312 13966 -1280
rect 18290 -1008 18324 -990
rect 18290 -1024 18324 -1008
rect 18290 -1076 18324 -1062
rect 18290 -1096 18324 -1076
rect 18290 -1144 18324 -1134
rect 18290 -1168 18324 -1144
rect 18290 -1212 18324 -1206
rect 18290 -1240 18324 -1212
rect 18290 -1280 18324 -1278
rect 5214 -1450 5248 -1422
rect 5214 -1456 5248 -1450
rect 5214 -1518 5248 -1494
rect 5214 -1528 5248 -1518
rect 856 -1600 890 -1586
rect 856 -1654 890 -1638
rect 856 -1672 890 -1654
rect 856 -1722 890 -1710
rect 856 -1744 890 -1722
rect 856 -1790 890 -1782
rect 856 -1816 890 -1790
rect 856 -1888 890 -1854
rect 5214 -1586 5248 -1566
rect 5214 -1600 5248 -1586
rect 5328 -1416 5362 -1414
rect 5328 -1448 5362 -1416
rect 5328 -1518 5362 -1486
rect 5328 -1520 5362 -1518
rect 5586 -1416 5620 -1414
rect 5586 -1448 5620 -1416
rect 5586 -1518 5620 -1486
rect 5586 -1520 5620 -1518
rect 5780 -1416 5814 -1414
rect 5780 -1448 5814 -1416
rect 5780 -1518 5814 -1486
rect 5780 -1520 5814 -1518
rect 6038 -1416 6072 -1414
rect 6038 -1448 6072 -1416
rect 6038 -1518 6072 -1486
rect 6038 -1520 6072 -1518
rect 6296 -1416 6330 -1414
rect 6296 -1448 6330 -1416
rect 6296 -1518 6330 -1486
rect 6296 -1520 6330 -1518
rect 6554 -1416 6588 -1414
rect 6554 -1448 6588 -1416
rect 6554 -1518 6588 -1486
rect 6554 -1520 6588 -1518
rect 6812 -1416 6846 -1414
rect 6812 -1448 6846 -1416
rect 6812 -1518 6846 -1486
rect 6812 -1520 6846 -1518
rect 7006 -1416 7040 -1414
rect 7006 -1448 7040 -1416
rect 7006 -1518 7040 -1486
rect 7006 -1520 7040 -1518
rect 7264 -1416 7298 -1414
rect 7264 -1448 7298 -1416
rect 7264 -1518 7298 -1486
rect 7264 -1520 7298 -1518
rect 7522 -1416 7556 -1414
rect 7522 -1448 7556 -1416
rect 7522 -1518 7556 -1486
rect 7522 -1520 7556 -1518
rect 7780 -1416 7814 -1414
rect 7780 -1448 7814 -1416
rect 7780 -1518 7814 -1486
rect 7780 -1520 7814 -1518
rect 7974 -1416 8008 -1414
rect 7974 -1448 8008 -1416
rect 7974 -1518 8008 -1486
rect 7974 -1520 8008 -1518
rect 8232 -1416 8266 -1414
rect 8232 -1448 8266 -1416
rect 8232 -1518 8266 -1486
rect 8232 -1520 8266 -1518
rect 8490 -1416 8524 -1414
rect 8490 -1448 8524 -1416
rect 8490 -1518 8524 -1486
rect 8490 -1520 8524 -1518
rect 8748 -1416 8782 -1414
rect 8748 -1448 8782 -1416
rect 8748 -1518 8782 -1486
rect 8748 -1520 8782 -1518
rect 9006 -1416 9040 -1414
rect 9006 -1448 9040 -1416
rect 9006 -1518 9040 -1486
rect 9006 -1520 9040 -1518
rect 9200 -1416 9234 -1414
rect 9200 -1448 9234 -1416
rect 9200 -1518 9234 -1486
rect 9200 -1520 9234 -1518
rect 9458 -1416 9492 -1414
rect 9458 -1448 9492 -1416
rect 9458 -1518 9492 -1486
rect 9458 -1520 9492 -1518
rect 9573 -1382 9607 -1350
rect 14139 -1320 14141 -1286
rect 14141 -1320 14173 -1286
rect 14211 -1320 14243 -1286
rect 14243 -1320 14245 -1286
rect 14590 -1320 14592 -1286
rect 14592 -1320 14624 -1286
rect 14662 -1320 14694 -1286
rect 14694 -1320 14696 -1286
rect 14848 -1320 14850 -1286
rect 14850 -1320 14882 -1286
rect 14920 -1320 14952 -1286
rect 14952 -1320 14954 -1286
rect 15106 -1320 15108 -1286
rect 15108 -1320 15140 -1286
rect 15178 -1320 15210 -1286
rect 15210 -1320 15212 -1286
rect 15364 -1320 15366 -1286
rect 15366 -1320 15398 -1286
rect 15436 -1320 15468 -1286
rect 15468 -1320 15470 -1286
rect 15816 -1320 15818 -1286
rect 15818 -1320 15850 -1286
rect 15888 -1320 15920 -1286
rect 15920 -1320 15922 -1286
rect 16074 -1320 16076 -1286
rect 16076 -1320 16108 -1286
rect 16146 -1320 16178 -1286
rect 16178 -1320 16180 -1286
rect 16332 -1320 16334 -1286
rect 16334 -1320 16366 -1286
rect 16404 -1320 16436 -1286
rect 16436 -1320 16438 -1286
rect 16784 -1320 16786 -1286
rect 16786 -1320 16818 -1286
rect 16856 -1320 16888 -1286
rect 16888 -1320 16890 -1286
rect 17042 -1320 17044 -1286
rect 17044 -1320 17076 -1286
rect 17114 -1320 17146 -1286
rect 17146 -1320 17148 -1286
rect 17300 -1320 17302 -1286
rect 17302 -1320 17334 -1286
rect 17372 -1320 17404 -1286
rect 17404 -1320 17406 -1286
rect 17558 -1320 17560 -1286
rect 17560 -1320 17592 -1286
rect 17630 -1320 17662 -1286
rect 17662 -1320 17664 -1286
rect 18010 -1320 18012 -1286
rect 18012 -1320 18044 -1286
rect 18082 -1320 18114 -1286
rect 18114 -1320 18116 -1286
rect 18290 -1312 18324 -1280
rect 9573 -1384 9607 -1382
rect 9573 -1450 9607 -1422
rect 9573 -1456 9607 -1450
rect 9573 -1518 9607 -1494
rect 9573 -1528 9607 -1518
rect 5214 -1654 5248 -1638
rect 5214 -1672 5248 -1654
rect 5214 -1722 5248 -1710
rect 5214 -1744 5248 -1722
rect 5214 -1790 5248 -1782
rect 5214 -1816 5248 -1790
rect 5214 -1888 5248 -1854
rect 9573 -1586 9607 -1566
rect 9688 -1416 9722 -1414
rect 9688 -1448 9722 -1416
rect 9688 -1518 9722 -1486
rect 9688 -1520 9722 -1518
rect 9946 -1416 9980 -1414
rect 9946 -1448 9980 -1416
rect 9946 -1518 9980 -1486
rect 9946 -1520 9980 -1518
rect 10140 -1416 10174 -1414
rect 10140 -1448 10174 -1416
rect 10140 -1518 10174 -1486
rect 10140 -1520 10174 -1518
rect 10398 -1416 10432 -1414
rect 10398 -1448 10432 -1416
rect 10398 -1518 10432 -1486
rect 10398 -1520 10432 -1518
rect 10656 -1416 10690 -1414
rect 10656 -1448 10690 -1416
rect 10656 -1518 10690 -1486
rect 10656 -1520 10690 -1518
rect 10914 -1416 10948 -1414
rect 10914 -1448 10948 -1416
rect 10914 -1518 10948 -1486
rect 10914 -1520 10948 -1518
rect 11172 -1416 11206 -1414
rect 11172 -1448 11206 -1416
rect 11172 -1518 11206 -1486
rect 11172 -1520 11206 -1518
rect 11366 -1416 11400 -1414
rect 11366 -1448 11400 -1416
rect 11366 -1518 11400 -1486
rect 11366 -1520 11400 -1518
rect 11624 -1416 11658 -1414
rect 11624 -1448 11658 -1416
rect 11624 -1518 11658 -1486
rect 11624 -1520 11658 -1518
rect 11882 -1416 11916 -1414
rect 11882 -1448 11916 -1416
rect 11882 -1518 11916 -1486
rect 11882 -1520 11916 -1518
rect 12140 -1416 12174 -1414
rect 12140 -1448 12174 -1416
rect 12140 -1518 12174 -1486
rect 12140 -1520 12174 -1518
rect 12334 -1416 12368 -1414
rect 12334 -1448 12368 -1416
rect 12334 -1518 12368 -1486
rect 12334 -1520 12368 -1518
rect 12592 -1416 12626 -1414
rect 12592 -1448 12626 -1416
rect 12592 -1518 12626 -1486
rect 12592 -1520 12626 -1518
rect 12850 -1416 12884 -1414
rect 12850 -1448 12884 -1416
rect 12850 -1518 12884 -1486
rect 12850 -1520 12884 -1518
rect 13108 -1416 13142 -1414
rect 13108 -1448 13142 -1416
rect 13108 -1518 13142 -1486
rect 13108 -1520 13142 -1518
rect 13366 -1416 13400 -1414
rect 13366 -1448 13400 -1416
rect 13366 -1518 13400 -1486
rect 13366 -1520 13400 -1518
rect 13560 -1416 13594 -1414
rect 13560 -1448 13594 -1416
rect 13560 -1518 13594 -1486
rect 13560 -1520 13594 -1518
rect 13818 -1416 13852 -1414
rect 13818 -1448 13852 -1416
rect 13818 -1518 13852 -1486
rect 13818 -1520 13852 -1518
rect 13932 -1382 13966 -1350
rect 13932 -1384 13966 -1382
rect 13932 -1450 13966 -1422
rect 13932 -1456 13966 -1450
rect 13932 -1518 13966 -1494
rect 13932 -1528 13966 -1518
rect 9573 -1600 9607 -1586
rect 9573 -1654 9607 -1638
rect 9573 -1672 9607 -1654
rect 9573 -1722 9607 -1710
rect 9573 -1744 9607 -1722
rect 9573 -1790 9607 -1782
rect 9573 -1816 9607 -1790
rect 9573 -1888 9607 -1854
rect 13932 -1586 13966 -1566
rect 14046 -1416 14080 -1414
rect 14046 -1448 14080 -1416
rect 14046 -1518 14080 -1486
rect 14046 -1520 14080 -1518
rect 14304 -1416 14338 -1414
rect 14304 -1448 14338 -1416
rect 14304 -1518 14338 -1486
rect 14304 -1520 14338 -1518
rect 14497 -1416 14531 -1414
rect 14497 -1448 14531 -1416
rect 14497 -1518 14531 -1486
rect 14497 -1520 14531 -1518
rect 14755 -1416 14789 -1414
rect 14755 -1448 14789 -1416
rect 14755 -1518 14789 -1486
rect 14755 -1520 14789 -1518
rect 15013 -1416 15047 -1414
rect 15013 -1448 15047 -1416
rect 15013 -1518 15047 -1486
rect 15013 -1520 15047 -1518
rect 15271 -1416 15305 -1414
rect 15271 -1448 15305 -1416
rect 15271 -1518 15305 -1486
rect 15271 -1520 15305 -1518
rect 15529 -1416 15563 -1414
rect 15529 -1448 15563 -1416
rect 15529 -1518 15563 -1486
rect 15529 -1520 15563 -1518
rect 15723 -1416 15757 -1414
rect 15723 -1448 15757 -1416
rect 15723 -1518 15757 -1486
rect 15723 -1520 15757 -1518
rect 15981 -1416 16015 -1414
rect 15981 -1448 16015 -1416
rect 15981 -1518 16015 -1486
rect 15981 -1520 16015 -1518
rect 16239 -1416 16273 -1414
rect 16239 -1448 16273 -1416
rect 16239 -1518 16273 -1486
rect 16239 -1520 16273 -1518
rect 16497 -1416 16531 -1414
rect 16497 -1448 16531 -1416
rect 16497 -1518 16531 -1486
rect 16497 -1520 16531 -1518
rect 16691 -1416 16725 -1414
rect 16691 -1448 16725 -1416
rect 16691 -1518 16725 -1486
rect 16691 -1520 16725 -1518
rect 16949 -1416 16983 -1414
rect 16949 -1448 16983 -1416
rect 16949 -1518 16983 -1486
rect 16949 -1520 16983 -1518
rect 17207 -1416 17241 -1414
rect 17207 -1448 17241 -1416
rect 17207 -1518 17241 -1486
rect 17207 -1520 17241 -1518
rect 17465 -1416 17499 -1414
rect 17465 -1448 17499 -1416
rect 17465 -1518 17499 -1486
rect 17465 -1520 17499 -1518
rect 17723 -1416 17757 -1414
rect 17723 -1448 17757 -1416
rect 17723 -1518 17757 -1486
rect 17723 -1520 17757 -1518
rect 17917 -1416 17951 -1414
rect 17917 -1448 17951 -1416
rect 17917 -1518 17951 -1486
rect 17917 -1520 17951 -1518
rect 18175 -1416 18209 -1414
rect 18175 -1448 18209 -1416
rect 18175 -1518 18209 -1486
rect 18175 -1520 18209 -1518
rect 18290 -1382 18324 -1350
rect 18290 -1384 18324 -1382
rect 18290 -1450 18324 -1422
rect 18290 -1456 18324 -1450
rect 18290 -1518 18324 -1494
rect 18290 -1528 18324 -1518
rect 13932 -1600 13966 -1586
rect 13932 -1654 13966 -1638
rect 13932 -1672 13966 -1654
rect 13932 -1722 13966 -1710
rect 13932 -1744 13966 -1722
rect 13932 -1790 13966 -1782
rect 13932 -1816 13966 -1790
rect 13932 -1888 13966 -1854
rect 18290 -1586 18324 -1566
rect 18290 -1600 18324 -1586
rect 18290 -1654 18324 -1638
rect 18290 -1672 18324 -1654
rect 18290 -1722 18324 -1710
rect 18290 -1744 18324 -1722
rect 18290 -1790 18324 -1782
rect 18290 -1816 18324 -1790
rect 18290 -1888 18324 -1854
rect 856 -1960 890 -1926
rect 5214 -1960 5248 -1926
rect 9573 -1960 9607 -1926
rect 13932 -1960 13966 -1926
rect 18290 -1960 18324 -1926
rect 856 -2032 890 -1998
rect 856 -2096 890 -2070
rect 856 -2104 890 -2096
rect 856 -2164 890 -2142
rect 856 -2176 890 -2164
rect 856 -2232 890 -2214
rect 856 -2248 890 -2232
rect 856 -2300 890 -2286
rect 856 -2320 890 -2300
rect 5214 -2032 5248 -1998
rect 5214 -2096 5248 -2070
rect 5214 -2104 5248 -2096
rect 5214 -2164 5248 -2142
rect 5214 -2176 5248 -2164
rect 5214 -2232 5248 -2214
rect 5214 -2248 5248 -2232
rect 5214 -2300 5248 -2286
rect 856 -2368 890 -2358
rect 856 -2392 890 -2368
rect 856 -2436 890 -2430
rect 856 -2464 890 -2436
rect 856 -2504 890 -2502
rect 856 -2536 890 -2504
rect 971 -2372 1005 -2370
rect 971 -2404 1005 -2372
rect 971 -2474 1005 -2442
rect 971 -2476 1005 -2474
rect 1229 -2372 1263 -2370
rect 1229 -2404 1263 -2372
rect 1229 -2474 1263 -2442
rect 1229 -2476 1263 -2474
rect 1423 -2372 1457 -2370
rect 1423 -2404 1457 -2372
rect 1423 -2474 1457 -2442
rect 1423 -2476 1457 -2474
rect 1681 -2372 1715 -2370
rect 1681 -2404 1715 -2372
rect 1681 -2474 1715 -2442
rect 1681 -2476 1715 -2474
rect 1939 -2372 1973 -2370
rect 1939 -2404 1973 -2372
rect 1939 -2474 1973 -2442
rect 1939 -2476 1973 -2474
rect 2197 -2372 2231 -2370
rect 2197 -2404 2231 -2372
rect 2197 -2474 2231 -2442
rect 2197 -2476 2231 -2474
rect 2455 -2372 2489 -2370
rect 2455 -2404 2489 -2372
rect 2455 -2474 2489 -2442
rect 2455 -2476 2489 -2474
rect 2649 -2372 2683 -2370
rect 2649 -2404 2683 -2372
rect 2649 -2474 2683 -2442
rect 2649 -2476 2683 -2474
rect 2907 -2372 2941 -2370
rect 2907 -2404 2941 -2372
rect 2907 -2474 2941 -2442
rect 2907 -2476 2941 -2474
rect 3165 -2372 3199 -2370
rect 3165 -2404 3199 -2372
rect 3165 -2474 3199 -2442
rect 3165 -2476 3199 -2474
rect 3423 -2372 3457 -2370
rect 3423 -2404 3457 -2372
rect 3423 -2474 3457 -2442
rect 3423 -2476 3457 -2474
rect 3617 -2372 3651 -2370
rect 3617 -2404 3651 -2372
rect 3617 -2474 3651 -2442
rect 3617 -2476 3651 -2474
rect 3875 -2372 3909 -2370
rect 3875 -2404 3909 -2372
rect 3875 -2474 3909 -2442
rect 3875 -2476 3909 -2474
rect 4133 -2372 4167 -2370
rect 4133 -2404 4167 -2372
rect 4133 -2474 4167 -2442
rect 4133 -2476 4167 -2474
rect 4391 -2372 4425 -2370
rect 4391 -2404 4425 -2372
rect 4391 -2474 4425 -2442
rect 4391 -2476 4425 -2474
rect 4649 -2372 4683 -2370
rect 4649 -2404 4683 -2372
rect 4649 -2474 4683 -2442
rect 4649 -2476 4683 -2474
rect 4842 -2372 4876 -2370
rect 4842 -2404 4876 -2372
rect 4842 -2474 4876 -2442
rect 4842 -2476 4876 -2474
rect 5100 -2372 5134 -2370
rect 5100 -2404 5134 -2372
rect 5100 -2474 5134 -2442
rect 5100 -2476 5134 -2474
rect 5214 -2320 5248 -2300
rect 9573 -2032 9607 -1998
rect 9573 -2096 9607 -2070
rect 9573 -2104 9607 -2096
rect 9573 -2164 9607 -2142
rect 9573 -2176 9607 -2164
rect 9573 -2232 9607 -2214
rect 9573 -2248 9607 -2232
rect 9573 -2300 9607 -2286
rect 5214 -2368 5248 -2358
rect 5214 -2392 5248 -2368
rect 5214 -2436 5248 -2430
rect 5214 -2464 5248 -2436
rect 5214 -2504 5248 -2502
rect 5214 -2536 5248 -2504
rect 5328 -2372 5362 -2370
rect 5328 -2404 5362 -2372
rect 5328 -2474 5362 -2442
rect 5328 -2476 5362 -2474
rect 5586 -2372 5620 -2370
rect 5586 -2404 5620 -2372
rect 5586 -2474 5620 -2442
rect 5586 -2476 5620 -2474
rect 5780 -2372 5814 -2370
rect 5780 -2404 5814 -2372
rect 5780 -2474 5814 -2442
rect 5780 -2476 5814 -2474
rect 6038 -2372 6072 -2370
rect 6038 -2404 6072 -2372
rect 6038 -2474 6072 -2442
rect 6038 -2476 6072 -2474
rect 6296 -2372 6330 -2370
rect 6296 -2404 6330 -2372
rect 6296 -2474 6330 -2442
rect 6296 -2476 6330 -2474
rect 6554 -2372 6588 -2370
rect 6554 -2404 6588 -2372
rect 6554 -2474 6588 -2442
rect 6554 -2476 6588 -2474
rect 6812 -2372 6846 -2370
rect 6812 -2404 6846 -2372
rect 6812 -2474 6846 -2442
rect 6812 -2476 6846 -2474
rect 7006 -2372 7040 -2370
rect 7006 -2404 7040 -2372
rect 7006 -2474 7040 -2442
rect 7006 -2476 7040 -2474
rect 7264 -2372 7298 -2370
rect 7264 -2404 7298 -2372
rect 7264 -2474 7298 -2442
rect 7264 -2476 7298 -2474
rect 7522 -2372 7556 -2370
rect 7522 -2404 7556 -2372
rect 7522 -2474 7556 -2442
rect 7522 -2476 7556 -2474
rect 7780 -2372 7814 -2370
rect 7780 -2404 7814 -2372
rect 7780 -2474 7814 -2442
rect 7780 -2476 7814 -2474
rect 7974 -2372 8008 -2370
rect 7974 -2404 8008 -2372
rect 7974 -2474 8008 -2442
rect 7974 -2476 8008 -2474
rect 8232 -2372 8266 -2370
rect 8232 -2404 8266 -2372
rect 8232 -2474 8266 -2442
rect 8232 -2476 8266 -2474
rect 8490 -2372 8524 -2370
rect 8490 -2404 8524 -2372
rect 8490 -2474 8524 -2442
rect 8490 -2476 8524 -2474
rect 8748 -2372 8782 -2370
rect 8748 -2404 8782 -2372
rect 8748 -2474 8782 -2442
rect 8748 -2476 8782 -2474
rect 9006 -2372 9040 -2370
rect 9006 -2404 9040 -2372
rect 9006 -2474 9040 -2442
rect 9006 -2476 9040 -2474
rect 9200 -2372 9234 -2370
rect 9200 -2404 9234 -2372
rect 9200 -2474 9234 -2442
rect 9200 -2476 9234 -2474
rect 9458 -2372 9492 -2370
rect 9458 -2404 9492 -2372
rect 9458 -2474 9492 -2442
rect 9458 -2476 9492 -2474
rect 9573 -2320 9607 -2300
rect 13932 -2032 13966 -1998
rect 13932 -2096 13966 -2070
rect 13932 -2104 13966 -2096
rect 13932 -2164 13966 -2142
rect 13932 -2176 13966 -2164
rect 13932 -2232 13966 -2214
rect 13932 -2248 13966 -2232
rect 9573 -2368 9607 -2358
rect 9573 -2392 9607 -2368
rect 9573 -2436 9607 -2430
rect 9573 -2464 9607 -2436
rect 9573 -2504 9607 -2502
rect 856 -2606 890 -2574
rect 1064 -2604 1066 -2570
rect 1066 -2604 1098 -2570
rect 1136 -2604 1168 -2570
rect 1168 -2604 1170 -2570
rect 1516 -2604 1518 -2570
rect 1518 -2604 1550 -2570
rect 1588 -2604 1620 -2570
rect 1620 -2604 1622 -2570
rect 1774 -2604 1776 -2570
rect 1776 -2604 1808 -2570
rect 1846 -2604 1878 -2570
rect 1878 -2604 1880 -2570
rect 2032 -2604 2034 -2570
rect 2034 -2604 2066 -2570
rect 2104 -2604 2136 -2570
rect 2136 -2604 2138 -2570
rect 2290 -2604 2292 -2570
rect 2292 -2604 2324 -2570
rect 2362 -2604 2394 -2570
rect 2394 -2604 2396 -2570
rect 2742 -2604 2744 -2570
rect 2744 -2604 2776 -2570
rect 2814 -2604 2846 -2570
rect 2846 -2604 2848 -2570
rect 3000 -2604 3002 -2570
rect 3002 -2604 3034 -2570
rect 3072 -2604 3104 -2570
rect 3104 -2604 3106 -2570
rect 3258 -2604 3260 -2570
rect 3260 -2604 3292 -2570
rect 3330 -2604 3362 -2570
rect 3362 -2604 3364 -2570
rect 3710 -2604 3712 -2570
rect 3712 -2604 3744 -2570
rect 3782 -2604 3814 -2570
rect 3814 -2604 3816 -2570
rect 3968 -2604 3970 -2570
rect 3970 -2604 4002 -2570
rect 4040 -2604 4072 -2570
rect 4072 -2604 4074 -2570
rect 4226 -2604 4228 -2570
rect 4228 -2604 4260 -2570
rect 4298 -2604 4330 -2570
rect 4330 -2604 4332 -2570
rect 4484 -2604 4486 -2570
rect 4486 -2604 4518 -2570
rect 4556 -2604 4588 -2570
rect 4588 -2604 4590 -2570
rect 4935 -2604 4937 -2570
rect 4937 -2604 4969 -2570
rect 5007 -2604 5039 -2570
rect 5039 -2604 5041 -2570
rect 9573 -2536 9607 -2504
rect 9688 -2372 9722 -2370
rect 9688 -2404 9722 -2372
rect 9688 -2474 9722 -2442
rect 9688 -2476 9722 -2474
rect 9946 -2372 9980 -2370
rect 9946 -2404 9980 -2372
rect 9946 -2474 9980 -2442
rect 9946 -2476 9980 -2474
rect 10140 -2372 10174 -2370
rect 10140 -2404 10174 -2372
rect 10140 -2474 10174 -2442
rect 10140 -2476 10174 -2474
rect 10398 -2372 10432 -2370
rect 10398 -2404 10432 -2372
rect 10398 -2474 10432 -2442
rect 10398 -2476 10432 -2474
rect 10656 -2372 10690 -2370
rect 10656 -2404 10690 -2372
rect 10656 -2474 10690 -2442
rect 10656 -2476 10690 -2474
rect 10914 -2372 10948 -2370
rect 10914 -2404 10948 -2372
rect 10914 -2474 10948 -2442
rect 10914 -2476 10948 -2474
rect 11172 -2372 11206 -2370
rect 11172 -2404 11206 -2372
rect 11172 -2474 11206 -2442
rect 11172 -2476 11206 -2474
rect 11366 -2372 11400 -2370
rect 11366 -2404 11400 -2372
rect 11366 -2474 11400 -2442
rect 11366 -2476 11400 -2474
rect 11624 -2372 11658 -2370
rect 11624 -2404 11658 -2372
rect 11624 -2474 11658 -2442
rect 11624 -2476 11658 -2474
rect 11882 -2372 11916 -2370
rect 11882 -2404 11916 -2372
rect 11882 -2474 11916 -2442
rect 11882 -2476 11916 -2474
rect 12140 -2372 12174 -2370
rect 12140 -2404 12174 -2372
rect 12140 -2474 12174 -2442
rect 12140 -2476 12174 -2474
rect 12334 -2372 12368 -2370
rect 12334 -2404 12368 -2372
rect 12334 -2474 12368 -2442
rect 12334 -2476 12368 -2474
rect 12592 -2372 12626 -2370
rect 12592 -2404 12626 -2372
rect 12592 -2474 12626 -2442
rect 12592 -2476 12626 -2474
rect 12850 -2372 12884 -2370
rect 12850 -2404 12884 -2372
rect 12850 -2474 12884 -2442
rect 12850 -2476 12884 -2474
rect 13108 -2372 13142 -2370
rect 13108 -2404 13142 -2372
rect 13108 -2474 13142 -2442
rect 13108 -2476 13142 -2474
rect 13366 -2372 13400 -2370
rect 13366 -2404 13400 -2372
rect 13366 -2474 13400 -2442
rect 13366 -2476 13400 -2474
rect 13560 -2372 13594 -2370
rect 13560 -2404 13594 -2372
rect 13560 -2474 13594 -2442
rect 13560 -2476 13594 -2474
rect 13818 -2372 13852 -2370
rect 13818 -2404 13852 -2372
rect 13818 -2474 13852 -2442
rect 13818 -2476 13852 -2474
rect 13932 -2300 13966 -2286
rect 13932 -2320 13966 -2300
rect 18290 -2032 18324 -1998
rect 18290 -2096 18324 -2070
rect 18290 -2104 18324 -2096
rect 18290 -2164 18324 -2142
rect 18290 -2176 18324 -2164
rect 18290 -2232 18324 -2214
rect 18290 -2248 18324 -2232
rect 18290 -2300 18324 -2286
rect 13932 -2368 13966 -2358
rect 13932 -2392 13966 -2368
rect 13932 -2436 13966 -2430
rect 13932 -2464 13966 -2436
rect 856 -2608 890 -2606
rect 856 -2674 890 -2646
rect 856 -2680 890 -2674
rect 856 -2742 890 -2718
rect 856 -2752 890 -2742
rect 856 -2810 890 -2790
rect 856 -2824 890 -2810
rect 856 -2878 890 -2862
rect 856 -2896 890 -2878
rect 5214 -2606 5248 -2574
rect 5214 -2608 5248 -2606
rect 5421 -2604 5423 -2570
rect 5423 -2604 5455 -2570
rect 5493 -2604 5525 -2570
rect 5525 -2604 5527 -2570
rect 5873 -2604 5875 -2570
rect 5875 -2604 5907 -2570
rect 5945 -2604 5977 -2570
rect 5977 -2604 5979 -2570
rect 6131 -2604 6133 -2570
rect 6133 -2604 6165 -2570
rect 6203 -2604 6235 -2570
rect 6235 -2604 6237 -2570
rect 6389 -2604 6391 -2570
rect 6391 -2604 6423 -2570
rect 6461 -2604 6493 -2570
rect 6493 -2604 6495 -2570
rect 6647 -2604 6649 -2570
rect 6649 -2604 6681 -2570
rect 6719 -2604 6751 -2570
rect 6751 -2604 6753 -2570
rect 7099 -2604 7101 -2570
rect 7101 -2604 7133 -2570
rect 7171 -2604 7203 -2570
rect 7203 -2604 7205 -2570
rect 7357 -2604 7359 -2570
rect 7359 -2604 7391 -2570
rect 7429 -2604 7461 -2570
rect 7461 -2604 7463 -2570
rect 7615 -2604 7617 -2570
rect 7617 -2604 7649 -2570
rect 7687 -2604 7719 -2570
rect 7719 -2604 7721 -2570
rect 8067 -2604 8069 -2570
rect 8069 -2604 8101 -2570
rect 8139 -2604 8171 -2570
rect 8171 -2604 8173 -2570
rect 8325 -2604 8327 -2570
rect 8327 -2604 8359 -2570
rect 8397 -2604 8429 -2570
rect 8429 -2604 8431 -2570
rect 8583 -2604 8585 -2570
rect 8585 -2604 8617 -2570
rect 8655 -2604 8687 -2570
rect 8687 -2604 8689 -2570
rect 8841 -2604 8843 -2570
rect 8843 -2604 8875 -2570
rect 8913 -2604 8945 -2570
rect 8945 -2604 8947 -2570
rect 9293 -2604 9295 -2570
rect 9295 -2604 9327 -2570
rect 9365 -2604 9397 -2570
rect 9397 -2604 9399 -2570
rect 13932 -2504 13966 -2502
rect 13932 -2536 13966 -2504
rect 14046 -2372 14080 -2370
rect 14046 -2404 14080 -2372
rect 14046 -2474 14080 -2442
rect 14046 -2476 14080 -2474
rect 14304 -2372 14338 -2370
rect 14304 -2404 14338 -2372
rect 14304 -2474 14338 -2442
rect 14304 -2476 14338 -2474
rect 14497 -2372 14531 -2370
rect 14497 -2404 14531 -2372
rect 14497 -2474 14531 -2442
rect 14497 -2476 14531 -2474
rect 14755 -2372 14789 -2370
rect 14755 -2404 14789 -2372
rect 14755 -2474 14789 -2442
rect 14755 -2476 14789 -2474
rect 15013 -2372 15047 -2370
rect 15013 -2404 15047 -2372
rect 15013 -2474 15047 -2442
rect 15013 -2476 15047 -2474
rect 15271 -2372 15305 -2370
rect 15271 -2404 15305 -2372
rect 15271 -2474 15305 -2442
rect 15271 -2476 15305 -2474
rect 15529 -2372 15563 -2370
rect 15529 -2404 15563 -2372
rect 15529 -2474 15563 -2442
rect 15529 -2476 15563 -2474
rect 15723 -2372 15757 -2370
rect 15723 -2404 15757 -2372
rect 15723 -2474 15757 -2442
rect 15723 -2476 15757 -2474
rect 15981 -2372 16015 -2370
rect 15981 -2404 16015 -2372
rect 15981 -2474 16015 -2442
rect 15981 -2476 16015 -2474
rect 16239 -2372 16273 -2370
rect 16239 -2404 16273 -2372
rect 16239 -2474 16273 -2442
rect 16239 -2476 16273 -2474
rect 16497 -2372 16531 -2370
rect 16497 -2404 16531 -2372
rect 16497 -2474 16531 -2442
rect 16497 -2476 16531 -2474
rect 16691 -2372 16725 -2370
rect 16691 -2404 16725 -2372
rect 16691 -2474 16725 -2442
rect 16691 -2476 16725 -2474
rect 16949 -2372 16983 -2370
rect 16949 -2404 16983 -2372
rect 16949 -2474 16983 -2442
rect 16949 -2476 16983 -2474
rect 17207 -2372 17241 -2370
rect 17207 -2404 17241 -2372
rect 17207 -2474 17241 -2442
rect 17207 -2476 17241 -2474
rect 17465 -2372 17499 -2370
rect 17465 -2404 17499 -2372
rect 17465 -2474 17499 -2442
rect 17465 -2476 17499 -2474
rect 17723 -2372 17757 -2370
rect 17723 -2404 17757 -2372
rect 17723 -2474 17757 -2442
rect 17723 -2476 17757 -2474
rect 17917 -2372 17951 -2370
rect 17917 -2404 17951 -2372
rect 17917 -2474 17951 -2442
rect 17917 -2476 17951 -2474
rect 18175 -2372 18209 -2370
rect 18175 -2404 18209 -2372
rect 18175 -2474 18209 -2442
rect 18175 -2476 18209 -2474
rect 18290 -2320 18324 -2300
rect 18290 -2368 18324 -2358
rect 18290 -2392 18324 -2368
rect 18290 -2436 18324 -2430
rect 18290 -2464 18324 -2436
rect 18290 -2504 18324 -2502
rect 5214 -2674 5248 -2646
rect 5214 -2680 5248 -2674
rect 5214 -2742 5248 -2718
rect 5214 -2752 5248 -2742
rect 5214 -2810 5248 -2790
rect 5214 -2824 5248 -2810
rect 5214 -2878 5248 -2862
rect 5214 -2896 5248 -2878
rect 856 -2946 890 -2934
rect 856 -2968 890 -2946
rect 1064 -2967 1066 -2933
rect 1066 -2967 1098 -2933
rect 1136 -2967 1168 -2933
rect 1168 -2967 1170 -2933
rect 1516 -2967 1518 -2933
rect 1518 -2967 1550 -2933
rect 1588 -2967 1620 -2933
rect 1620 -2967 1622 -2933
rect 1774 -2967 1776 -2933
rect 1776 -2967 1808 -2933
rect 1846 -2967 1878 -2933
rect 1878 -2967 1880 -2933
rect 2032 -2967 2034 -2933
rect 2034 -2967 2066 -2933
rect 2104 -2967 2136 -2933
rect 2136 -2967 2138 -2933
rect 2290 -2967 2292 -2933
rect 2292 -2967 2324 -2933
rect 2362 -2967 2394 -2933
rect 2394 -2967 2396 -2933
rect 2742 -2967 2744 -2933
rect 2744 -2967 2776 -2933
rect 2814 -2967 2846 -2933
rect 2846 -2967 2848 -2933
rect 3000 -2967 3002 -2933
rect 3002 -2967 3034 -2933
rect 3072 -2967 3104 -2933
rect 3104 -2967 3106 -2933
rect 3258 -2967 3260 -2933
rect 3260 -2967 3292 -2933
rect 3330 -2967 3362 -2933
rect 3362 -2967 3364 -2933
rect 3710 -2967 3712 -2933
rect 3712 -2967 3744 -2933
rect 3782 -2967 3814 -2933
rect 3814 -2967 3816 -2933
rect 3968 -2967 3970 -2933
rect 3970 -2967 4002 -2933
rect 4040 -2967 4072 -2933
rect 4072 -2967 4074 -2933
rect 4226 -2967 4228 -2933
rect 4228 -2967 4260 -2933
rect 4298 -2967 4330 -2933
rect 4330 -2967 4332 -2933
rect 4484 -2967 4486 -2933
rect 4486 -2967 4518 -2933
rect 4556 -2967 4588 -2933
rect 4588 -2967 4590 -2933
rect 4935 -2967 4937 -2933
rect 4937 -2967 4969 -2933
rect 5007 -2967 5039 -2933
rect 5039 -2967 5041 -2933
rect 9573 -2606 9607 -2574
rect 9781 -2604 9783 -2570
rect 9783 -2604 9815 -2570
rect 9853 -2604 9885 -2570
rect 9885 -2604 9887 -2570
rect 10233 -2604 10235 -2570
rect 10235 -2604 10267 -2570
rect 10305 -2604 10337 -2570
rect 10337 -2604 10339 -2570
rect 10491 -2604 10493 -2570
rect 10493 -2604 10525 -2570
rect 10563 -2604 10595 -2570
rect 10595 -2604 10597 -2570
rect 10749 -2604 10751 -2570
rect 10751 -2604 10783 -2570
rect 10821 -2604 10853 -2570
rect 10853 -2604 10855 -2570
rect 11007 -2604 11009 -2570
rect 11009 -2604 11041 -2570
rect 11079 -2604 11111 -2570
rect 11111 -2604 11113 -2570
rect 11459 -2604 11461 -2570
rect 11461 -2604 11493 -2570
rect 11531 -2604 11563 -2570
rect 11563 -2604 11565 -2570
rect 11717 -2604 11719 -2570
rect 11719 -2604 11751 -2570
rect 11789 -2604 11821 -2570
rect 11821 -2604 11823 -2570
rect 11975 -2604 11977 -2570
rect 11977 -2604 12009 -2570
rect 12047 -2604 12079 -2570
rect 12079 -2604 12081 -2570
rect 12427 -2604 12429 -2570
rect 12429 -2604 12461 -2570
rect 12499 -2604 12531 -2570
rect 12531 -2604 12533 -2570
rect 12685 -2604 12687 -2570
rect 12687 -2604 12719 -2570
rect 12757 -2604 12789 -2570
rect 12789 -2604 12791 -2570
rect 12943 -2604 12945 -2570
rect 12945 -2604 12977 -2570
rect 13015 -2604 13047 -2570
rect 13047 -2604 13049 -2570
rect 13201 -2604 13203 -2570
rect 13203 -2604 13235 -2570
rect 13273 -2604 13305 -2570
rect 13305 -2604 13307 -2570
rect 13653 -2604 13655 -2570
rect 13655 -2604 13687 -2570
rect 13725 -2604 13757 -2570
rect 13757 -2604 13759 -2570
rect 18290 -2536 18324 -2504
rect 9573 -2608 9607 -2606
rect 9573 -2674 9607 -2646
rect 9573 -2680 9607 -2674
rect 9573 -2742 9607 -2718
rect 9573 -2752 9607 -2742
rect 9573 -2810 9607 -2790
rect 9573 -2824 9607 -2810
rect 9573 -2878 9607 -2862
rect 9573 -2896 9607 -2878
rect 5214 -2946 5248 -2934
rect 856 -3014 890 -3006
rect 5214 -2968 5248 -2946
rect 5421 -2967 5423 -2933
rect 5423 -2967 5455 -2933
rect 5493 -2967 5525 -2933
rect 5525 -2967 5527 -2933
rect 5873 -2967 5875 -2933
rect 5875 -2967 5907 -2933
rect 5945 -2967 5977 -2933
rect 5977 -2967 5979 -2933
rect 6131 -2967 6133 -2933
rect 6133 -2967 6165 -2933
rect 6203 -2967 6235 -2933
rect 6235 -2967 6237 -2933
rect 6389 -2967 6391 -2933
rect 6391 -2967 6423 -2933
rect 6461 -2967 6493 -2933
rect 6493 -2967 6495 -2933
rect 6647 -2967 6649 -2933
rect 6649 -2967 6681 -2933
rect 6719 -2967 6751 -2933
rect 6751 -2967 6753 -2933
rect 7099 -2967 7101 -2933
rect 7101 -2967 7133 -2933
rect 7171 -2967 7203 -2933
rect 7203 -2967 7205 -2933
rect 7357 -2967 7359 -2933
rect 7359 -2967 7391 -2933
rect 7429 -2967 7461 -2933
rect 7461 -2967 7463 -2933
rect 7615 -2967 7617 -2933
rect 7617 -2967 7649 -2933
rect 7687 -2967 7719 -2933
rect 7719 -2967 7721 -2933
rect 8067 -2967 8069 -2933
rect 8069 -2967 8101 -2933
rect 8139 -2967 8171 -2933
rect 8171 -2967 8173 -2933
rect 8325 -2967 8327 -2933
rect 8327 -2967 8359 -2933
rect 8397 -2967 8429 -2933
rect 8429 -2967 8431 -2933
rect 8583 -2967 8585 -2933
rect 8585 -2967 8617 -2933
rect 8655 -2967 8687 -2933
rect 8687 -2967 8689 -2933
rect 8841 -2967 8843 -2933
rect 8843 -2967 8875 -2933
rect 8913 -2967 8945 -2933
rect 8945 -2967 8947 -2933
rect 9293 -2967 9295 -2933
rect 9295 -2967 9327 -2933
rect 9365 -2967 9397 -2933
rect 9397 -2967 9399 -2933
rect 13932 -2606 13966 -2574
rect 14139 -2604 14141 -2570
rect 14141 -2604 14173 -2570
rect 14211 -2604 14243 -2570
rect 14243 -2604 14245 -2570
rect 14590 -2604 14592 -2570
rect 14592 -2604 14624 -2570
rect 14662 -2604 14694 -2570
rect 14694 -2604 14696 -2570
rect 14848 -2604 14850 -2570
rect 14850 -2604 14882 -2570
rect 14920 -2604 14952 -2570
rect 14952 -2604 14954 -2570
rect 15106 -2604 15108 -2570
rect 15108 -2604 15140 -2570
rect 15178 -2604 15210 -2570
rect 15210 -2604 15212 -2570
rect 15364 -2604 15366 -2570
rect 15366 -2604 15398 -2570
rect 15436 -2604 15468 -2570
rect 15468 -2604 15470 -2570
rect 15816 -2604 15818 -2570
rect 15818 -2604 15850 -2570
rect 15888 -2604 15920 -2570
rect 15920 -2604 15922 -2570
rect 16074 -2604 16076 -2570
rect 16076 -2604 16108 -2570
rect 16146 -2604 16178 -2570
rect 16178 -2604 16180 -2570
rect 16332 -2604 16334 -2570
rect 16334 -2604 16366 -2570
rect 16404 -2604 16436 -2570
rect 16436 -2604 16438 -2570
rect 16784 -2604 16786 -2570
rect 16786 -2604 16818 -2570
rect 16856 -2604 16888 -2570
rect 16888 -2604 16890 -2570
rect 17042 -2604 17044 -2570
rect 17044 -2604 17076 -2570
rect 17114 -2604 17146 -2570
rect 17146 -2604 17148 -2570
rect 17300 -2604 17302 -2570
rect 17302 -2604 17334 -2570
rect 17372 -2604 17404 -2570
rect 17404 -2604 17406 -2570
rect 17558 -2604 17560 -2570
rect 17560 -2604 17592 -2570
rect 17630 -2604 17662 -2570
rect 17662 -2604 17664 -2570
rect 18010 -2604 18012 -2570
rect 18012 -2604 18044 -2570
rect 18082 -2604 18114 -2570
rect 18114 -2604 18116 -2570
rect 13932 -2608 13966 -2606
rect 13932 -2674 13966 -2646
rect 13932 -2680 13966 -2674
rect 13932 -2742 13966 -2718
rect 13932 -2752 13966 -2742
rect 13932 -2810 13966 -2790
rect 13932 -2824 13966 -2810
rect 13932 -2878 13966 -2862
rect 13932 -2896 13966 -2878
rect 9573 -2946 9607 -2934
rect 856 -3040 890 -3014
rect 856 -3082 890 -3078
rect 856 -3112 890 -3082
rect 856 -3184 890 -3150
rect 971 -3063 1005 -3061
rect 971 -3095 1005 -3063
rect 971 -3165 1005 -3133
rect 971 -3167 1005 -3165
rect 1229 -3063 1263 -3061
rect 1229 -3095 1263 -3063
rect 1229 -3165 1263 -3133
rect 1229 -3167 1263 -3165
rect 1423 -3063 1457 -3061
rect 1423 -3095 1457 -3063
rect 1423 -3165 1457 -3133
rect 1423 -3167 1457 -3165
rect 1681 -3063 1715 -3061
rect 1681 -3095 1715 -3063
rect 1681 -3165 1715 -3133
rect 1681 -3167 1715 -3165
rect 1939 -3063 1973 -3061
rect 1939 -3095 1973 -3063
rect 1939 -3165 1973 -3133
rect 1939 -3167 1973 -3165
rect 2197 -3063 2231 -3061
rect 2197 -3095 2231 -3063
rect 2197 -3165 2231 -3133
rect 2197 -3167 2231 -3165
rect 2455 -3063 2489 -3061
rect 2455 -3095 2489 -3063
rect 2455 -3165 2489 -3133
rect 2455 -3167 2489 -3165
rect 2649 -3063 2683 -3061
rect 2649 -3095 2683 -3063
rect 2649 -3165 2683 -3133
rect 2649 -3167 2683 -3165
rect 2907 -3063 2941 -3061
rect 2907 -3095 2941 -3063
rect 2907 -3165 2941 -3133
rect 2907 -3167 2941 -3165
rect 3165 -3063 3199 -3061
rect 3165 -3095 3199 -3063
rect 3165 -3165 3199 -3133
rect 3165 -3167 3199 -3165
rect 3423 -3063 3457 -3061
rect 3423 -3095 3457 -3063
rect 3423 -3165 3457 -3133
rect 3423 -3167 3457 -3165
rect 3617 -3063 3651 -3061
rect 3617 -3095 3651 -3063
rect 3617 -3165 3651 -3133
rect 3617 -3167 3651 -3165
rect 3875 -3063 3909 -3061
rect 3875 -3095 3909 -3063
rect 3875 -3165 3909 -3133
rect 3875 -3167 3909 -3165
rect 4133 -3063 4167 -3061
rect 4133 -3095 4167 -3063
rect 4133 -3165 4167 -3133
rect 4133 -3167 4167 -3165
rect 4391 -3063 4425 -3061
rect 4391 -3095 4425 -3063
rect 4391 -3165 4425 -3133
rect 4391 -3167 4425 -3165
rect 4649 -3063 4683 -3061
rect 4649 -3095 4683 -3063
rect 4649 -3165 4683 -3133
rect 4649 -3167 4683 -3165
rect 4842 -3063 4876 -3061
rect 4842 -3095 4876 -3063
rect 4842 -3165 4876 -3133
rect 4842 -3167 4876 -3165
rect 5100 -3063 5134 -3061
rect 5100 -3095 5134 -3063
rect 5100 -3165 5134 -3133
rect 5100 -3167 5134 -3165
rect 5214 -3014 5248 -3006
rect 5214 -3040 5248 -3014
rect 9573 -2968 9607 -2946
rect 9781 -2967 9783 -2933
rect 9783 -2967 9815 -2933
rect 9853 -2967 9885 -2933
rect 9885 -2967 9887 -2933
rect 10233 -2967 10235 -2933
rect 10235 -2967 10267 -2933
rect 10305 -2967 10337 -2933
rect 10337 -2967 10339 -2933
rect 10491 -2967 10493 -2933
rect 10493 -2967 10525 -2933
rect 10563 -2967 10595 -2933
rect 10595 -2967 10597 -2933
rect 10749 -2967 10751 -2933
rect 10751 -2967 10783 -2933
rect 10821 -2967 10853 -2933
rect 10853 -2967 10855 -2933
rect 11007 -2967 11009 -2933
rect 11009 -2967 11041 -2933
rect 11079 -2967 11111 -2933
rect 11111 -2967 11113 -2933
rect 11459 -2967 11461 -2933
rect 11461 -2967 11493 -2933
rect 11531 -2967 11563 -2933
rect 11563 -2967 11565 -2933
rect 11717 -2967 11719 -2933
rect 11719 -2967 11751 -2933
rect 11789 -2967 11821 -2933
rect 11821 -2967 11823 -2933
rect 11975 -2967 11977 -2933
rect 11977 -2967 12009 -2933
rect 12047 -2967 12079 -2933
rect 12079 -2967 12081 -2933
rect 12427 -2967 12429 -2933
rect 12429 -2967 12461 -2933
rect 12499 -2967 12531 -2933
rect 12531 -2967 12533 -2933
rect 12685 -2967 12687 -2933
rect 12687 -2967 12719 -2933
rect 12757 -2967 12789 -2933
rect 12789 -2967 12791 -2933
rect 12943 -2967 12945 -2933
rect 12945 -2967 12977 -2933
rect 13015 -2967 13047 -2933
rect 13047 -2967 13049 -2933
rect 13201 -2967 13203 -2933
rect 13203 -2967 13235 -2933
rect 13273 -2967 13305 -2933
rect 13305 -2967 13307 -2933
rect 13653 -2967 13655 -2933
rect 13655 -2967 13687 -2933
rect 13725 -2967 13757 -2933
rect 13757 -2967 13759 -2933
rect 18290 -2606 18324 -2574
rect 18290 -2608 18324 -2606
rect 18290 -2674 18324 -2646
rect 18290 -2680 18324 -2674
rect 18290 -2742 18324 -2718
rect 18290 -2752 18324 -2742
rect 18290 -2810 18324 -2790
rect 18290 -2824 18324 -2810
rect 18290 -2878 18324 -2862
rect 18290 -2896 18324 -2878
rect 5214 -3082 5248 -3078
rect 5214 -3112 5248 -3082
rect 5214 -3184 5248 -3150
rect 5328 -3063 5362 -3061
rect 5328 -3095 5362 -3063
rect 5328 -3165 5362 -3133
rect 5328 -3167 5362 -3165
rect 5586 -3063 5620 -3061
rect 5586 -3095 5620 -3063
rect 5586 -3165 5620 -3133
rect 5586 -3167 5620 -3165
rect 5780 -3063 5814 -3061
rect 5780 -3095 5814 -3063
rect 5780 -3165 5814 -3133
rect 5780 -3167 5814 -3165
rect 6038 -3063 6072 -3061
rect 6038 -3095 6072 -3063
rect 6038 -3165 6072 -3133
rect 6038 -3167 6072 -3165
rect 6296 -3063 6330 -3061
rect 6296 -3095 6330 -3063
rect 6296 -3165 6330 -3133
rect 6296 -3167 6330 -3165
rect 6554 -3063 6588 -3061
rect 6554 -3095 6588 -3063
rect 6554 -3165 6588 -3133
rect 6554 -3167 6588 -3165
rect 6812 -3063 6846 -3061
rect 6812 -3095 6846 -3063
rect 6812 -3165 6846 -3133
rect 6812 -3167 6846 -3165
rect 7006 -3063 7040 -3061
rect 7006 -3095 7040 -3063
rect 7006 -3165 7040 -3133
rect 7006 -3167 7040 -3165
rect 7264 -3063 7298 -3061
rect 7264 -3095 7298 -3063
rect 7264 -3165 7298 -3133
rect 7264 -3167 7298 -3165
rect 7522 -3063 7556 -3061
rect 7522 -3095 7556 -3063
rect 7522 -3165 7556 -3133
rect 7522 -3167 7556 -3165
rect 7780 -3063 7814 -3061
rect 7780 -3095 7814 -3063
rect 7780 -3165 7814 -3133
rect 7780 -3167 7814 -3165
rect 7974 -3063 8008 -3061
rect 7974 -3095 8008 -3063
rect 7974 -3165 8008 -3133
rect 7974 -3167 8008 -3165
rect 8232 -3063 8266 -3061
rect 8232 -3095 8266 -3063
rect 8232 -3165 8266 -3133
rect 8232 -3167 8266 -3165
rect 8490 -3063 8524 -3061
rect 8490 -3095 8524 -3063
rect 8490 -3165 8524 -3133
rect 8490 -3167 8524 -3165
rect 8748 -3063 8782 -3061
rect 8748 -3095 8782 -3063
rect 8748 -3165 8782 -3133
rect 8748 -3167 8782 -3165
rect 9006 -3063 9040 -3061
rect 9006 -3095 9040 -3063
rect 9006 -3165 9040 -3133
rect 9006 -3167 9040 -3165
rect 9200 -3063 9234 -3061
rect 9200 -3095 9234 -3063
rect 9200 -3165 9234 -3133
rect 9200 -3167 9234 -3165
rect 9458 -3063 9492 -3061
rect 9458 -3095 9492 -3063
rect 9458 -3165 9492 -3133
rect 9458 -3167 9492 -3165
rect 9573 -3014 9607 -3006
rect 13932 -2946 13966 -2934
rect 13932 -2968 13966 -2946
rect 14139 -2967 14141 -2933
rect 14141 -2967 14173 -2933
rect 14211 -2967 14243 -2933
rect 14243 -2967 14245 -2933
rect 14590 -2967 14592 -2933
rect 14592 -2967 14624 -2933
rect 14662 -2967 14694 -2933
rect 14694 -2967 14696 -2933
rect 14848 -2967 14850 -2933
rect 14850 -2967 14882 -2933
rect 14920 -2967 14952 -2933
rect 14952 -2967 14954 -2933
rect 15106 -2967 15108 -2933
rect 15108 -2967 15140 -2933
rect 15178 -2967 15210 -2933
rect 15210 -2967 15212 -2933
rect 15364 -2967 15366 -2933
rect 15366 -2967 15398 -2933
rect 15436 -2967 15468 -2933
rect 15468 -2967 15470 -2933
rect 15816 -2967 15818 -2933
rect 15818 -2967 15850 -2933
rect 15888 -2967 15920 -2933
rect 15920 -2967 15922 -2933
rect 16074 -2967 16076 -2933
rect 16076 -2967 16108 -2933
rect 16146 -2967 16178 -2933
rect 16178 -2967 16180 -2933
rect 16332 -2967 16334 -2933
rect 16334 -2967 16366 -2933
rect 16404 -2967 16436 -2933
rect 16436 -2967 16438 -2933
rect 16784 -2967 16786 -2933
rect 16786 -2967 16818 -2933
rect 16856 -2967 16888 -2933
rect 16888 -2967 16890 -2933
rect 17042 -2967 17044 -2933
rect 17044 -2967 17076 -2933
rect 17114 -2967 17146 -2933
rect 17146 -2967 17148 -2933
rect 17300 -2967 17302 -2933
rect 17302 -2967 17334 -2933
rect 17372 -2967 17404 -2933
rect 17404 -2967 17406 -2933
rect 17558 -2967 17560 -2933
rect 17560 -2967 17592 -2933
rect 17630 -2967 17662 -2933
rect 17662 -2967 17664 -2933
rect 18010 -2967 18012 -2933
rect 18012 -2967 18044 -2933
rect 18082 -2967 18114 -2933
rect 18114 -2967 18116 -2933
rect 18290 -2946 18324 -2934
rect 9573 -3040 9607 -3014
rect 9573 -3082 9607 -3078
rect 9573 -3112 9607 -3082
rect 9573 -3184 9607 -3150
rect 9688 -3063 9722 -3061
rect 9688 -3095 9722 -3063
rect 9688 -3165 9722 -3133
rect 9688 -3167 9722 -3165
rect 9946 -3063 9980 -3061
rect 9946 -3095 9980 -3063
rect 9946 -3165 9980 -3133
rect 9946 -3167 9980 -3165
rect 10140 -3063 10174 -3061
rect 10140 -3095 10174 -3063
rect 10140 -3165 10174 -3133
rect 10140 -3167 10174 -3165
rect 10398 -3063 10432 -3061
rect 10398 -3095 10432 -3063
rect 10398 -3165 10432 -3133
rect 10398 -3167 10432 -3165
rect 10656 -3063 10690 -3061
rect 10656 -3095 10690 -3063
rect 10656 -3165 10690 -3133
rect 10656 -3167 10690 -3165
rect 10914 -3063 10948 -3061
rect 10914 -3095 10948 -3063
rect 10914 -3165 10948 -3133
rect 10914 -3167 10948 -3165
rect 11172 -3063 11206 -3061
rect 11172 -3095 11206 -3063
rect 11172 -3165 11206 -3133
rect 11172 -3167 11206 -3165
rect 11366 -3063 11400 -3061
rect 11366 -3095 11400 -3063
rect 11366 -3165 11400 -3133
rect 11366 -3167 11400 -3165
rect 11624 -3063 11658 -3061
rect 11624 -3095 11658 -3063
rect 11624 -3165 11658 -3133
rect 11624 -3167 11658 -3165
rect 11882 -3063 11916 -3061
rect 11882 -3095 11916 -3063
rect 11882 -3165 11916 -3133
rect 11882 -3167 11916 -3165
rect 12140 -3063 12174 -3061
rect 12140 -3095 12174 -3063
rect 12140 -3165 12174 -3133
rect 12140 -3167 12174 -3165
rect 12334 -3063 12368 -3061
rect 12334 -3095 12368 -3063
rect 12334 -3165 12368 -3133
rect 12334 -3167 12368 -3165
rect 12592 -3063 12626 -3061
rect 12592 -3095 12626 -3063
rect 12592 -3165 12626 -3133
rect 12592 -3167 12626 -3165
rect 12850 -3063 12884 -3061
rect 12850 -3095 12884 -3063
rect 12850 -3165 12884 -3133
rect 12850 -3167 12884 -3165
rect 13108 -3063 13142 -3061
rect 13108 -3095 13142 -3063
rect 13108 -3165 13142 -3133
rect 13108 -3167 13142 -3165
rect 13366 -3063 13400 -3061
rect 13366 -3095 13400 -3063
rect 13366 -3165 13400 -3133
rect 13366 -3167 13400 -3165
rect 13560 -3063 13594 -3061
rect 13560 -3095 13594 -3063
rect 13560 -3165 13594 -3133
rect 13560 -3167 13594 -3165
rect 13818 -3063 13852 -3061
rect 13818 -3095 13852 -3063
rect 13818 -3165 13852 -3133
rect 13818 -3167 13852 -3165
rect 13932 -3014 13966 -3006
rect 18290 -2968 18324 -2946
rect 13932 -3040 13966 -3014
rect 13932 -3082 13966 -3078
rect 13932 -3112 13966 -3082
rect 13932 -3184 13966 -3150
rect 14046 -3063 14080 -3061
rect 14046 -3095 14080 -3063
rect 14046 -3165 14080 -3133
rect 14046 -3167 14080 -3165
rect 14304 -3063 14338 -3061
rect 14304 -3095 14338 -3063
rect 14304 -3165 14338 -3133
rect 14304 -3167 14338 -3165
rect 14497 -3063 14531 -3061
rect 14497 -3095 14531 -3063
rect 14497 -3165 14531 -3133
rect 14497 -3167 14531 -3165
rect 14755 -3063 14789 -3061
rect 14755 -3095 14789 -3063
rect 14755 -3165 14789 -3133
rect 14755 -3167 14789 -3165
rect 15013 -3063 15047 -3061
rect 15013 -3095 15047 -3063
rect 15013 -3165 15047 -3133
rect 15013 -3167 15047 -3165
rect 15271 -3063 15305 -3061
rect 15271 -3095 15305 -3063
rect 15271 -3165 15305 -3133
rect 15271 -3167 15305 -3165
rect 15529 -3063 15563 -3061
rect 15529 -3095 15563 -3063
rect 15529 -3165 15563 -3133
rect 15529 -3167 15563 -3165
rect 15723 -3063 15757 -3061
rect 15723 -3095 15757 -3063
rect 15723 -3165 15757 -3133
rect 15723 -3167 15757 -3165
rect 15981 -3063 16015 -3061
rect 15981 -3095 16015 -3063
rect 15981 -3165 16015 -3133
rect 15981 -3167 16015 -3165
rect 16239 -3063 16273 -3061
rect 16239 -3095 16273 -3063
rect 16239 -3165 16273 -3133
rect 16239 -3167 16273 -3165
rect 16497 -3063 16531 -3061
rect 16497 -3095 16531 -3063
rect 16497 -3165 16531 -3133
rect 16497 -3167 16531 -3165
rect 16691 -3063 16725 -3061
rect 16691 -3095 16725 -3063
rect 16691 -3165 16725 -3133
rect 16691 -3167 16725 -3165
rect 16949 -3063 16983 -3061
rect 16949 -3095 16983 -3063
rect 16949 -3165 16983 -3133
rect 16949 -3167 16983 -3165
rect 17207 -3063 17241 -3061
rect 17207 -3095 17241 -3063
rect 17207 -3165 17241 -3133
rect 17207 -3167 17241 -3165
rect 17465 -3063 17499 -3061
rect 17465 -3095 17499 -3063
rect 17465 -3165 17499 -3133
rect 17465 -3167 17499 -3165
rect 17723 -3063 17757 -3061
rect 17723 -3095 17757 -3063
rect 17723 -3165 17757 -3133
rect 17723 -3167 17757 -3165
rect 17917 -3063 17951 -3061
rect 17917 -3095 17951 -3063
rect 17917 -3165 17951 -3133
rect 17917 -3167 17951 -3165
rect 18175 -3063 18209 -3061
rect 18175 -3095 18209 -3063
rect 18175 -3165 18209 -3133
rect 18175 -3167 18209 -3165
rect 18290 -3014 18324 -3006
rect 18290 -3040 18324 -3014
rect 18290 -3082 18324 -3078
rect 18290 -3112 18324 -3082
rect 18290 -3184 18324 -3150
rect 856 -3252 890 -3222
rect 856 -3256 890 -3252
rect 856 -3320 890 -3294
rect 856 -3328 890 -3320
rect 856 -3388 890 -3366
rect 856 -3400 890 -3388
rect 856 -3456 890 -3438
rect 856 -3472 890 -3456
rect 856 -3524 890 -3510
rect 856 -3544 890 -3524
rect 856 -3592 890 -3582
rect 5214 -3252 5248 -3222
rect 5214 -3256 5248 -3252
rect 5214 -3320 5248 -3294
rect 5214 -3328 5248 -3320
rect 5214 -3388 5248 -3366
rect 5214 -3400 5248 -3388
rect 5214 -3456 5248 -3438
rect 5214 -3472 5248 -3456
rect 5214 -3524 5248 -3510
rect 5214 -3544 5248 -3524
rect 5214 -3592 5248 -3582
rect 9573 -3252 9607 -3222
rect 9573 -3256 9607 -3252
rect 9573 -3320 9607 -3294
rect 9573 -3328 9607 -3320
rect 9573 -3388 9607 -3366
rect 9573 -3400 9607 -3388
rect 9573 -3456 9607 -3438
rect 9573 -3472 9607 -3456
rect 9573 -3524 9607 -3510
rect 9573 -3544 9607 -3524
rect 9573 -3592 9607 -3582
rect 13932 -3252 13966 -3222
rect 13932 -3256 13966 -3252
rect 13932 -3320 13966 -3294
rect 13932 -3328 13966 -3320
rect 13932 -3388 13966 -3366
rect 13932 -3400 13966 -3388
rect 13932 -3456 13966 -3438
rect 13932 -3472 13966 -3456
rect 13932 -3524 13966 -3510
rect 13932 -3544 13966 -3524
rect 13932 -3592 13966 -3582
rect 18290 -3252 18324 -3222
rect 18290 -3256 18324 -3252
rect 18290 -3320 18324 -3294
rect 18290 -3328 18324 -3320
rect 18290 -3388 18324 -3366
rect 18290 -3400 18324 -3388
rect 18290 -3456 18324 -3438
rect 18290 -3472 18324 -3456
rect 18290 -3524 18324 -3510
rect 18290 -3544 18324 -3524
rect 18290 -3592 18324 -3582
rect 856 -3616 890 -3592
rect 5214 -3616 5248 -3592
rect 9573 -3616 9607 -3592
rect 13932 -3616 13966 -3592
rect 18290 -3616 18324 -3592
rect 856 -3660 890 -3654
rect 856 -3688 890 -3660
rect 856 -3728 890 -3726
rect 856 -3760 890 -3728
rect 856 -3830 890 -3798
rect 856 -3832 890 -3830
rect 856 -3898 890 -3870
rect 856 -3904 890 -3898
rect 856 -3966 890 -3942
rect 856 -3976 890 -3966
rect 5214 -3660 5248 -3654
rect 5214 -3688 5248 -3660
rect 5214 -3728 5248 -3726
rect 5214 -3760 5248 -3728
rect 5214 -3830 5248 -3798
rect 5214 -3832 5248 -3830
rect 5214 -3898 5248 -3870
rect 5214 -3904 5248 -3898
rect 5214 -3966 5248 -3942
rect 5214 -3976 5248 -3966
rect 9573 -3660 9607 -3654
rect 9573 -3688 9607 -3660
rect 9573 -3728 9607 -3726
rect 9573 -3760 9607 -3728
rect 9573 -3830 9607 -3798
rect 9573 -3832 9607 -3830
rect 9573 -3898 9607 -3870
rect 9573 -3904 9607 -3898
rect 9573 -3966 9607 -3942
rect 9573 -3976 9607 -3966
rect 13932 -3660 13966 -3654
rect 13932 -3688 13966 -3660
rect 13932 -3728 13966 -3726
rect 13932 -3760 13966 -3728
rect 13932 -3830 13966 -3798
rect 13932 -3832 13966 -3830
rect 13932 -3898 13966 -3870
rect 13932 -3904 13966 -3898
rect 13932 -3966 13966 -3942
rect 13932 -3976 13966 -3966
rect 18290 -3660 18324 -3654
rect 18290 -3688 18324 -3660
rect 18290 -3728 18324 -3726
rect 18290 -3760 18324 -3728
rect 18290 -3830 18324 -3798
rect 18290 -3832 18324 -3830
rect 18290 -3898 18324 -3870
rect 18290 -3904 18324 -3898
rect 18290 -3966 18324 -3942
rect 18290 -3976 18324 -3966
rect 856 -4034 890 -4014
rect 856 -4048 890 -4034
rect 856 -4102 890 -4086
rect 856 -4120 890 -4102
rect 856 -4192 890 -4158
rect 971 -4053 1005 -4051
rect 971 -4085 1005 -4053
rect 971 -4155 1005 -4123
rect 971 -4157 1005 -4155
rect 1229 -4053 1263 -4051
rect 1229 -4085 1263 -4053
rect 1229 -4155 1263 -4123
rect 1229 -4157 1263 -4155
rect 1423 -4053 1457 -4051
rect 1423 -4085 1457 -4053
rect 1423 -4155 1457 -4123
rect 1423 -4157 1457 -4155
rect 1681 -4053 1715 -4051
rect 1681 -4085 1715 -4053
rect 1681 -4155 1715 -4123
rect 1681 -4157 1715 -4155
rect 1939 -4053 1973 -4051
rect 1939 -4085 1973 -4053
rect 1939 -4155 1973 -4123
rect 1939 -4157 1973 -4155
rect 2197 -4053 2231 -4051
rect 2197 -4085 2231 -4053
rect 2197 -4155 2231 -4123
rect 2197 -4157 2231 -4155
rect 2455 -4053 2489 -4051
rect 2455 -4085 2489 -4053
rect 2455 -4155 2489 -4123
rect 2455 -4157 2489 -4155
rect 2649 -4053 2683 -4051
rect 2649 -4085 2683 -4053
rect 2649 -4155 2683 -4123
rect 2649 -4157 2683 -4155
rect 2907 -4053 2941 -4051
rect 2907 -4085 2941 -4053
rect 2907 -4155 2941 -4123
rect 2907 -4157 2941 -4155
rect 3165 -4053 3199 -4051
rect 3165 -4085 3199 -4053
rect 3165 -4155 3199 -4123
rect 3165 -4157 3199 -4155
rect 3423 -4053 3457 -4051
rect 3423 -4085 3457 -4053
rect 3423 -4155 3457 -4123
rect 3423 -4157 3457 -4155
rect 3617 -4053 3651 -4051
rect 3617 -4085 3651 -4053
rect 3617 -4155 3651 -4123
rect 3617 -4157 3651 -4155
rect 3875 -4053 3909 -4051
rect 3875 -4085 3909 -4053
rect 3875 -4155 3909 -4123
rect 3875 -4157 3909 -4155
rect 4133 -4053 4167 -4051
rect 4133 -4085 4167 -4053
rect 4133 -4155 4167 -4123
rect 4133 -4157 4167 -4155
rect 4391 -4053 4425 -4051
rect 4391 -4085 4425 -4053
rect 4391 -4155 4425 -4123
rect 4391 -4157 4425 -4155
rect 4649 -4053 4683 -4051
rect 4649 -4085 4683 -4053
rect 4649 -4155 4683 -4123
rect 4649 -4157 4683 -4155
rect 4842 -4053 4876 -4051
rect 4842 -4085 4876 -4053
rect 4842 -4155 4876 -4123
rect 4842 -4157 4876 -4155
rect 5100 -4053 5134 -4051
rect 5100 -4085 5134 -4053
rect 5100 -4155 5134 -4123
rect 5100 -4157 5134 -4155
rect 5214 -4034 5248 -4014
rect 5214 -4048 5248 -4034
rect 5214 -4102 5248 -4086
rect 5214 -4120 5248 -4102
rect 5214 -4192 5248 -4158
rect 856 -4264 890 -4230
rect 5328 -4053 5362 -4051
rect 5328 -4085 5362 -4053
rect 5328 -4155 5362 -4123
rect 5328 -4157 5362 -4155
rect 5586 -4053 5620 -4051
rect 5586 -4085 5620 -4053
rect 5586 -4155 5620 -4123
rect 5586 -4157 5620 -4155
rect 5780 -4053 5814 -4051
rect 5780 -4085 5814 -4053
rect 5780 -4155 5814 -4123
rect 5780 -4157 5814 -4155
rect 6038 -4053 6072 -4051
rect 6038 -4085 6072 -4053
rect 6038 -4155 6072 -4123
rect 6038 -4157 6072 -4155
rect 6296 -4053 6330 -4051
rect 6296 -4085 6330 -4053
rect 6296 -4155 6330 -4123
rect 6296 -4157 6330 -4155
rect 6554 -4053 6588 -4051
rect 6554 -4085 6588 -4053
rect 6554 -4155 6588 -4123
rect 6554 -4157 6588 -4155
rect 6812 -4053 6846 -4051
rect 6812 -4085 6846 -4053
rect 6812 -4155 6846 -4123
rect 6812 -4157 6846 -4155
rect 7006 -4053 7040 -4051
rect 7006 -4085 7040 -4053
rect 7006 -4155 7040 -4123
rect 7006 -4157 7040 -4155
rect 7264 -4053 7298 -4051
rect 7264 -4085 7298 -4053
rect 7264 -4155 7298 -4123
rect 7264 -4157 7298 -4155
rect 7522 -4053 7556 -4051
rect 7522 -4085 7556 -4053
rect 7522 -4155 7556 -4123
rect 7522 -4157 7556 -4155
rect 7780 -4053 7814 -4051
rect 7780 -4085 7814 -4053
rect 7780 -4155 7814 -4123
rect 7780 -4157 7814 -4155
rect 7974 -4053 8008 -4051
rect 7974 -4085 8008 -4053
rect 7974 -4155 8008 -4123
rect 7974 -4157 8008 -4155
rect 8232 -4053 8266 -4051
rect 8232 -4085 8266 -4053
rect 8232 -4155 8266 -4123
rect 8232 -4157 8266 -4155
rect 8490 -4053 8524 -4051
rect 8490 -4085 8524 -4053
rect 8490 -4155 8524 -4123
rect 8490 -4157 8524 -4155
rect 8748 -4053 8782 -4051
rect 8748 -4085 8782 -4053
rect 8748 -4155 8782 -4123
rect 8748 -4157 8782 -4155
rect 9006 -4053 9040 -4051
rect 9006 -4085 9040 -4053
rect 9006 -4155 9040 -4123
rect 9006 -4157 9040 -4155
rect 9200 -4053 9234 -4051
rect 9200 -4085 9234 -4053
rect 9200 -4155 9234 -4123
rect 9200 -4157 9234 -4155
rect 9458 -4053 9492 -4051
rect 9458 -4085 9492 -4053
rect 9458 -4155 9492 -4123
rect 9458 -4157 9492 -4155
rect 9573 -4034 9607 -4014
rect 9573 -4048 9607 -4034
rect 9573 -4102 9607 -4086
rect 9573 -4120 9607 -4102
rect 9573 -4192 9607 -4158
rect 1064 -4285 1066 -4251
rect 1066 -4285 1098 -4251
rect 1136 -4285 1168 -4251
rect 1168 -4285 1170 -4251
rect 1516 -4285 1518 -4251
rect 1518 -4285 1550 -4251
rect 1588 -4285 1620 -4251
rect 1620 -4285 1622 -4251
rect 1774 -4285 1776 -4251
rect 1776 -4285 1808 -4251
rect 1846 -4285 1878 -4251
rect 1878 -4285 1880 -4251
rect 2032 -4285 2034 -4251
rect 2034 -4285 2066 -4251
rect 2104 -4285 2136 -4251
rect 2136 -4285 2138 -4251
rect 2290 -4285 2292 -4251
rect 2292 -4285 2324 -4251
rect 2362 -4285 2394 -4251
rect 2394 -4285 2396 -4251
rect 2742 -4285 2744 -4251
rect 2744 -4285 2776 -4251
rect 2814 -4285 2846 -4251
rect 2846 -4285 2848 -4251
rect 3000 -4285 3002 -4251
rect 3002 -4285 3034 -4251
rect 3072 -4285 3104 -4251
rect 3104 -4285 3106 -4251
rect 3258 -4285 3260 -4251
rect 3260 -4285 3292 -4251
rect 3330 -4285 3362 -4251
rect 3362 -4285 3364 -4251
rect 3710 -4285 3712 -4251
rect 3712 -4285 3744 -4251
rect 3782 -4285 3814 -4251
rect 3814 -4285 3816 -4251
rect 3968 -4285 3970 -4251
rect 3970 -4285 4002 -4251
rect 4040 -4285 4072 -4251
rect 4072 -4285 4074 -4251
rect 4226 -4285 4228 -4251
rect 4228 -4285 4260 -4251
rect 4298 -4285 4330 -4251
rect 4330 -4285 4332 -4251
rect 4484 -4285 4486 -4251
rect 4486 -4285 4518 -4251
rect 4556 -4285 4588 -4251
rect 4588 -4285 4590 -4251
rect 4935 -4285 4937 -4251
rect 4937 -4285 4969 -4251
rect 5007 -4285 5039 -4251
rect 5039 -4285 5041 -4251
rect 5214 -4264 5248 -4230
rect 9688 -4053 9722 -4051
rect 9688 -4085 9722 -4053
rect 9688 -4155 9722 -4123
rect 9688 -4157 9722 -4155
rect 9946 -4053 9980 -4051
rect 9946 -4085 9980 -4053
rect 9946 -4155 9980 -4123
rect 9946 -4157 9980 -4155
rect 10140 -4053 10174 -4051
rect 10140 -4085 10174 -4053
rect 10140 -4155 10174 -4123
rect 10140 -4157 10174 -4155
rect 10398 -4053 10432 -4051
rect 10398 -4085 10432 -4053
rect 10398 -4155 10432 -4123
rect 10398 -4157 10432 -4155
rect 10656 -4053 10690 -4051
rect 10656 -4085 10690 -4053
rect 10656 -4155 10690 -4123
rect 10656 -4157 10690 -4155
rect 10914 -4053 10948 -4051
rect 10914 -4085 10948 -4053
rect 10914 -4155 10948 -4123
rect 10914 -4157 10948 -4155
rect 11172 -4053 11206 -4051
rect 11172 -4085 11206 -4053
rect 11172 -4155 11206 -4123
rect 11172 -4157 11206 -4155
rect 11366 -4053 11400 -4051
rect 11366 -4085 11400 -4053
rect 11366 -4155 11400 -4123
rect 11366 -4157 11400 -4155
rect 11624 -4053 11658 -4051
rect 11624 -4085 11658 -4053
rect 11624 -4155 11658 -4123
rect 11624 -4157 11658 -4155
rect 11882 -4053 11916 -4051
rect 11882 -4085 11916 -4053
rect 11882 -4155 11916 -4123
rect 11882 -4157 11916 -4155
rect 12140 -4053 12174 -4051
rect 12140 -4085 12174 -4053
rect 12140 -4155 12174 -4123
rect 12140 -4157 12174 -4155
rect 12334 -4053 12368 -4051
rect 12334 -4085 12368 -4053
rect 12334 -4155 12368 -4123
rect 12334 -4157 12368 -4155
rect 12592 -4053 12626 -4051
rect 12592 -4085 12626 -4053
rect 12592 -4155 12626 -4123
rect 12592 -4157 12626 -4155
rect 12850 -4053 12884 -4051
rect 12850 -4085 12884 -4053
rect 12850 -4155 12884 -4123
rect 12850 -4157 12884 -4155
rect 13108 -4053 13142 -4051
rect 13108 -4085 13142 -4053
rect 13108 -4155 13142 -4123
rect 13108 -4157 13142 -4155
rect 13366 -4053 13400 -4051
rect 13366 -4085 13400 -4053
rect 13366 -4155 13400 -4123
rect 13366 -4157 13400 -4155
rect 13560 -4053 13594 -4051
rect 13560 -4085 13594 -4053
rect 13560 -4155 13594 -4123
rect 13560 -4157 13594 -4155
rect 13818 -4053 13852 -4051
rect 13818 -4085 13852 -4053
rect 13818 -4155 13852 -4123
rect 13818 -4157 13852 -4155
rect 13932 -4034 13966 -4014
rect 13932 -4048 13966 -4034
rect 13932 -4102 13966 -4086
rect 13932 -4120 13966 -4102
rect 13932 -4192 13966 -4158
rect 856 -4336 890 -4302
rect 5421 -4285 5423 -4251
rect 5423 -4285 5455 -4251
rect 5493 -4285 5525 -4251
rect 5525 -4285 5527 -4251
rect 5873 -4285 5875 -4251
rect 5875 -4285 5907 -4251
rect 5945 -4285 5977 -4251
rect 5977 -4285 5979 -4251
rect 6131 -4285 6133 -4251
rect 6133 -4285 6165 -4251
rect 6203 -4285 6235 -4251
rect 6235 -4285 6237 -4251
rect 6389 -4285 6391 -4251
rect 6391 -4285 6423 -4251
rect 6461 -4285 6493 -4251
rect 6493 -4285 6495 -4251
rect 6647 -4285 6649 -4251
rect 6649 -4285 6681 -4251
rect 6719 -4285 6751 -4251
rect 6751 -4285 6753 -4251
rect 7099 -4285 7101 -4251
rect 7101 -4285 7133 -4251
rect 7171 -4285 7203 -4251
rect 7203 -4285 7205 -4251
rect 7357 -4285 7359 -4251
rect 7359 -4285 7391 -4251
rect 7429 -4285 7461 -4251
rect 7461 -4285 7463 -4251
rect 7615 -4285 7617 -4251
rect 7617 -4285 7649 -4251
rect 7687 -4285 7719 -4251
rect 7719 -4285 7721 -4251
rect 8067 -4285 8069 -4251
rect 8069 -4285 8101 -4251
rect 8139 -4285 8171 -4251
rect 8171 -4285 8173 -4251
rect 8325 -4285 8327 -4251
rect 8327 -4285 8359 -4251
rect 8397 -4285 8429 -4251
rect 8429 -4285 8431 -4251
rect 8583 -4285 8585 -4251
rect 8585 -4285 8617 -4251
rect 8655 -4285 8687 -4251
rect 8687 -4285 8689 -4251
rect 8841 -4285 8843 -4251
rect 8843 -4285 8875 -4251
rect 8913 -4285 8945 -4251
rect 8945 -4285 8947 -4251
rect 9293 -4285 9295 -4251
rect 9295 -4285 9327 -4251
rect 9365 -4285 9397 -4251
rect 9397 -4285 9399 -4251
rect 9573 -4264 9607 -4230
rect 14046 -4053 14080 -4051
rect 14046 -4085 14080 -4053
rect 14046 -4155 14080 -4123
rect 14046 -4157 14080 -4155
rect 14304 -4053 14338 -4051
rect 14304 -4085 14338 -4053
rect 14304 -4155 14338 -4123
rect 14304 -4157 14338 -4155
rect 14497 -4053 14531 -4051
rect 14497 -4085 14531 -4053
rect 14497 -4155 14531 -4123
rect 14497 -4157 14531 -4155
rect 14755 -4053 14789 -4051
rect 14755 -4085 14789 -4053
rect 14755 -4155 14789 -4123
rect 14755 -4157 14789 -4155
rect 15013 -4053 15047 -4051
rect 15013 -4085 15047 -4053
rect 15013 -4155 15047 -4123
rect 15013 -4157 15047 -4155
rect 15271 -4053 15305 -4051
rect 15271 -4085 15305 -4053
rect 15271 -4155 15305 -4123
rect 15271 -4157 15305 -4155
rect 15529 -4053 15563 -4051
rect 15529 -4085 15563 -4053
rect 15529 -4155 15563 -4123
rect 15529 -4157 15563 -4155
rect 15723 -4053 15757 -4051
rect 15723 -4085 15757 -4053
rect 15723 -4155 15757 -4123
rect 15723 -4157 15757 -4155
rect 15981 -4053 16015 -4051
rect 15981 -4085 16015 -4053
rect 15981 -4155 16015 -4123
rect 15981 -4157 16015 -4155
rect 16239 -4053 16273 -4051
rect 16239 -4085 16273 -4053
rect 16239 -4155 16273 -4123
rect 16239 -4157 16273 -4155
rect 16497 -4053 16531 -4051
rect 16497 -4085 16531 -4053
rect 16497 -4155 16531 -4123
rect 16497 -4157 16531 -4155
rect 16691 -4053 16725 -4051
rect 16691 -4085 16725 -4053
rect 16691 -4155 16725 -4123
rect 16691 -4157 16725 -4155
rect 16949 -4053 16983 -4051
rect 16949 -4085 16983 -4053
rect 16949 -4155 16983 -4123
rect 16949 -4157 16983 -4155
rect 17207 -4053 17241 -4051
rect 17207 -4085 17241 -4053
rect 17207 -4155 17241 -4123
rect 17207 -4157 17241 -4155
rect 17465 -4053 17499 -4051
rect 17465 -4085 17499 -4053
rect 17465 -4155 17499 -4123
rect 17465 -4157 17499 -4155
rect 17723 -4053 17757 -4051
rect 17723 -4085 17757 -4053
rect 17723 -4155 17757 -4123
rect 17723 -4157 17757 -4155
rect 17917 -4053 17951 -4051
rect 17917 -4085 17951 -4053
rect 17917 -4155 17951 -4123
rect 17917 -4157 17951 -4155
rect 18175 -4053 18209 -4051
rect 18175 -4085 18209 -4053
rect 18175 -4155 18209 -4123
rect 18175 -4157 18209 -4155
rect 18290 -4034 18324 -4014
rect 18290 -4048 18324 -4034
rect 18290 -4102 18324 -4086
rect 18290 -4120 18324 -4102
rect 18290 -4192 18324 -4158
rect 5214 -4336 5248 -4302
rect 9781 -4285 9783 -4251
rect 9783 -4285 9815 -4251
rect 9853 -4285 9885 -4251
rect 9885 -4285 9887 -4251
rect 10233 -4285 10235 -4251
rect 10235 -4285 10267 -4251
rect 10305 -4285 10337 -4251
rect 10337 -4285 10339 -4251
rect 10491 -4285 10493 -4251
rect 10493 -4285 10525 -4251
rect 10563 -4285 10595 -4251
rect 10595 -4285 10597 -4251
rect 10749 -4285 10751 -4251
rect 10751 -4285 10783 -4251
rect 10821 -4285 10853 -4251
rect 10853 -4285 10855 -4251
rect 11007 -4285 11009 -4251
rect 11009 -4285 11041 -4251
rect 11079 -4285 11111 -4251
rect 11111 -4285 11113 -4251
rect 11459 -4285 11461 -4251
rect 11461 -4285 11493 -4251
rect 11531 -4285 11563 -4251
rect 11563 -4285 11565 -4251
rect 11717 -4285 11719 -4251
rect 11719 -4285 11751 -4251
rect 11789 -4285 11821 -4251
rect 11821 -4285 11823 -4251
rect 11975 -4285 11977 -4251
rect 11977 -4285 12009 -4251
rect 12047 -4285 12079 -4251
rect 12079 -4285 12081 -4251
rect 12427 -4285 12429 -4251
rect 12429 -4285 12461 -4251
rect 12499 -4285 12531 -4251
rect 12531 -4285 12533 -4251
rect 12685 -4285 12687 -4251
rect 12687 -4285 12719 -4251
rect 12757 -4285 12789 -4251
rect 12789 -4285 12791 -4251
rect 12943 -4285 12945 -4251
rect 12945 -4285 12977 -4251
rect 13015 -4285 13047 -4251
rect 13047 -4285 13049 -4251
rect 13201 -4285 13203 -4251
rect 13203 -4285 13235 -4251
rect 13273 -4285 13305 -4251
rect 13305 -4285 13307 -4251
rect 13653 -4285 13655 -4251
rect 13655 -4285 13687 -4251
rect 13725 -4285 13757 -4251
rect 13757 -4285 13759 -4251
rect 13932 -4264 13966 -4230
rect 9573 -4336 9607 -4302
rect 14139 -4285 14141 -4251
rect 14141 -4285 14173 -4251
rect 14211 -4285 14243 -4251
rect 14243 -4285 14245 -4251
rect 14590 -4285 14592 -4251
rect 14592 -4285 14624 -4251
rect 14662 -4285 14694 -4251
rect 14694 -4285 14696 -4251
rect 14848 -4285 14850 -4251
rect 14850 -4285 14882 -4251
rect 14920 -4285 14952 -4251
rect 14952 -4285 14954 -4251
rect 15106 -4285 15108 -4251
rect 15108 -4285 15140 -4251
rect 15178 -4285 15210 -4251
rect 15210 -4285 15212 -4251
rect 15364 -4285 15366 -4251
rect 15366 -4285 15398 -4251
rect 15436 -4285 15468 -4251
rect 15468 -4285 15470 -4251
rect 15816 -4285 15818 -4251
rect 15818 -4285 15850 -4251
rect 15888 -4285 15920 -4251
rect 15920 -4285 15922 -4251
rect 16074 -4285 16076 -4251
rect 16076 -4285 16108 -4251
rect 16146 -4285 16178 -4251
rect 16178 -4285 16180 -4251
rect 16332 -4285 16334 -4251
rect 16334 -4285 16366 -4251
rect 16404 -4285 16436 -4251
rect 16436 -4285 16438 -4251
rect 16784 -4285 16786 -4251
rect 16786 -4285 16818 -4251
rect 16856 -4285 16888 -4251
rect 16888 -4285 16890 -4251
rect 17042 -4285 17044 -4251
rect 17044 -4285 17076 -4251
rect 17114 -4285 17146 -4251
rect 17146 -4285 17148 -4251
rect 17300 -4285 17302 -4251
rect 17302 -4285 17334 -4251
rect 17372 -4285 17404 -4251
rect 17404 -4285 17406 -4251
rect 17558 -4285 17560 -4251
rect 17560 -4285 17592 -4251
rect 17630 -4285 17662 -4251
rect 17662 -4285 17664 -4251
rect 18010 -4285 18012 -4251
rect 18012 -4285 18044 -4251
rect 18082 -4285 18114 -4251
rect 18114 -4285 18116 -4251
rect 18290 -4264 18324 -4230
rect 13932 -4336 13966 -4302
rect 18290 -4336 18324 -4302
rect 930 -4399 964 -4365
rect 1002 -4399 1011 -4365
rect 1011 -4399 1036 -4365
rect 1074 -4399 1079 -4365
rect 1079 -4399 1108 -4365
rect 1146 -4399 1147 -4365
rect 1147 -4399 1180 -4365
rect 1218 -4399 1249 -4365
rect 1249 -4399 1252 -4365
rect 1290 -4399 1317 -4365
rect 1317 -4399 1324 -4365
rect 1362 -4399 1385 -4365
rect 1385 -4399 1396 -4365
rect 1434 -4399 1453 -4365
rect 1453 -4399 1468 -4365
rect 1506 -4399 1521 -4365
rect 1521 -4399 1540 -4365
rect 1578 -4399 1589 -4365
rect 1589 -4399 1612 -4365
rect 1650 -4399 1657 -4365
rect 1657 -4399 1684 -4365
rect 1722 -4399 1725 -4365
rect 1725 -4399 1756 -4365
rect 1794 -4399 1827 -4365
rect 1827 -4399 1828 -4365
rect 1866 -4399 1895 -4365
rect 1895 -4399 1900 -4365
rect 1938 -4399 1963 -4365
rect 1963 -4399 1972 -4365
rect 2010 -4399 2031 -4365
rect 2031 -4399 2044 -4365
rect 2082 -4399 2099 -4365
rect 2099 -4399 2116 -4365
rect 2154 -4399 2167 -4365
rect 2167 -4399 2188 -4365
rect 2226 -4399 2235 -4365
rect 2235 -4399 2260 -4365
rect 2298 -4399 2303 -4365
rect 2303 -4399 2332 -4365
rect 2370 -4399 2371 -4365
rect 2371 -4399 2404 -4365
rect 2442 -4399 2473 -4365
rect 2473 -4399 2476 -4365
rect 2514 -4399 2541 -4365
rect 2541 -4399 2548 -4365
rect 2586 -4399 2609 -4365
rect 2609 -4399 2620 -4365
rect 2658 -4399 2677 -4365
rect 2677 -4399 2692 -4365
rect 2730 -4399 2745 -4365
rect 2745 -4399 2764 -4365
rect 2802 -4399 2813 -4365
rect 2813 -4399 2836 -4365
rect 2874 -4399 2881 -4365
rect 2881 -4399 2908 -4365
rect 2946 -4399 2949 -4365
rect 2949 -4399 2980 -4365
rect 3018 -4399 3051 -4365
rect 3051 -4399 3052 -4365
rect 3090 -4399 3119 -4365
rect 3119 -4399 3124 -4365
rect 3162 -4399 3187 -4365
rect 3187 -4399 3196 -4365
rect 3234 -4399 3255 -4365
rect 3255 -4399 3268 -4365
rect 3306 -4399 3323 -4365
rect 3323 -4399 3340 -4365
rect 3378 -4399 3391 -4365
rect 3391 -4399 3412 -4365
rect 3450 -4399 3459 -4365
rect 3459 -4399 3484 -4365
rect 3522 -4399 3527 -4365
rect 3527 -4399 3556 -4365
rect 3594 -4399 3595 -4365
rect 3595 -4399 3628 -4365
rect 3666 -4399 3697 -4365
rect 3697 -4399 3700 -4365
rect 3738 -4399 3765 -4365
rect 3765 -4399 3772 -4365
rect 3810 -4399 3833 -4365
rect 3833 -4399 3844 -4365
rect 3882 -4399 3901 -4365
rect 3901 -4399 3916 -4365
rect 3954 -4399 3969 -4365
rect 3969 -4399 3988 -4365
rect 4026 -4399 4037 -4365
rect 4037 -4399 4060 -4365
rect 4098 -4399 4105 -4365
rect 4105 -4399 4132 -4365
rect 4170 -4399 4173 -4365
rect 4173 -4399 4204 -4365
rect 4242 -4399 4275 -4365
rect 4275 -4399 4276 -4365
rect 4314 -4399 4343 -4365
rect 4343 -4399 4348 -4365
rect 4386 -4399 4411 -4365
rect 4411 -4399 4420 -4365
rect 4458 -4399 4479 -4365
rect 4479 -4399 4492 -4365
rect 4530 -4399 4547 -4365
rect 4547 -4399 4564 -4365
rect 4602 -4399 4615 -4365
rect 4615 -4399 4636 -4365
rect 4674 -4399 4683 -4365
rect 4683 -4399 4708 -4365
rect 4746 -4399 4751 -4365
rect 4751 -4399 4780 -4365
rect 4818 -4399 4819 -4365
rect 4819 -4399 4852 -4365
rect 4890 -4399 4921 -4365
rect 4921 -4399 4924 -4365
rect 4962 -4399 4989 -4365
rect 4989 -4399 4996 -4365
rect 5034 -4399 5057 -4365
rect 5057 -4399 5068 -4365
rect 5106 -4399 5140 -4365
rect 5323 -4399 5357 -4365
rect 5395 -4399 5406 -4365
rect 5406 -4399 5429 -4365
rect 5467 -4399 5474 -4365
rect 5474 -4399 5501 -4365
rect 5539 -4399 5542 -4365
rect 5542 -4399 5573 -4365
rect 5611 -4399 5644 -4365
rect 5644 -4399 5645 -4365
rect 5683 -4399 5712 -4365
rect 5712 -4399 5717 -4365
rect 5755 -4399 5780 -4365
rect 5780 -4399 5789 -4365
rect 5827 -4399 5848 -4365
rect 5848 -4399 5861 -4365
rect 5899 -4399 5916 -4365
rect 5916 -4399 5933 -4365
rect 5971 -4399 5984 -4365
rect 5984 -4399 6005 -4365
rect 6043 -4399 6052 -4365
rect 6052 -4399 6077 -4365
rect 6115 -4399 6120 -4365
rect 6120 -4399 6149 -4365
rect 6187 -4399 6188 -4365
rect 6188 -4399 6221 -4365
rect 6259 -4399 6290 -4365
rect 6290 -4399 6293 -4365
rect 6331 -4399 6358 -4365
rect 6358 -4399 6365 -4365
rect 6403 -4399 6426 -4365
rect 6426 -4399 6437 -4365
rect 6475 -4399 6494 -4365
rect 6494 -4399 6509 -4365
rect 6547 -4399 6562 -4365
rect 6562 -4399 6581 -4365
rect 6619 -4399 6630 -4365
rect 6630 -4399 6653 -4365
rect 6691 -4399 6698 -4365
rect 6698 -4399 6725 -4365
rect 6763 -4399 6766 -4365
rect 6766 -4399 6797 -4365
rect 6835 -4399 6868 -4365
rect 6868 -4399 6869 -4365
rect 6907 -4399 6936 -4365
rect 6936 -4399 6941 -4365
rect 6979 -4399 7004 -4365
rect 7004 -4399 7013 -4365
rect 7051 -4399 7072 -4365
rect 7072 -4399 7085 -4365
rect 7123 -4399 7140 -4365
rect 7140 -4399 7157 -4365
rect 7195 -4399 7208 -4365
rect 7208 -4399 7229 -4365
rect 7267 -4399 7276 -4365
rect 7276 -4399 7301 -4365
rect 7339 -4399 7344 -4365
rect 7344 -4399 7373 -4365
rect 7411 -4399 7412 -4365
rect 7412 -4399 7445 -4365
rect 7483 -4399 7514 -4365
rect 7514 -4399 7517 -4365
rect 7555 -4399 7582 -4365
rect 7582 -4399 7589 -4365
rect 7627 -4399 7650 -4365
rect 7650 -4399 7661 -4365
rect 7699 -4399 7718 -4365
rect 7718 -4399 7733 -4365
rect 7771 -4399 7786 -4365
rect 7786 -4399 7805 -4365
rect 7843 -4399 7854 -4365
rect 7854 -4399 7877 -4365
rect 7915 -4399 7922 -4365
rect 7922 -4399 7949 -4365
rect 7987 -4399 7990 -4365
rect 7990 -4399 8021 -4365
rect 8059 -4399 8092 -4365
rect 8092 -4399 8093 -4365
rect 8131 -4399 8160 -4365
rect 8160 -4399 8165 -4365
rect 8203 -4399 8228 -4365
rect 8228 -4399 8237 -4365
rect 8275 -4399 8296 -4365
rect 8296 -4399 8309 -4365
rect 8347 -4399 8364 -4365
rect 8364 -4399 8381 -4365
rect 8419 -4399 8432 -4365
rect 8432 -4399 8453 -4365
rect 8491 -4399 8500 -4365
rect 8500 -4399 8525 -4365
rect 8563 -4399 8568 -4365
rect 8568 -4399 8597 -4365
rect 8635 -4399 8636 -4365
rect 8636 -4399 8669 -4365
rect 8707 -4399 8738 -4365
rect 8738 -4399 8741 -4365
rect 8779 -4399 8806 -4365
rect 8806 -4399 8813 -4365
rect 8851 -4399 8874 -4365
rect 8874 -4399 8885 -4365
rect 8923 -4399 8942 -4365
rect 8942 -4399 8957 -4365
rect 8995 -4399 9010 -4365
rect 9010 -4399 9029 -4365
rect 9067 -4399 9078 -4365
rect 9078 -4399 9101 -4365
rect 9139 -4399 9146 -4365
rect 9146 -4399 9173 -4365
rect 9211 -4399 9214 -4365
rect 9214 -4399 9245 -4365
rect 9283 -4399 9316 -4365
rect 9316 -4399 9317 -4365
rect 9355 -4399 9384 -4365
rect 9384 -4399 9389 -4365
rect 9427 -4399 9452 -4365
rect 9452 -4399 9461 -4365
rect 9499 -4399 9533 -4365
rect 9647 -4399 9681 -4365
rect 9719 -4399 9728 -4365
rect 9728 -4399 9753 -4365
rect 9791 -4399 9796 -4365
rect 9796 -4399 9825 -4365
rect 9863 -4399 9864 -4365
rect 9864 -4399 9897 -4365
rect 9935 -4399 9966 -4365
rect 9966 -4399 9969 -4365
rect 10007 -4399 10034 -4365
rect 10034 -4399 10041 -4365
rect 10079 -4399 10102 -4365
rect 10102 -4399 10113 -4365
rect 10151 -4399 10170 -4365
rect 10170 -4399 10185 -4365
rect 10223 -4399 10238 -4365
rect 10238 -4399 10257 -4365
rect 10295 -4399 10306 -4365
rect 10306 -4399 10329 -4365
rect 10367 -4399 10374 -4365
rect 10374 -4399 10401 -4365
rect 10439 -4399 10442 -4365
rect 10442 -4399 10473 -4365
rect 10511 -4399 10544 -4365
rect 10544 -4399 10545 -4365
rect 10583 -4399 10612 -4365
rect 10612 -4399 10617 -4365
rect 10655 -4399 10680 -4365
rect 10680 -4399 10689 -4365
rect 10727 -4399 10748 -4365
rect 10748 -4399 10761 -4365
rect 10799 -4399 10816 -4365
rect 10816 -4399 10833 -4365
rect 10871 -4399 10884 -4365
rect 10884 -4399 10905 -4365
rect 10943 -4399 10952 -4365
rect 10952 -4399 10977 -4365
rect 11015 -4399 11020 -4365
rect 11020 -4399 11049 -4365
rect 11087 -4399 11088 -4365
rect 11088 -4399 11121 -4365
rect 11159 -4399 11190 -4365
rect 11190 -4399 11193 -4365
rect 11231 -4399 11258 -4365
rect 11258 -4399 11265 -4365
rect 11303 -4399 11326 -4365
rect 11326 -4399 11337 -4365
rect 11375 -4399 11394 -4365
rect 11394 -4399 11409 -4365
rect 11447 -4399 11462 -4365
rect 11462 -4399 11481 -4365
rect 11519 -4399 11530 -4365
rect 11530 -4399 11553 -4365
rect 11591 -4399 11598 -4365
rect 11598 -4399 11625 -4365
rect 11663 -4399 11666 -4365
rect 11666 -4399 11697 -4365
rect 11735 -4399 11768 -4365
rect 11768 -4399 11769 -4365
rect 11807 -4399 11836 -4365
rect 11836 -4399 11841 -4365
rect 11879 -4399 11904 -4365
rect 11904 -4399 11913 -4365
rect 11951 -4399 11972 -4365
rect 11972 -4399 11985 -4365
rect 12023 -4399 12040 -4365
rect 12040 -4399 12057 -4365
rect 12095 -4399 12108 -4365
rect 12108 -4399 12129 -4365
rect 12167 -4399 12176 -4365
rect 12176 -4399 12201 -4365
rect 12239 -4399 12244 -4365
rect 12244 -4399 12273 -4365
rect 12311 -4399 12312 -4365
rect 12312 -4399 12345 -4365
rect 12383 -4399 12414 -4365
rect 12414 -4399 12417 -4365
rect 12455 -4399 12482 -4365
rect 12482 -4399 12489 -4365
rect 12527 -4399 12550 -4365
rect 12550 -4399 12561 -4365
rect 12599 -4399 12618 -4365
rect 12618 -4399 12633 -4365
rect 12671 -4399 12686 -4365
rect 12686 -4399 12705 -4365
rect 12743 -4399 12754 -4365
rect 12754 -4399 12777 -4365
rect 12815 -4399 12822 -4365
rect 12822 -4399 12849 -4365
rect 12887 -4399 12890 -4365
rect 12890 -4399 12921 -4365
rect 12959 -4399 12992 -4365
rect 12992 -4399 12993 -4365
rect 13031 -4399 13060 -4365
rect 13060 -4399 13065 -4365
rect 13103 -4399 13128 -4365
rect 13128 -4399 13137 -4365
rect 13175 -4399 13196 -4365
rect 13196 -4399 13209 -4365
rect 13247 -4399 13264 -4365
rect 13264 -4399 13281 -4365
rect 13319 -4399 13332 -4365
rect 13332 -4399 13353 -4365
rect 13391 -4399 13400 -4365
rect 13400 -4399 13425 -4365
rect 13463 -4399 13468 -4365
rect 13468 -4399 13497 -4365
rect 13535 -4399 13536 -4365
rect 13536 -4399 13569 -4365
rect 13607 -4399 13638 -4365
rect 13638 -4399 13641 -4365
rect 13679 -4399 13706 -4365
rect 13706 -4399 13713 -4365
rect 13751 -4399 13774 -4365
rect 13774 -4399 13785 -4365
rect 13823 -4399 13857 -4365
rect 14040 -4399 14074 -4365
rect 14112 -4399 14123 -4365
rect 14123 -4399 14146 -4365
rect 14184 -4399 14191 -4365
rect 14191 -4399 14218 -4365
rect 14256 -4399 14259 -4365
rect 14259 -4399 14290 -4365
rect 14328 -4399 14361 -4365
rect 14361 -4399 14362 -4365
rect 14400 -4399 14429 -4365
rect 14429 -4399 14434 -4365
rect 14472 -4399 14497 -4365
rect 14497 -4399 14506 -4365
rect 14544 -4399 14565 -4365
rect 14565 -4399 14578 -4365
rect 14616 -4399 14633 -4365
rect 14633 -4399 14650 -4365
rect 14688 -4399 14701 -4365
rect 14701 -4399 14722 -4365
rect 14760 -4399 14769 -4365
rect 14769 -4399 14794 -4365
rect 14832 -4399 14837 -4365
rect 14837 -4399 14866 -4365
rect 14904 -4399 14905 -4365
rect 14905 -4399 14938 -4365
rect 14976 -4399 15007 -4365
rect 15007 -4399 15010 -4365
rect 15048 -4399 15075 -4365
rect 15075 -4399 15082 -4365
rect 15120 -4399 15143 -4365
rect 15143 -4399 15154 -4365
rect 15192 -4399 15211 -4365
rect 15211 -4399 15226 -4365
rect 15264 -4399 15279 -4365
rect 15279 -4399 15298 -4365
rect 15336 -4399 15347 -4365
rect 15347 -4399 15370 -4365
rect 15408 -4399 15415 -4365
rect 15415 -4399 15442 -4365
rect 15480 -4399 15483 -4365
rect 15483 -4399 15514 -4365
rect 15552 -4399 15585 -4365
rect 15585 -4399 15586 -4365
rect 15624 -4399 15653 -4365
rect 15653 -4399 15658 -4365
rect 15696 -4399 15721 -4365
rect 15721 -4399 15730 -4365
rect 15768 -4399 15789 -4365
rect 15789 -4399 15802 -4365
rect 15840 -4399 15857 -4365
rect 15857 -4399 15874 -4365
rect 15912 -4399 15925 -4365
rect 15925 -4399 15946 -4365
rect 15984 -4399 15993 -4365
rect 15993 -4399 16018 -4365
rect 16056 -4399 16061 -4365
rect 16061 -4399 16090 -4365
rect 16128 -4399 16129 -4365
rect 16129 -4399 16162 -4365
rect 16200 -4399 16231 -4365
rect 16231 -4399 16234 -4365
rect 16272 -4399 16299 -4365
rect 16299 -4399 16306 -4365
rect 16344 -4399 16367 -4365
rect 16367 -4399 16378 -4365
rect 16416 -4399 16435 -4365
rect 16435 -4399 16450 -4365
rect 16488 -4399 16503 -4365
rect 16503 -4399 16522 -4365
rect 16560 -4399 16571 -4365
rect 16571 -4399 16594 -4365
rect 16632 -4399 16639 -4365
rect 16639 -4399 16666 -4365
rect 16704 -4399 16707 -4365
rect 16707 -4399 16738 -4365
rect 16776 -4399 16809 -4365
rect 16809 -4399 16810 -4365
rect 16848 -4399 16877 -4365
rect 16877 -4399 16882 -4365
rect 16920 -4399 16945 -4365
rect 16945 -4399 16954 -4365
rect 16992 -4399 17013 -4365
rect 17013 -4399 17026 -4365
rect 17064 -4399 17081 -4365
rect 17081 -4399 17098 -4365
rect 17136 -4399 17149 -4365
rect 17149 -4399 17170 -4365
rect 17208 -4399 17217 -4365
rect 17217 -4399 17242 -4365
rect 17280 -4399 17285 -4365
rect 17285 -4399 17314 -4365
rect 17352 -4399 17353 -4365
rect 17353 -4399 17386 -4365
rect 17424 -4399 17455 -4365
rect 17455 -4399 17458 -4365
rect 17496 -4399 17523 -4365
rect 17523 -4399 17530 -4365
rect 17568 -4399 17591 -4365
rect 17591 -4399 17602 -4365
rect 17640 -4399 17659 -4365
rect 17659 -4399 17674 -4365
rect 17712 -4399 17727 -4365
rect 17727 -4399 17746 -4365
rect 17784 -4399 17795 -4365
rect 17795 -4399 17818 -4365
rect 17856 -4399 17863 -4365
rect 17863 -4399 17890 -4365
rect 17928 -4399 17931 -4365
rect 17931 -4399 17962 -4365
rect 18000 -4399 18033 -4365
rect 18033 -4399 18034 -4365
rect 18072 -4399 18101 -4365
rect 18101 -4399 18106 -4365
rect 18144 -4399 18169 -4365
rect 18169 -4399 18178 -4365
rect 18216 -4399 18250 -4365
rect 856 -4462 890 -4428
rect 5214 -4462 5248 -4428
rect 856 -4534 890 -4500
rect 1064 -4513 1066 -4479
rect 1066 -4513 1098 -4479
rect 1136 -4513 1168 -4479
rect 1168 -4513 1170 -4479
rect 1516 -4513 1518 -4479
rect 1518 -4513 1550 -4479
rect 1588 -4513 1620 -4479
rect 1620 -4513 1622 -4479
rect 1774 -4513 1776 -4479
rect 1776 -4513 1808 -4479
rect 1846 -4513 1878 -4479
rect 1878 -4513 1880 -4479
rect 2032 -4513 2034 -4479
rect 2034 -4513 2066 -4479
rect 2104 -4513 2136 -4479
rect 2136 -4513 2138 -4479
rect 2290 -4513 2292 -4479
rect 2292 -4513 2324 -4479
rect 2362 -4513 2394 -4479
rect 2394 -4513 2396 -4479
rect 2742 -4513 2744 -4479
rect 2744 -4513 2776 -4479
rect 2814 -4513 2846 -4479
rect 2846 -4513 2848 -4479
rect 3000 -4513 3002 -4479
rect 3002 -4513 3034 -4479
rect 3072 -4513 3104 -4479
rect 3104 -4513 3106 -4479
rect 3258 -4513 3260 -4479
rect 3260 -4513 3292 -4479
rect 3330 -4513 3362 -4479
rect 3362 -4513 3364 -4479
rect 3710 -4513 3712 -4479
rect 3712 -4513 3744 -4479
rect 3782 -4513 3814 -4479
rect 3814 -4513 3816 -4479
rect 3968 -4513 3970 -4479
rect 3970 -4513 4002 -4479
rect 4040 -4513 4072 -4479
rect 4072 -4513 4074 -4479
rect 4226 -4513 4228 -4479
rect 4228 -4513 4260 -4479
rect 4298 -4513 4330 -4479
rect 4330 -4513 4332 -4479
rect 4484 -4513 4486 -4479
rect 4486 -4513 4518 -4479
rect 4556 -4513 4588 -4479
rect 4588 -4513 4590 -4479
rect 4935 -4513 4937 -4479
rect 4937 -4513 4969 -4479
rect 5007 -4513 5039 -4479
rect 5039 -4513 5041 -4479
rect 9573 -4462 9607 -4428
rect 5214 -4534 5248 -4500
rect 5421 -4513 5423 -4479
rect 5423 -4513 5455 -4479
rect 5493 -4513 5525 -4479
rect 5525 -4513 5527 -4479
rect 5873 -4513 5875 -4479
rect 5875 -4513 5907 -4479
rect 5945 -4513 5977 -4479
rect 5977 -4513 5979 -4479
rect 6131 -4513 6133 -4479
rect 6133 -4513 6165 -4479
rect 6203 -4513 6235 -4479
rect 6235 -4513 6237 -4479
rect 6389 -4513 6391 -4479
rect 6391 -4513 6423 -4479
rect 6461 -4513 6493 -4479
rect 6493 -4513 6495 -4479
rect 6647 -4513 6649 -4479
rect 6649 -4513 6681 -4479
rect 6719 -4513 6751 -4479
rect 6751 -4513 6753 -4479
rect 7099 -4513 7101 -4479
rect 7101 -4513 7133 -4479
rect 7171 -4513 7203 -4479
rect 7203 -4513 7205 -4479
rect 7357 -4513 7359 -4479
rect 7359 -4513 7391 -4479
rect 7429 -4513 7461 -4479
rect 7461 -4513 7463 -4479
rect 7615 -4513 7617 -4479
rect 7617 -4513 7649 -4479
rect 7687 -4513 7719 -4479
rect 7719 -4513 7721 -4479
rect 8067 -4513 8069 -4479
rect 8069 -4513 8101 -4479
rect 8139 -4513 8171 -4479
rect 8171 -4513 8173 -4479
rect 8325 -4513 8327 -4479
rect 8327 -4513 8359 -4479
rect 8397 -4513 8429 -4479
rect 8429 -4513 8431 -4479
rect 8583 -4513 8585 -4479
rect 8585 -4513 8617 -4479
rect 8655 -4513 8687 -4479
rect 8687 -4513 8689 -4479
rect 8841 -4513 8843 -4479
rect 8843 -4513 8875 -4479
rect 8913 -4513 8945 -4479
rect 8945 -4513 8947 -4479
rect 9293 -4513 9295 -4479
rect 9295 -4513 9327 -4479
rect 9365 -4513 9397 -4479
rect 9397 -4513 9399 -4479
rect 13932 -4462 13966 -4428
rect 856 -4606 890 -4572
rect 856 -4662 890 -4644
rect 856 -4678 890 -4662
rect 856 -4730 890 -4716
rect 856 -4750 890 -4730
rect 971 -4609 1005 -4607
rect 971 -4641 1005 -4609
rect 971 -4711 1005 -4679
rect 971 -4713 1005 -4711
rect 1229 -4609 1263 -4607
rect 1229 -4641 1263 -4609
rect 1229 -4711 1263 -4679
rect 1229 -4713 1263 -4711
rect 1423 -4609 1457 -4607
rect 1423 -4641 1457 -4609
rect 1423 -4711 1457 -4679
rect 1423 -4713 1457 -4711
rect 1681 -4609 1715 -4607
rect 1681 -4641 1715 -4609
rect 1681 -4711 1715 -4679
rect 1681 -4713 1715 -4711
rect 1939 -4609 1973 -4607
rect 1939 -4641 1973 -4609
rect 1939 -4711 1973 -4679
rect 1939 -4713 1973 -4711
rect 2197 -4609 2231 -4607
rect 2197 -4641 2231 -4609
rect 2197 -4711 2231 -4679
rect 2197 -4713 2231 -4711
rect 2455 -4609 2489 -4607
rect 2455 -4641 2489 -4609
rect 2455 -4711 2489 -4679
rect 2455 -4713 2489 -4711
rect 2649 -4609 2683 -4607
rect 2649 -4641 2683 -4609
rect 2649 -4711 2683 -4679
rect 2649 -4713 2683 -4711
rect 2907 -4609 2941 -4607
rect 2907 -4641 2941 -4609
rect 2907 -4711 2941 -4679
rect 2907 -4713 2941 -4711
rect 3165 -4609 3199 -4607
rect 3165 -4641 3199 -4609
rect 3165 -4711 3199 -4679
rect 3165 -4713 3199 -4711
rect 3423 -4609 3457 -4607
rect 3423 -4641 3457 -4609
rect 3423 -4711 3457 -4679
rect 3423 -4713 3457 -4711
rect 3617 -4609 3651 -4607
rect 3617 -4641 3651 -4609
rect 3617 -4711 3651 -4679
rect 3617 -4713 3651 -4711
rect 3875 -4609 3909 -4607
rect 3875 -4641 3909 -4609
rect 3875 -4711 3909 -4679
rect 3875 -4713 3909 -4711
rect 4133 -4609 4167 -4607
rect 4133 -4641 4167 -4609
rect 4133 -4711 4167 -4679
rect 4133 -4713 4167 -4711
rect 4391 -4609 4425 -4607
rect 4391 -4641 4425 -4609
rect 4391 -4711 4425 -4679
rect 4391 -4713 4425 -4711
rect 4649 -4609 4683 -4607
rect 4649 -4641 4683 -4609
rect 4649 -4711 4683 -4679
rect 4649 -4713 4683 -4711
rect 4842 -4609 4876 -4607
rect 4842 -4641 4876 -4609
rect 4842 -4711 4876 -4679
rect 4842 -4713 4876 -4711
rect 5100 -4609 5134 -4607
rect 5100 -4641 5134 -4609
rect 5100 -4711 5134 -4679
rect 5100 -4713 5134 -4711
rect 9573 -4534 9607 -4500
rect 9781 -4513 9783 -4479
rect 9783 -4513 9815 -4479
rect 9853 -4513 9885 -4479
rect 9885 -4513 9887 -4479
rect 10233 -4513 10235 -4479
rect 10235 -4513 10267 -4479
rect 10305 -4513 10337 -4479
rect 10337 -4513 10339 -4479
rect 10491 -4513 10493 -4479
rect 10493 -4513 10525 -4479
rect 10563 -4513 10595 -4479
rect 10595 -4513 10597 -4479
rect 10749 -4513 10751 -4479
rect 10751 -4513 10783 -4479
rect 10821 -4513 10853 -4479
rect 10853 -4513 10855 -4479
rect 11007 -4513 11009 -4479
rect 11009 -4513 11041 -4479
rect 11079 -4513 11111 -4479
rect 11111 -4513 11113 -4479
rect 11459 -4513 11461 -4479
rect 11461 -4513 11493 -4479
rect 11531 -4513 11563 -4479
rect 11563 -4513 11565 -4479
rect 11717 -4513 11719 -4479
rect 11719 -4513 11751 -4479
rect 11789 -4513 11821 -4479
rect 11821 -4513 11823 -4479
rect 11975 -4513 11977 -4479
rect 11977 -4513 12009 -4479
rect 12047 -4513 12079 -4479
rect 12079 -4513 12081 -4479
rect 12427 -4513 12429 -4479
rect 12429 -4513 12461 -4479
rect 12499 -4513 12531 -4479
rect 12531 -4513 12533 -4479
rect 12685 -4513 12687 -4479
rect 12687 -4513 12719 -4479
rect 12757 -4513 12789 -4479
rect 12789 -4513 12791 -4479
rect 12943 -4513 12945 -4479
rect 12945 -4513 12977 -4479
rect 13015 -4513 13047 -4479
rect 13047 -4513 13049 -4479
rect 13201 -4513 13203 -4479
rect 13203 -4513 13235 -4479
rect 13273 -4513 13305 -4479
rect 13305 -4513 13307 -4479
rect 13653 -4513 13655 -4479
rect 13655 -4513 13687 -4479
rect 13725 -4513 13757 -4479
rect 13757 -4513 13759 -4479
rect 18290 -4462 18324 -4428
rect 5214 -4606 5248 -4572
rect 5214 -4662 5248 -4644
rect 5214 -4678 5248 -4662
rect 5214 -4730 5248 -4716
rect 5214 -4750 5248 -4730
rect 5328 -4609 5362 -4607
rect 5328 -4641 5362 -4609
rect 5328 -4711 5362 -4679
rect 5328 -4713 5362 -4711
rect 5586 -4609 5620 -4607
rect 5586 -4641 5620 -4609
rect 5586 -4711 5620 -4679
rect 5586 -4713 5620 -4711
rect 5780 -4609 5814 -4607
rect 5780 -4641 5814 -4609
rect 5780 -4711 5814 -4679
rect 5780 -4713 5814 -4711
rect 6038 -4609 6072 -4607
rect 6038 -4641 6072 -4609
rect 6038 -4711 6072 -4679
rect 6038 -4713 6072 -4711
rect 6296 -4609 6330 -4607
rect 6296 -4641 6330 -4609
rect 6296 -4711 6330 -4679
rect 6296 -4713 6330 -4711
rect 6554 -4609 6588 -4607
rect 6554 -4641 6588 -4609
rect 6554 -4711 6588 -4679
rect 6554 -4713 6588 -4711
rect 6812 -4609 6846 -4607
rect 6812 -4641 6846 -4609
rect 6812 -4711 6846 -4679
rect 6812 -4713 6846 -4711
rect 7006 -4609 7040 -4607
rect 7006 -4641 7040 -4609
rect 7006 -4711 7040 -4679
rect 7006 -4713 7040 -4711
rect 7264 -4609 7298 -4607
rect 7264 -4641 7298 -4609
rect 7264 -4711 7298 -4679
rect 7264 -4713 7298 -4711
rect 7522 -4609 7556 -4607
rect 7522 -4641 7556 -4609
rect 7522 -4711 7556 -4679
rect 7522 -4713 7556 -4711
rect 7780 -4609 7814 -4607
rect 7780 -4641 7814 -4609
rect 7780 -4711 7814 -4679
rect 7780 -4713 7814 -4711
rect 7974 -4609 8008 -4607
rect 7974 -4641 8008 -4609
rect 7974 -4711 8008 -4679
rect 7974 -4713 8008 -4711
rect 8232 -4609 8266 -4607
rect 8232 -4641 8266 -4609
rect 8232 -4711 8266 -4679
rect 8232 -4713 8266 -4711
rect 8490 -4609 8524 -4607
rect 8490 -4641 8524 -4609
rect 8490 -4711 8524 -4679
rect 8490 -4713 8524 -4711
rect 8748 -4609 8782 -4607
rect 8748 -4641 8782 -4609
rect 8748 -4711 8782 -4679
rect 8748 -4713 8782 -4711
rect 9006 -4609 9040 -4607
rect 9006 -4641 9040 -4609
rect 9006 -4711 9040 -4679
rect 9006 -4713 9040 -4711
rect 9200 -4609 9234 -4607
rect 9200 -4641 9234 -4609
rect 9200 -4711 9234 -4679
rect 9200 -4713 9234 -4711
rect 9458 -4609 9492 -4607
rect 9458 -4641 9492 -4609
rect 9458 -4711 9492 -4679
rect 9458 -4713 9492 -4711
rect 13932 -4534 13966 -4500
rect 14139 -4513 14141 -4479
rect 14141 -4513 14173 -4479
rect 14211 -4513 14243 -4479
rect 14243 -4513 14245 -4479
rect 14590 -4513 14592 -4479
rect 14592 -4513 14624 -4479
rect 14662 -4513 14694 -4479
rect 14694 -4513 14696 -4479
rect 14848 -4513 14850 -4479
rect 14850 -4513 14882 -4479
rect 14920 -4513 14952 -4479
rect 14952 -4513 14954 -4479
rect 15106 -4513 15108 -4479
rect 15108 -4513 15140 -4479
rect 15178 -4513 15210 -4479
rect 15210 -4513 15212 -4479
rect 15364 -4513 15366 -4479
rect 15366 -4513 15398 -4479
rect 15436 -4513 15468 -4479
rect 15468 -4513 15470 -4479
rect 15816 -4513 15818 -4479
rect 15818 -4513 15850 -4479
rect 15888 -4513 15920 -4479
rect 15920 -4513 15922 -4479
rect 16074 -4513 16076 -4479
rect 16076 -4513 16108 -4479
rect 16146 -4513 16178 -4479
rect 16178 -4513 16180 -4479
rect 16332 -4513 16334 -4479
rect 16334 -4513 16366 -4479
rect 16404 -4513 16436 -4479
rect 16436 -4513 16438 -4479
rect 16784 -4513 16786 -4479
rect 16786 -4513 16818 -4479
rect 16856 -4513 16888 -4479
rect 16888 -4513 16890 -4479
rect 17042 -4513 17044 -4479
rect 17044 -4513 17076 -4479
rect 17114 -4513 17146 -4479
rect 17146 -4513 17148 -4479
rect 17300 -4513 17302 -4479
rect 17302 -4513 17334 -4479
rect 17372 -4513 17404 -4479
rect 17404 -4513 17406 -4479
rect 17558 -4513 17560 -4479
rect 17560 -4513 17592 -4479
rect 17630 -4513 17662 -4479
rect 17662 -4513 17664 -4479
rect 18010 -4513 18012 -4479
rect 18012 -4513 18044 -4479
rect 18082 -4513 18114 -4479
rect 18114 -4513 18116 -4479
rect 9573 -4606 9607 -4572
rect 9573 -4662 9607 -4644
rect 9573 -4678 9607 -4662
rect 9573 -4730 9607 -4716
rect 9573 -4750 9607 -4730
rect 9688 -4609 9722 -4607
rect 9688 -4641 9722 -4609
rect 9688 -4711 9722 -4679
rect 9688 -4713 9722 -4711
rect 9946 -4609 9980 -4607
rect 9946 -4641 9980 -4609
rect 9946 -4711 9980 -4679
rect 9946 -4713 9980 -4711
rect 10140 -4609 10174 -4607
rect 10140 -4641 10174 -4609
rect 10140 -4711 10174 -4679
rect 10140 -4713 10174 -4711
rect 10398 -4609 10432 -4607
rect 10398 -4641 10432 -4609
rect 10398 -4711 10432 -4679
rect 10398 -4713 10432 -4711
rect 10656 -4609 10690 -4607
rect 10656 -4641 10690 -4609
rect 10656 -4711 10690 -4679
rect 10656 -4713 10690 -4711
rect 10914 -4609 10948 -4607
rect 10914 -4641 10948 -4609
rect 10914 -4711 10948 -4679
rect 10914 -4713 10948 -4711
rect 11172 -4609 11206 -4607
rect 11172 -4641 11206 -4609
rect 11172 -4711 11206 -4679
rect 11172 -4713 11206 -4711
rect 11366 -4609 11400 -4607
rect 11366 -4641 11400 -4609
rect 11366 -4711 11400 -4679
rect 11366 -4713 11400 -4711
rect 11624 -4609 11658 -4607
rect 11624 -4641 11658 -4609
rect 11624 -4711 11658 -4679
rect 11624 -4713 11658 -4711
rect 11882 -4609 11916 -4607
rect 11882 -4641 11916 -4609
rect 11882 -4711 11916 -4679
rect 11882 -4713 11916 -4711
rect 12140 -4609 12174 -4607
rect 12140 -4641 12174 -4609
rect 12140 -4711 12174 -4679
rect 12140 -4713 12174 -4711
rect 12334 -4609 12368 -4607
rect 12334 -4641 12368 -4609
rect 12334 -4711 12368 -4679
rect 12334 -4713 12368 -4711
rect 12592 -4609 12626 -4607
rect 12592 -4641 12626 -4609
rect 12592 -4711 12626 -4679
rect 12592 -4713 12626 -4711
rect 12850 -4609 12884 -4607
rect 12850 -4641 12884 -4609
rect 12850 -4711 12884 -4679
rect 12850 -4713 12884 -4711
rect 13108 -4609 13142 -4607
rect 13108 -4641 13142 -4609
rect 13108 -4711 13142 -4679
rect 13108 -4713 13142 -4711
rect 13366 -4609 13400 -4607
rect 13366 -4641 13400 -4609
rect 13366 -4711 13400 -4679
rect 13366 -4713 13400 -4711
rect 13560 -4609 13594 -4607
rect 13560 -4641 13594 -4609
rect 13560 -4711 13594 -4679
rect 13560 -4713 13594 -4711
rect 13818 -4609 13852 -4607
rect 13818 -4641 13852 -4609
rect 13818 -4711 13852 -4679
rect 13818 -4713 13852 -4711
rect 18290 -4534 18324 -4500
rect 13932 -4606 13966 -4572
rect 13932 -4662 13966 -4644
rect 13932 -4678 13966 -4662
rect 13932 -4730 13966 -4716
rect 13932 -4750 13966 -4730
rect 14046 -4609 14080 -4607
rect 14046 -4641 14080 -4609
rect 14046 -4711 14080 -4679
rect 14046 -4713 14080 -4711
rect 14304 -4609 14338 -4607
rect 14304 -4641 14338 -4609
rect 14304 -4711 14338 -4679
rect 14304 -4713 14338 -4711
rect 14497 -4609 14531 -4607
rect 14497 -4641 14531 -4609
rect 14497 -4711 14531 -4679
rect 14497 -4713 14531 -4711
rect 14755 -4609 14789 -4607
rect 14755 -4641 14789 -4609
rect 14755 -4711 14789 -4679
rect 14755 -4713 14789 -4711
rect 15013 -4609 15047 -4607
rect 15013 -4641 15047 -4609
rect 15013 -4711 15047 -4679
rect 15013 -4713 15047 -4711
rect 15271 -4609 15305 -4607
rect 15271 -4641 15305 -4609
rect 15271 -4711 15305 -4679
rect 15271 -4713 15305 -4711
rect 15529 -4609 15563 -4607
rect 15529 -4641 15563 -4609
rect 15529 -4711 15563 -4679
rect 15529 -4713 15563 -4711
rect 15723 -4609 15757 -4607
rect 15723 -4641 15757 -4609
rect 15723 -4711 15757 -4679
rect 15723 -4713 15757 -4711
rect 15981 -4609 16015 -4607
rect 15981 -4641 16015 -4609
rect 15981 -4711 16015 -4679
rect 15981 -4713 16015 -4711
rect 16239 -4609 16273 -4607
rect 16239 -4641 16273 -4609
rect 16239 -4711 16273 -4679
rect 16239 -4713 16273 -4711
rect 16497 -4609 16531 -4607
rect 16497 -4641 16531 -4609
rect 16497 -4711 16531 -4679
rect 16497 -4713 16531 -4711
rect 16691 -4609 16725 -4607
rect 16691 -4641 16725 -4609
rect 16691 -4711 16725 -4679
rect 16691 -4713 16725 -4711
rect 16949 -4609 16983 -4607
rect 16949 -4641 16983 -4609
rect 16949 -4711 16983 -4679
rect 16949 -4713 16983 -4711
rect 17207 -4609 17241 -4607
rect 17207 -4641 17241 -4609
rect 17207 -4711 17241 -4679
rect 17207 -4713 17241 -4711
rect 17465 -4609 17499 -4607
rect 17465 -4641 17499 -4609
rect 17465 -4711 17499 -4679
rect 17465 -4713 17499 -4711
rect 17723 -4609 17757 -4607
rect 17723 -4641 17757 -4609
rect 17723 -4711 17757 -4679
rect 17723 -4713 17757 -4711
rect 17917 -4609 17951 -4607
rect 17917 -4641 17951 -4609
rect 17917 -4711 17951 -4679
rect 17917 -4713 17951 -4711
rect 18175 -4609 18209 -4607
rect 18175 -4641 18209 -4609
rect 18175 -4711 18209 -4679
rect 18175 -4713 18209 -4711
rect 18290 -4606 18324 -4572
rect 18290 -4662 18324 -4644
rect 18290 -4678 18324 -4662
rect 18290 -4730 18324 -4716
rect 18290 -4750 18324 -4730
rect 856 -4798 890 -4788
rect 856 -4822 890 -4798
rect 856 -4866 890 -4860
rect 856 -4894 890 -4866
rect 856 -4934 890 -4932
rect 856 -4966 890 -4934
rect 856 -5036 890 -5004
rect 856 -5038 890 -5036
rect 856 -5104 890 -5076
rect 856 -5110 890 -5104
rect 5214 -4798 5248 -4788
rect 5214 -4822 5248 -4798
rect 5214 -4866 5248 -4860
rect 5214 -4894 5248 -4866
rect 5214 -4934 5248 -4932
rect 5214 -4966 5248 -4934
rect 5214 -5036 5248 -5004
rect 5214 -5038 5248 -5036
rect 5214 -5104 5248 -5076
rect 5214 -5110 5248 -5104
rect 9573 -4798 9607 -4788
rect 9573 -4822 9607 -4798
rect 9573 -4866 9607 -4860
rect 9573 -4894 9607 -4866
rect 9573 -4934 9607 -4932
rect 9573 -4966 9607 -4934
rect 9573 -5036 9607 -5004
rect 9573 -5038 9607 -5036
rect 9573 -5104 9607 -5076
rect 9573 -5110 9607 -5104
rect 13932 -4798 13966 -4788
rect 13932 -4822 13966 -4798
rect 13932 -4866 13966 -4860
rect 13932 -4894 13966 -4866
rect 13932 -4934 13966 -4932
rect 13932 -4966 13966 -4934
rect 13932 -5036 13966 -5004
rect 13932 -5038 13966 -5036
rect 13932 -5104 13966 -5076
rect 13932 -5110 13966 -5104
rect 18290 -4798 18324 -4788
rect 18290 -4822 18324 -4798
rect 18290 -4866 18324 -4860
rect 18290 -4894 18324 -4866
rect 18290 -4934 18324 -4932
rect 18290 -4966 18324 -4934
rect 18290 -5036 18324 -5004
rect 18290 -5038 18324 -5036
rect 18290 -5104 18324 -5076
rect 18290 -5110 18324 -5104
rect 856 -5172 890 -5148
rect 5214 -5172 5248 -5148
rect 9573 -5172 9607 -5148
rect 13932 -5172 13966 -5148
rect 18290 -5172 18324 -5148
rect 856 -5182 890 -5172
rect 856 -5240 890 -5220
rect 856 -5254 890 -5240
rect 856 -5308 890 -5292
rect 856 -5326 890 -5308
rect 856 -5376 890 -5364
rect 856 -5398 890 -5376
rect 856 -5444 890 -5436
rect 856 -5470 890 -5444
rect 856 -5512 890 -5508
rect 856 -5542 890 -5512
rect 5214 -5182 5248 -5172
rect 5214 -5240 5248 -5220
rect 5214 -5254 5248 -5240
rect 5214 -5308 5248 -5292
rect 5214 -5326 5248 -5308
rect 5214 -5376 5248 -5364
rect 5214 -5398 5248 -5376
rect 5214 -5444 5248 -5436
rect 5214 -5470 5248 -5444
rect 5214 -5512 5248 -5508
rect 5214 -5542 5248 -5512
rect 9573 -5182 9607 -5172
rect 9573 -5240 9607 -5220
rect 9573 -5254 9607 -5240
rect 9573 -5308 9607 -5292
rect 9573 -5326 9607 -5308
rect 9573 -5376 9607 -5364
rect 9573 -5398 9607 -5376
rect 9573 -5444 9607 -5436
rect 9573 -5470 9607 -5444
rect 9573 -5512 9607 -5508
rect 9573 -5542 9607 -5512
rect 13932 -5182 13966 -5172
rect 13932 -5240 13966 -5220
rect 13932 -5254 13966 -5240
rect 13932 -5308 13966 -5292
rect 13932 -5326 13966 -5308
rect 13932 -5376 13966 -5364
rect 13932 -5398 13966 -5376
rect 13932 -5444 13966 -5436
rect 13932 -5470 13966 -5444
rect 13932 -5512 13966 -5508
rect 13932 -5542 13966 -5512
rect 18290 -5182 18324 -5172
rect 18290 -5240 18324 -5220
rect 18290 -5254 18324 -5240
rect 18290 -5308 18324 -5292
rect 18290 -5326 18324 -5308
rect 18290 -5376 18324 -5364
rect 18290 -5398 18324 -5376
rect 18290 -5444 18324 -5436
rect 18290 -5470 18324 -5444
rect 18290 -5512 18324 -5508
rect 18290 -5542 18324 -5512
rect 856 -5614 890 -5580
rect 856 -5682 890 -5652
rect 856 -5686 890 -5682
rect 856 -5750 890 -5724
rect 856 -5758 890 -5750
rect 971 -5599 1005 -5597
rect 971 -5631 1005 -5599
rect 971 -5701 1005 -5669
rect 971 -5703 1005 -5701
rect 1229 -5599 1263 -5597
rect 1229 -5631 1263 -5599
rect 1229 -5701 1263 -5669
rect 1229 -5703 1263 -5701
rect 1423 -5599 1457 -5597
rect 1423 -5631 1457 -5599
rect 1423 -5701 1457 -5669
rect 1423 -5703 1457 -5701
rect 1681 -5599 1715 -5597
rect 1681 -5631 1715 -5599
rect 1681 -5701 1715 -5669
rect 1681 -5703 1715 -5701
rect 1939 -5599 1973 -5597
rect 1939 -5631 1973 -5599
rect 1939 -5701 1973 -5669
rect 1939 -5703 1973 -5701
rect 2197 -5599 2231 -5597
rect 2197 -5631 2231 -5599
rect 2197 -5701 2231 -5669
rect 2197 -5703 2231 -5701
rect 2455 -5599 2489 -5597
rect 2455 -5631 2489 -5599
rect 2455 -5701 2489 -5669
rect 2455 -5703 2489 -5701
rect 2649 -5599 2683 -5597
rect 2649 -5631 2683 -5599
rect 2649 -5701 2683 -5669
rect 2649 -5703 2683 -5701
rect 2907 -5599 2941 -5597
rect 2907 -5631 2941 -5599
rect 2907 -5701 2941 -5669
rect 2907 -5703 2941 -5701
rect 3165 -5599 3199 -5597
rect 3165 -5631 3199 -5599
rect 3165 -5701 3199 -5669
rect 3165 -5703 3199 -5701
rect 3423 -5599 3457 -5597
rect 3423 -5631 3457 -5599
rect 3423 -5701 3457 -5669
rect 3423 -5703 3457 -5701
rect 3617 -5599 3651 -5597
rect 3617 -5631 3651 -5599
rect 3617 -5701 3651 -5669
rect 3617 -5703 3651 -5701
rect 3875 -5599 3909 -5597
rect 3875 -5631 3909 -5599
rect 3875 -5701 3909 -5669
rect 3875 -5703 3909 -5701
rect 4133 -5599 4167 -5597
rect 4133 -5631 4167 -5599
rect 4133 -5701 4167 -5669
rect 4133 -5703 4167 -5701
rect 4391 -5599 4425 -5597
rect 4391 -5631 4425 -5599
rect 4391 -5701 4425 -5669
rect 4391 -5703 4425 -5701
rect 4649 -5599 4683 -5597
rect 4649 -5631 4683 -5599
rect 4649 -5701 4683 -5669
rect 4649 -5703 4683 -5701
rect 4842 -5599 4876 -5597
rect 4842 -5631 4876 -5599
rect 4842 -5701 4876 -5669
rect 4842 -5703 4876 -5701
rect 5100 -5599 5134 -5597
rect 5100 -5631 5134 -5599
rect 5100 -5701 5134 -5669
rect 5100 -5703 5134 -5701
rect 5214 -5614 5248 -5580
rect 5214 -5682 5248 -5652
rect 5214 -5686 5248 -5682
rect 5214 -5750 5248 -5724
rect 856 -5818 890 -5796
rect 5214 -5758 5248 -5750
rect 5328 -5599 5362 -5597
rect 5328 -5631 5362 -5599
rect 5328 -5701 5362 -5669
rect 5328 -5703 5362 -5701
rect 5586 -5599 5620 -5597
rect 5586 -5631 5620 -5599
rect 5586 -5701 5620 -5669
rect 5586 -5703 5620 -5701
rect 5780 -5599 5814 -5597
rect 5780 -5631 5814 -5599
rect 5780 -5701 5814 -5669
rect 5780 -5703 5814 -5701
rect 6038 -5599 6072 -5597
rect 6038 -5631 6072 -5599
rect 6038 -5701 6072 -5669
rect 6038 -5703 6072 -5701
rect 6296 -5599 6330 -5597
rect 6296 -5631 6330 -5599
rect 6296 -5701 6330 -5669
rect 6296 -5703 6330 -5701
rect 6554 -5599 6588 -5597
rect 6554 -5631 6588 -5599
rect 6554 -5701 6588 -5669
rect 6554 -5703 6588 -5701
rect 6812 -5599 6846 -5597
rect 6812 -5631 6846 -5599
rect 6812 -5701 6846 -5669
rect 6812 -5703 6846 -5701
rect 7006 -5599 7040 -5597
rect 7006 -5631 7040 -5599
rect 7006 -5701 7040 -5669
rect 7006 -5703 7040 -5701
rect 7264 -5599 7298 -5597
rect 7264 -5631 7298 -5599
rect 7264 -5701 7298 -5669
rect 7264 -5703 7298 -5701
rect 7522 -5599 7556 -5597
rect 7522 -5631 7556 -5599
rect 7522 -5701 7556 -5669
rect 7522 -5703 7556 -5701
rect 7780 -5599 7814 -5597
rect 7780 -5631 7814 -5599
rect 7780 -5701 7814 -5669
rect 7780 -5703 7814 -5701
rect 7974 -5599 8008 -5597
rect 7974 -5631 8008 -5599
rect 7974 -5701 8008 -5669
rect 7974 -5703 8008 -5701
rect 8232 -5599 8266 -5597
rect 8232 -5631 8266 -5599
rect 8232 -5701 8266 -5669
rect 8232 -5703 8266 -5701
rect 8490 -5599 8524 -5597
rect 8490 -5631 8524 -5599
rect 8490 -5701 8524 -5669
rect 8490 -5703 8524 -5701
rect 8748 -5599 8782 -5597
rect 8748 -5631 8782 -5599
rect 8748 -5701 8782 -5669
rect 8748 -5703 8782 -5701
rect 9006 -5599 9040 -5597
rect 9006 -5631 9040 -5599
rect 9006 -5701 9040 -5669
rect 9006 -5703 9040 -5701
rect 9200 -5599 9234 -5597
rect 9200 -5631 9234 -5599
rect 9200 -5701 9234 -5669
rect 9200 -5703 9234 -5701
rect 9458 -5599 9492 -5597
rect 9458 -5631 9492 -5599
rect 9458 -5701 9492 -5669
rect 9458 -5703 9492 -5701
rect 9573 -5614 9607 -5580
rect 9573 -5682 9607 -5652
rect 9573 -5686 9607 -5682
rect 9573 -5750 9607 -5724
rect 856 -5830 890 -5818
rect 1064 -5831 1066 -5797
rect 1066 -5831 1098 -5797
rect 1136 -5831 1168 -5797
rect 1168 -5831 1170 -5797
rect 1516 -5831 1518 -5797
rect 1518 -5831 1550 -5797
rect 1588 -5831 1620 -5797
rect 1620 -5831 1622 -5797
rect 1774 -5831 1776 -5797
rect 1776 -5831 1808 -5797
rect 1846 -5831 1878 -5797
rect 1878 -5831 1880 -5797
rect 2032 -5831 2034 -5797
rect 2034 -5831 2066 -5797
rect 2104 -5831 2136 -5797
rect 2136 -5831 2138 -5797
rect 2290 -5831 2292 -5797
rect 2292 -5831 2324 -5797
rect 2362 -5831 2394 -5797
rect 2394 -5831 2396 -5797
rect 2742 -5831 2744 -5797
rect 2744 -5831 2776 -5797
rect 2814 -5831 2846 -5797
rect 2846 -5831 2848 -5797
rect 3000 -5831 3002 -5797
rect 3002 -5831 3034 -5797
rect 3072 -5831 3104 -5797
rect 3104 -5831 3106 -5797
rect 3258 -5831 3260 -5797
rect 3260 -5831 3292 -5797
rect 3330 -5831 3362 -5797
rect 3362 -5831 3364 -5797
rect 3710 -5831 3712 -5797
rect 3712 -5831 3744 -5797
rect 3782 -5831 3814 -5797
rect 3814 -5831 3816 -5797
rect 3968 -5831 3970 -5797
rect 3970 -5831 4002 -5797
rect 4040 -5831 4072 -5797
rect 4072 -5831 4074 -5797
rect 4226 -5831 4228 -5797
rect 4228 -5831 4260 -5797
rect 4298 -5831 4330 -5797
rect 4330 -5831 4332 -5797
rect 4484 -5831 4486 -5797
rect 4486 -5831 4518 -5797
rect 4556 -5831 4588 -5797
rect 4588 -5831 4590 -5797
rect 4935 -5831 4937 -5797
rect 4937 -5831 4969 -5797
rect 5007 -5831 5039 -5797
rect 5039 -5831 5041 -5797
rect 5214 -5818 5248 -5796
rect 5214 -5830 5248 -5818
rect 9573 -5758 9607 -5750
rect 9688 -5599 9722 -5597
rect 9688 -5631 9722 -5599
rect 9688 -5701 9722 -5669
rect 9688 -5703 9722 -5701
rect 9946 -5599 9980 -5597
rect 9946 -5631 9980 -5599
rect 9946 -5701 9980 -5669
rect 9946 -5703 9980 -5701
rect 10140 -5599 10174 -5597
rect 10140 -5631 10174 -5599
rect 10140 -5701 10174 -5669
rect 10140 -5703 10174 -5701
rect 10398 -5599 10432 -5597
rect 10398 -5631 10432 -5599
rect 10398 -5701 10432 -5669
rect 10398 -5703 10432 -5701
rect 10656 -5599 10690 -5597
rect 10656 -5631 10690 -5599
rect 10656 -5701 10690 -5669
rect 10656 -5703 10690 -5701
rect 10914 -5599 10948 -5597
rect 10914 -5631 10948 -5599
rect 10914 -5701 10948 -5669
rect 10914 -5703 10948 -5701
rect 11172 -5599 11206 -5597
rect 11172 -5631 11206 -5599
rect 11172 -5701 11206 -5669
rect 11172 -5703 11206 -5701
rect 11366 -5599 11400 -5597
rect 11366 -5631 11400 -5599
rect 11366 -5701 11400 -5669
rect 11366 -5703 11400 -5701
rect 11624 -5599 11658 -5597
rect 11624 -5631 11658 -5599
rect 11624 -5701 11658 -5669
rect 11624 -5703 11658 -5701
rect 11882 -5599 11916 -5597
rect 11882 -5631 11916 -5599
rect 11882 -5701 11916 -5669
rect 11882 -5703 11916 -5701
rect 12140 -5599 12174 -5597
rect 12140 -5631 12174 -5599
rect 12140 -5701 12174 -5669
rect 12140 -5703 12174 -5701
rect 12334 -5599 12368 -5597
rect 12334 -5631 12368 -5599
rect 12334 -5701 12368 -5669
rect 12334 -5703 12368 -5701
rect 12592 -5599 12626 -5597
rect 12592 -5631 12626 -5599
rect 12592 -5701 12626 -5669
rect 12592 -5703 12626 -5701
rect 12850 -5599 12884 -5597
rect 12850 -5631 12884 -5599
rect 12850 -5701 12884 -5669
rect 12850 -5703 12884 -5701
rect 13108 -5599 13142 -5597
rect 13108 -5631 13142 -5599
rect 13108 -5701 13142 -5669
rect 13108 -5703 13142 -5701
rect 13366 -5599 13400 -5597
rect 13366 -5631 13400 -5599
rect 13366 -5701 13400 -5669
rect 13366 -5703 13400 -5701
rect 13560 -5599 13594 -5597
rect 13560 -5631 13594 -5599
rect 13560 -5701 13594 -5669
rect 13560 -5703 13594 -5701
rect 13818 -5599 13852 -5597
rect 13818 -5631 13852 -5599
rect 13818 -5701 13852 -5669
rect 13818 -5703 13852 -5701
rect 13932 -5614 13966 -5580
rect 13932 -5682 13966 -5652
rect 13932 -5686 13966 -5682
rect 856 -5886 890 -5868
rect 856 -5902 890 -5886
rect 856 -5954 890 -5940
rect 856 -5974 890 -5954
rect 856 -6022 890 -6012
rect 856 -6046 890 -6022
rect 856 -6090 890 -6084
rect 856 -6118 890 -6090
rect 856 -6158 890 -6156
rect 856 -6190 890 -6158
rect 5421 -5831 5423 -5797
rect 5423 -5831 5455 -5797
rect 5493 -5831 5525 -5797
rect 5525 -5831 5527 -5797
rect 5873 -5831 5875 -5797
rect 5875 -5831 5907 -5797
rect 5945 -5831 5977 -5797
rect 5977 -5831 5979 -5797
rect 6131 -5831 6133 -5797
rect 6133 -5831 6165 -5797
rect 6203 -5831 6235 -5797
rect 6235 -5831 6237 -5797
rect 6389 -5831 6391 -5797
rect 6391 -5831 6423 -5797
rect 6461 -5831 6493 -5797
rect 6493 -5831 6495 -5797
rect 6647 -5831 6649 -5797
rect 6649 -5831 6681 -5797
rect 6719 -5831 6751 -5797
rect 6751 -5831 6753 -5797
rect 7099 -5831 7101 -5797
rect 7101 -5831 7133 -5797
rect 7171 -5831 7203 -5797
rect 7203 -5831 7205 -5797
rect 7357 -5831 7359 -5797
rect 7359 -5831 7391 -5797
rect 7429 -5831 7461 -5797
rect 7461 -5831 7463 -5797
rect 7615 -5831 7617 -5797
rect 7617 -5831 7649 -5797
rect 7687 -5831 7719 -5797
rect 7719 -5831 7721 -5797
rect 8067 -5831 8069 -5797
rect 8069 -5831 8101 -5797
rect 8139 -5831 8171 -5797
rect 8171 -5831 8173 -5797
rect 8325 -5831 8327 -5797
rect 8327 -5831 8359 -5797
rect 8397 -5831 8429 -5797
rect 8429 -5831 8431 -5797
rect 8583 -5831 8585 -5797
rect 8585 -5831 8617 -5797
rect 8655 -5831 8687 -5797
rect 8687 -5831 8689 -5797
rect 8841 -5831 8843 -5797
rect 8843 -5831 8875 -5797
rect 8913 -5831 8945 -5797
rect 8945 -5831 8947 -5797
rect 9293 -5831 9295 -5797
rect 9295 -5831 9327 -5797
rect 9365 -5831 9397 -5797
rect 9397 -5831 9399 -5797
rect 9573 -5818 9607 -5796
rect 13932 -5750 13966 -5724
rect 13932 -5758 13966 -5750
rect 14046 -5599 14080 -5597
rect 14046 -5631 14080 -5599
rect 14046 -5701 14080 -5669
rect 14046 -5703 14080 -5701
rect 14304 -5599 14338 -5597
rect 14304 -5631 14338 -5599
rect 14304 -5701 14338 -5669
rect 14304 -5703 14338 -5701
rect 14497 -5599 14531 -5597
rect 14497 -5631 14531 -5599
rect 14497 -5701 14531 -5669
rect 14497 -5703 14531 -5701
rect 14755 -5599 14789 -5597
rect 14755 -5631 14789 -5599
rect 14755 -5701 14789 -5669
rect 14755 -5703 14789 -5701
rect 15013 -5599 15047 -5597
rect 15013 -5631 15047 -5599
rect 15013 -5701 15047 -5669
rect 15013 -5703 15047 -5701
rect 15271 -5599 15305 -5597
rect 15271 -5631 15305 -5599
rect 15271 -5701 15305 -5669
rect 15271 -5703 15305 -5701
rect 15529 -5599 15563 -5597
rect 15529 -5631 15563 -5599
rect 15529 -5701 15563 -5669
rect 15529 -5703 15563 -5701
rect 15723 -5599 15757 -5597
rect 15723 -5631 15757 -5599
rect 15723 -5701 15757 -5669
rect 15723 -5703 15757 -5701
rect 15981 -5599 16015 -5597
rect 15981 -5631 16015 -5599
rect 15981 -5701 16015 -5669
rect 15981 -5703 16015 -5701
rect 16239 -5599 16273 -5597
rect 16239 -5631 16273 -5599
rect 16239 -5701 16273 -5669
rect 16239 -5703 16273 -5701
rect 16497 -5599 16531 -5597
rect 16497 -5631 16531 -5599
rect 16497 -5701 16531 -5669
rect 16497 -5703 16531 -5701
rect 16691 -5599 16725 -5597
rect 16691 -5631 16725 -5599
rect 16691 -5701 16725 -5669
rect 16691 -5703 16725 -5701
rect 16949 -5599 16983 -5597
rect 16949 -5631 16983 -5599
rect 16949 -5701 16983 -5669
rect 16949 -5703 16983 -5701
rect 17207 -5599 17241 -5597
rect 17207 -5631 17241 -5599
rect 17207 -5701 17241 -5669
rect 17207 -5703 17241 -5701
rect 17465 -5599 17499 -5597
rect 17465 -5631 17499 -5599
rect 17465 -5701 17499 -5669
rect 17465 -5703 17499 -5701
rect 17723 -5599 17757 -5597
rect 17723 -5631 17757 -5599
rect 17723 -5701 17757 -5669
rect 17723 -5703 17757 -5701
rect 17917 -5599 17951 -5597
rect 17917 -5631 17951 -5599
rect 17917 -5701 17951 -5669
rect 17917 -5703 17951 -5701
rect 18175 -5599 18209 -5597
rect 18175 -5631 18209 -5599
rect 18175 -5701 18209 -5669
rect 18175 -5703 18209 -5701
rect 18290 -5614 18324 -5580
rect 18290 -5682 18324 -5652
rect 18290 -5686 18324 -5682
rect 18290 -5750 18324 -5724
rect 9573 -5830 9607 -5818
rect 5214 -5886 5248 -5868
rect 5214 -5902 5248 -5886
rect 5214 -5954 5248 -5940
rect 5214 -5974 5248 -5954
rect 5214 -6022 5248 -6012
rect 5214 -6046 5248 -6022
rect 5214 -6090 5248 -6084
rect 5214 -6118 5248 -6090
rect 5214 -6158 5248 -6156
rect 1064 -6193 1066 -6159
rect 1066 -6193 1098 -6159
rect 1136 -6193 1168 -6159
rect 1168 -6193 1170 -6159
rect 1516 -6193 1518 -6159
rect 1518 -6193 1550 -6159
rect 1588 -6193 1620 -6159
rect 1620 -6193 1622 -6159
rect 1774 -6193 1776 -6159
rect 1776 -6193 1808 -6159
rect 1846 -6193 1878 -6159
rect 1878 -6193 1880 -6159
rect 2032 -6193 2034 -6159
rect 2034 -6193 2066 -6159
rect 2104 -6193 2136 -6159
rect 2136 -6193 2138 -6159
rect 2290 -6193 2292 -6159
rect 2292 -6193 2324 -6159
rect 2362 -6193 2394 -6159
rect 2394 -6193 2396 -6159
rect 2742 -6193 2744 -6159
rect 2744 -6193 2776 -6159
rect 2814 -6193 2846 -6159
rect 2846 -6193 2848 -6159
rect 3000 -6193 3002 -6159
rect 3002 -6193 3034 -6159
rect 3072 -6193 3104 -6159
rect 3104 -6193 3106 -6159
rect 3258 -6193 3260 -6159
rect 3260 -6193 3292 -6159
rect 3330 -6193 3362 -6159
rect 3362 -6193 3364 -6159
rect 3710 -6193 3712 -6159
rect 3712 -6193 3744 -6159
rect 3782 -6193 3814 -6159
rect 3814 -6193 3816 -6159
rect 3968 -6193 3970 -6159
rect 3970 -6193 4002 -6159
rect 4040 -6193 4072 -6159
rect 4072 -6193 4074 -6159
rect 4226 -6193 4228 -6159
rect 4228 -6193 4260 -6159
rect 4298 -6193 4330 -6159
rect 4330 -6193 4332 -6159
rect 4484 -6193 4486 -6159
rect 4486 -6193 4518 -6159
rect 4556 -6193 4588 -6159
rect 4588 -6193 4590 -6159
rect 4935 -6193 4937 -6159
rect 4937 -6193 4969 -6159
rect 5007 -6193 5039 -6159
rect 5039 -6193 5041 -6159
rect 5214 -6190 5248 -6158
rect 9781 -5831 9783 -5797
rect 9783 -5831 9815 -5797
rect 9853 -5831 9885 -5797
rect 9885 -5831 9887 -5797
rect 10233 -5831 10235 -5797
rect 10235 -5831 10267 -5797
rect 10305 -5831 10337 -5797
rect 10337 -5831 10339 -5797
rect 10491 -5831 10493 -5797
rect 10493 -5831 10525 -5797
rect 10563 -5831 10595 -5797
rect 10595 -5831 10597 -5797
rect 10749 -5831 10751 -5797
rect 10751 -5831 10783 -5797
rect 10821 -5831 10853 -5797
rect 10853 -5831 10855 -5797
rect 11007 -5831 11009 -5797
rect 11009 -5831 11041 -5797
rect 11079 -5831 11111 -5797
rect 11111 -5831 11113 -5797
rect 11459 -5831 11461 -5797
rect 11461 -5831 11493 -5797
rect 11531 -5831 11563 -5797
rect 11563 -5831 11565 -5797
rect 11717 -5831 11719 -5797
rect 11719 -5831 11751 -5797
rect 11789 -5831 11821 -5797
rect 11821 -5831 11823 -5797
rect 11975 -5831 11977 -5797
rect 11977 -5831 12009 -5797
rect 12047 -5831 12079 -5797
rect 12079 -5831 12081 -5797
rect 12427 -5831 12429 -5797
rect 12429 -5831 12461 -5797
rect 12499 -5831 12531 -5797
rect 12531 -5831 12533 -5797
rect 12685 -5831 12687 -5797
rect 12687 -5831 12719 -5797
rect 12757 -5831 12789 -5797
rect 12789 -5831 12791 -5797
rect 12943 -5831 12945 -5797
rect 12945 -5831 12977 -5797
rect 13015 -5831 13047 -5797
rect 13047 -5831 13049 -5797
rect 13201 -5831 13203 -5797
rect 13203 -5831 13235 -5797
rect 13273 -5831 13305 -5797
rect 13305 -5831 13307 -5797
rect 13653 -5831 13655 -5797
rect 13655 -5831 13687 -5797
rect 13725 -5831 13757 -5797
rect 13757 -5831 13759 -5797
rect 13932 -5818 13966 -5796
rect 18290 -5758 18324 -5750
rect 13932 -5830 13966 -5818
rect 9573 -5886 9607 -5868
rect 9573 -5902 9607 -5886
rect 9573 -5954 9607 -5940
rect 9573 -5974 9607 -5954
rect 9573 -6022 9607 -6012
rect 9573 -6046 9607 -6022
rect 9573 -6090 9607 -6084
rect 9573 -6118 9607 -6090
rect 9573 -6158 9607 -6156
rect 856 -6260 890 -6228
rect 5421 -6193 5423 -6159
rect 5423 -6193 5455 -6159
rect 5493 -6193 5525 -6159
rect 5525 -6193 5527 -6159
rect 5873 -6193 5875 -6159
rect 5875 -6193 5907 -6159
rect 5945 -6193 5977 -6159
rect 5977 -6193 5979 -6159
rect 6131 -6193 6133 -6159
rect 6133 -6193 6165 -6159
rect 6203 -6193 6235 -6159
rect 6235 -6193 6237 -6159
rect 6389 -6193 6391 -6159
rect 6391 -6193 6423 -6159
rect 6461 -6193 6493 -6159
rect 6493 -6193 6495 -6159
rect 6647 -6193 6649 -6159
rect 6649 -6193 6681 -6159
rect 6719 -6193 6751 -6159
rect 6751 -6193 6753 -6159
rect 7099 -6193 7101 -6159
rect 7101 -6193 7133 -6159
rect 7171 -6193 7203 -6159
rect 7203 -6193 7205 -6159
rect 7357 -6193 7359 -6159
rect 7359 -6193 7391 -6159
rect 7429 -6193 7461 -6159
rect 7461 -6193 7463 -6159
rect 7615 -6193 7617 -6159
rect 7617 -6193 7649 -6159
rect 7687 -6193 7719 -6159
rect 7719 -6193 7721 -6159
rect 8067 -6193 8069 -6159
rect 8069 -6193 8101 -6159
rect 8139 -6193 8171 -6159
rect 8171 -6193 8173 -6159
rect 8325 -6193 8327 -6159
rect 8327 -6193 8359 -6159
rect 8397 -6193 8429 -6159
rect 8429 -6193 8431 -6159
rect 8583 -6193 8585 -6159
rect 8585 -6193 8617 -6159
rect 8655 -6193 8687 -6159
rect 8687 -6193 8689 -6159
rect 8841 -6193 8843 -6159
rect 8843 -6193 8875 -6159
rect 8913 -6193 8945 -6159
rect 8945 -6193 8947 -6159
rect 9293 -6193 9295 -6159
rect 9295 -6193 9327 -6159
rect 9365 -6193 9397 -6159
rect 9397 -6193 9399 -6159
rect 9573 -6190 9607 -6158
rect 14139 -5831 14141 -5797
rect 14141 -5831 14173 -5797
rect 14211 -5831 14243 -5797
rect 14243 -5831 14245 -5797
rect 14590 -5831 14592 -5797
rect 14592 -5831 14624 -5797
rect 14662 -5831 14694 -5797
rect 14694 -5831 14696 -5797
rect 14848 -5831 14850 -5797
rect 14850 -5831 14882 -5797
rect 14920 -5831 14952 -5797
rect 14952 -5831 14954 -5797
rect 15106 -5831 15108 -5797
rect 15108 -5831 15140 -5797
rect 15178 -5831 15210 -5797
rect 15210 -5831 15212 -5797
rect 15364 -5831 15366 -5797
rect 15366 -5831 15398 -5797
rect 15436 -5831 15468 -5797
rect 15468 -5831 15470 -5797
rect 15816 -5831 15818 -5797
rect 15818 -5831 15850 -5797
rect 15888 -5831 15920 -5797
rect 15920 -5831 15922 -5797
rect 16074 -5831 16076 -5797
rect 16076 -5831 16108 -5797
rect 16146 -5831 16178 -5797
rect 16178 -5831 16180 -5797
rect 16332 -5831 16334 -5797
rect 16334 -5831 16366 -5797
rect 16404 -5831 16436 -5797
rect 16436 -5831 16438 -5797
rect 16784 -5831 16786 -5797
rect 16786 -5831 16818 -5797
rect 16856 -5831 16888 -5797
rect 16888 -5831 16890 -5797
rect 17042 -5831 17044 -5797
rect 17044 -5831 17076 -5797
rect 17114 -5831 17146 -5797
rect 17146 -5831 17148 -5797
rect 17300 -5831 17302 -5797
rect 17302 -5831 17334 -5797
rect 17372 -5831 17404 -5797
rect 17404 -5831 17406 -5797
rect 17558 -5831 17560 -5797
rect 17560 -5831 17592 -5797
rect 17630 -5831 17662 -5797
rect 17662 -5831 17664 -5797
rect 18010 -5831 18012 -5797
rect 18012 -5831 18044 -5797
rect 18082 -5831 18114 -5797
rect 18114 -5831 18116 -5797
rect 18290 -5818 18324 -5796
rect 18290 -5830 18324 -5818
rect 13932 -5886 13966 -5868
rect 13932 -5902 13966 -5886
rect 13932 -5954 13966 -5940
rect 13932 -5974 13966 -5954
rect 13932 -6022 13966 -6012
rect 13932 -6046 13966 -6022
rect 13932 -6090 13966 -6084
rect 13932 -6118 13966 -6090
rect 856 -6262 890 -6260
rect 856 -6328 890 -6300
rect 856 -6334 890 -6328
rect 856 -6396 890 -6372
rect 856 -6406 890 -6396
rect 971 -6289 1005 -6287
rect 971 -6321 1005 -6289
rect 971 -6391 1005 -6359
rect 971 -6393 1005 -6391
rect 1229 -6289 1263 -6287
rect 1229 -6321 1263 -6289
rect 1229 -6391 1263 -6359
rect 1229 -6393 1263 -6391
rect 1423 -6289 1457 -6287
rect 1423 -6321 1457 -6289
rect 1423 -6391 1457 -6359
rect 1423 -6393 1457 -6391
rect 1681 -6289 1715 -6287
rect 1681 -6321 1715 -6289
rect 1681 -6391 1715 -6359
rect 1681 -6393 1715 -6391
rect 1939 -6289 1973 -6287
rect 1939 -6321 1973 -6289
rect 1939 -6391 1973 -6359
rect 1939 -6393 1973 -6391
rect 2197 -6289 2231 -6287
rect 2197 -6321 2231 -6289
rect 2197 -6391 2231 -6359
rect 2197 -6393 2231 -6391
rect 2455 -6289 2489 -6287
rect 2455 -6321 2489 -6289
rect 2455 -6391 2489 -6359
rect 2455 -6393 2489 -6391
rect 2649 -6289 2683 -6287
rect 2649 -6321 2683 -6289
rect 2649 -6391 2683 -6359
rect 2649 -6393 2683 -6391
rect 2907 -6289 2941 -6287
rect 2907 -6321 2941 -6289
rect 2907 -6391 2941 -6359
rect 2907 -6393 2941 -6391
rect 3165 -6289 3199 -6287
rect 3165 -6321 3199 -6289
rect 3165 -6391 3199 -6359
rect 3165 -6393 3199 -6391
rect 3423 -6289 3457 -6287
rect 3423 -6321 3457 -6289
rect 3423 -6391 3457 -6359
rect 3423 -6393 3457 -6391
rect 3617 -6289 3651 -6287
rect 3617 -6321 3651 -6289
rect 3617 -6391 3651 -6359
rect 3617 -6393 3651 -6391
rect 3875 -6289 3909 -6287
rect 3875 -6321 3909 -6289
rect 3875 -6391 3909 -6359
rect 3875 -6393 3909 -6391
rect 4133 -6289 4167 -6287
rect 4133 -6321 4167 -6289
rect 4133 -6391 4167 -6359
rect 4133 -6393 4167 -6391
rect 4391 -6289 4425 -6287
rect 4391 -6321 4425 -6289
rect 4391 -6391 4425 -6359
rect 4391 -6393 4425 -6391
rect 4649 -6289 4683 -6287
rect 4649 -6321 4683 -6289
rect 4649 -6391 4683 -6359
rect 4649 -6393 4683 -6391
rect 4842 -6289 4876 -6287
rect 4842 -6321 4876 -6289
rect 4842 -6391 4876 -6359
rect 4842 -6393 4876 -6391
rect 5100 -6289 5134 -6287
rect 5100 -6321 5134 -6289
rect 5100 -6391 5134 -6359
rect 5100 -6393 5134 -6391
rect 5214 -6260 5248 -6228
rect 5214 -6262 5248 -6260
rect 9781 -6193 9783 -6159
rect 9783 -6193 9815 -6159
rect 9853 -6193 9885 -6159
rect 9885 -6193 9887 -6159
rect 10233 -6193 10235 -6159
rect 10235 -6193 10267 -6159
rect 10305 -6193 10337 -6159
rect 10337 -6193 10339 -6159
rect 10491 -6193 10493 -6159
rect 10493 -6193 10525 -6159
rect 10563 -6193 10595 -6159
rect 10595 -6193 10597 -6159
rect 10749 -6193 10751 -6159
rect 10751 -6193 10783 -6159
rect 10821 -6193 10853 -6159
rect 10853 -6193 10855 -6159
rect 11007 -6193 11009 -6159
rect 11009 -6193 11041 -6159
rect 11079 -6193 11111 -6159
rect 11111 -6193 11113 -6159
rect 11459 -6193 11461 -6159
rect 11461 -6193 11493 -6159
rect 11531 -6193 11563 -6159
rect 11563 -6193 11565 -6159
rect 11717 -6193 11719 -6159
rect 11719 -6193 11751 -6159
rect 11789 -6193 11821 -6159
rect 11821 -6193 11823 -6159
rect 11975 -6193 11977 -6159
rect 11977 -6193 12009 -6159
rect 12047 -6193 12079 -6159
rect 12079 -6193 12081 -6159
rect 12427 -6193 12429 -6159
rect 12429 -6193 12461 -6159
rect 12499 -6193 12531 -6159
rect 12531 -6193 12533 -6159
rect 12685 -6193 12687 -6159
rect 12687 -6193 12719 -6159
rect 12757 -6193 12789 -6159
rect 12789 -6193 12791 -6159
rect 12943 -6193 12945 -6159
rect 12945 -6193 12977 -6159
rect 13015 -6193 13047 -6159
rect 13047 -6193 13049 -6159
rect 13201 -6193 13203 -6159
rect 13203 -6193 13235 -6159
rect 13273 -6193 13305 -6159
rect 13305 -6193 13307 -6159
rect 13653 -6193 13655 -6159
rect 13655 -6193 13687 -6159
rect 13725 -6193 13757 -6159
rect 13757 -6193 13759 -6159
rect 13932 -6158 13966 -6156
rect 13932 -6190 13966 -6158
rect 18290 -5886 18324 -5868
rect 18290 -5902 18324 -5886
rect 18290 -5954 18324 -5940
rect 18290 -5974 18324 -5954
rect 18290 -6022 18324 -6012
rect 18290 -6046 18324 -6022
rect 18290 -6090 18324 -6084
rect 18290 -6118 18324 -6090
rect 18290 -6158 18324 -6156
rect 5214 -6328 5248 -6300
rect 5214 -6334 5248 -6328
rect 5214 -6396 5248 -6372
rect 5214 -6406 5248 -6396
rect 5328 -6289 5362 -6287
rect 5328 -6321 5362 -6289
rect 5328 -6391 5362 -6359
rect 5328 -6393 5362 -6391
rect 5586 -6289 5620 -6287
rect 5586 -6321 5620 -6289
rect 5586 -6391 5620 -6359
rect 5586 -6393 5620 -6391
rect 5780 -6289 5814 -6287
rect 5780 -6321 5814 -6289
rect 5780 -6391 5814 -6359
rect 5780 -6393 5814 -6391
rect 6038 -6289 6072 -6287
rect 6038 -6321 6072 -6289
rect 6038 -6391 6072 -6359
rect 6038 -6393 6072 -6391
rect 6296 -6289 6330 -6287
rect 6296 -6321 6330 -6289
rect 6296 -6391 6330 -6359
rect 6296 -6393 6330 -6391
rect 6554 -6289 6588 -6287
rect 6554 -6321 6588 -6289
rect 6554 -6391 6588 -6359
rect 6554 -6393 6588 -6391
rect 6812 -6289 6846 -6287
rect 6812 -6321 6846 -6289
rect 6812 -6391 6846 -6359
rect 6812 -6393 6846 -6391
rect 7006 -6289 7040 -6287
rect 7006 -6321 7040 -6289
rect 7006 -6391 7040 -6359
rect 7006 -6393 7040 -6391
rect 7264 -6289 7298 -6287
rect 7264 -6321 7298 -6289
rect 7264 -6391 7298 -6359
rect 7264 -6393 7298 -6391
rect 7522 -6289 7556 -6287
rect 7522 -6321 7556 -6289
rect 7522 -6391 7556 -6359
rect 7522 -6393 7556 -6391
rect 7780 -6289 7814 -6287
rect 7780 -6321 7814 -6289
rect 7780 -6391 7814 -6359
rect 7780 -6393 7814 -6391
rect 7974 -6289 8008 -6287
rect 7974 -6321 8008 -6289
rect 7974 -6391 8008 -6359
rect 7974 -6393 8008 -6391
rect 8232 -6289 8266 -6287
rect 8232 -6321 8266 -6289
rect 8232 -6391 8266 -6359
rect 8232 -6393 8266 -6391
rect 8490 -6289 8524 -6287
rect 8490 -6321 8524 -6289
rect 8490 -6391 8524 -6359
rect 8490 -6393 8524 -6391
rect 8748 -6289 8782 -6287
rect 8748 -6321 8782 -6289
rect 8748 -6391 8782 -6359
rect 8748 -6393 8782 -6391
rect 9006 -6289 9040 -6287
rect 9006 -6321 9040 -6289
rect 9006 -6391 9040 -6359
rect 9006 -6393 9040 -6391
rect 9200 -6289 9234 -6287
rect 9200 -6321 9234 -6289
rect 9200 -6391 9234 -6359
rect 9200 -6393 9234 -6391
rect 9458 -6289 9492 -6287
rect 9458 -6321 9492 -6289
rect 9458 -6391 9492 -6359
rect 9458 -6393 9492 -6391
rect 9573 -6260 9607 -6228
rect 14139 -6193 14141 -6159
rect 14141 -6193 14173 -6159
rect 14211 -6193 14243 -6159
rect 14243 -6193 14245 -6159
rect 14590 -6193 14592 -6159
rect 14592 -6193 14624 -6159
rect 14662 -6193 14694 -6159
rect 14694 -6193 14696 -6159
rect 14848 -6193 14850 -6159
rect 14850 -6193 14882 -6159
rect 14920 -6193 14952 -6159
rect 14952 -6193 14954 -6159
rect 15106 -6193 15108 -6159
rect 15108 -6193 15140 -6159
rect 15178 -6193 15210 -6159
rect 15210 -6193 15212 -6159
rect 15364 -6193 15366 -6159
rect 15366 -6193 15398 -6159
rect 15436 -6193 15468 -6159
rect 15468 -6193 15470 -6159
rect 15816 -6193 15818 -6159
rect 15818 -6193 15850 -6159
rect 15888 -6193 15920 -6159
rect 15920 -6193 15922 -6159
rect 16074 -6193 16076 -6159
rect 16076 -6193 16108 -6159
rect 16146 -6193 16178 -6159
rect 16178 -6193 16180 -6159
rect 16332 -6193 16334 -6159
rect 16334 -6193 16366 -6159
rect 16404 -6193 16436 -6159
rect 16436 -6193 16438 -6159
rect 16784 -6193 16786 -6159
rect 16786 -6193 16818 -6159
rect 16856 -6193 16888 -6159
rect 16888 -6193 16890 -6159
rect 17042 -6193 17044 -6159
rect 17044 -6193 17076 -6159
rect 17114 -6193 17146 -6159
rect 17146 -6193 17148 -6159
rect 17300 -6193 17302 -6159
rect 17302 -6193 17334 -6159
rect 17372 -6193 17404 -6159
rect 17404 -6193 17406 -6159
rect 17558 -6193 17560 -6159
rect 17560 -6193 17592 -6159
rect 17630 -6193 17662 -6159
rect 17662 -6193 17664 -6159
rect 18010 -6193 18012 -6159
rect 18012 -6193 18044 -6159
rect 18082 -6193 18114 -6159
rect 18114 -6193 18116 -6159
rect 18290 -6190 18324 -6158
rect 9573 -6262 9607 -6260
rect 9573 -6328 9607 -6300
rect 9573 -6334 9607 -6328
rect 9573 -6396 9607 -6372
rect 9573 -6406 9607 -6396
rect 9688 -6289 9722 -6287
rect 9688 -6321 9722 -6289
rect 9688 -6391 9722 -6359
rect 9688 -6393 9722 -6391
rect 9946 -6289 9980 -6287
rect 9946 -6321 9980 -6289
rect 9946 -6391 9980 -6359
rect 9946 -6393 9980 -6391
rect 10140 -6289 10174 -6287
rect 10140 -6321 10174 -6289
rect 10140 -6391 10174 -6359
rect 10140 -6393 10174 -6391
rect 10398 -6289 10432 -6287
rect 10398 -6321 10432 -6289
rect 10398 -6391 10432 -6359
rect 10398 -6393 10432 -6391
rect 10656 -6289 10690 -6287
rect 10656 -6321 10690 -6289
rect 10656 -6391 10690 -6359
rect 10656 -6393 10690 -6391
rect 10914 -6289 10948 -6287
rect 10914 -6321 10948 -6289
rect 10914 -6391 10948 -6359
rect 10914 -6393 10948 -6391
rect 11172 -6289 11206 -6287
rect 11172 -6321 11206 -6289
rect 11172 -6391 11206 -6359
rect 11172 -6393 11206 -6391
rect 11366 -6289 11400 -6287
rect 11366 -6321 11400 -6289
rect 11366 -6391 11400 -6359
rect 11366 -6393 11400 -6391
rect 11624 -6289 11658 -6287
rect 11624 -6321 11658 -6289
rect 11624 -6391 11658 -6359
rect 11624 -6393 11658 -6391
rect 11882 -6289 11916 -6287
rect 11882 -6321 11916 -6289
rect 11882 -6391 11916 -6359
rect 11882 -6393 11916 -6391
rect 12140 -6289 12174 -6287
rect 12140 -6321 12174 -6289
rect 12140 -6391 12174 -6359
rect 12140 -6393 12174 -6391
rect 12334 -6289 12368 -6287
rect 12334 -6321 12368 -6289
rect 12334 -6391 12368 -6359
rect 12334 -6393 12368 -6391
rect 12592 -6289 12626 -6287
rect 12592 -6321 12626 -6289
rect 12592 -6391 12626 -6359
rect 12592 -6393 12626 -6391
rect 12850 -6289 12884 -6287
rect 12850 -6321 12884 -6289
rect 12850 -6391 12884 -6359
rect 12850 -6393 12884 -6391
rect 13108 -6289 13142 -6287
rect 13108 -6321 13142 -6289
rect 13108 -6391 13142 -6359
rect 13108 -6393 13142 -6391
rect 13366 -6289 13400 -6287
rect 13366 -6321 13400 -6289
rect 13366 -6391 13400 -6359
rect 13366 -6393 13400 -6391
rect 13560 -6289 13594 -6287
rect 13560 -6321 13594 -6289
rect 13560 -6391 13594 -6359
rect 13560 -6393 13594 -6391
rect 13818 -6289 13852 -6287
rect 13818 -6321 13852 -6289
rect 13818 -6391 13852 -6359
rect 13818 -6393 13852 -6391
rect 13932 -6260 13966 -6228
rect 13932 -6262 13966 -6260
rect 13932 -6328 13966 -6300
rect 13932 -6334 13966 -6328
rect 13932 -6396 13966 -6372
rect 13932 -6406 13966 -6396
rect 14046 -6289 14080 -6287
rect 14046 -6321 14080 -6289
rect 14046 -6391 14080 -6359
rect 14046 -6393 14080 -6391
rect 14304 -6289 14338 -6287
rect 14304 -6321 14338 -6289
rect 14304 -6391 14338 -6359
rect 14304 -6393 14338 -6391
rect 14497 -6289 14531 -6287
rect 14497 -6321 14531 -6289
rect 14497 -6391 14531 -6359
rect 14497 -6393 14531 -6391
rect 14755 -6289 14789 -6287
rect 14755 -6321 14789 -6289
rect 14755 -6391 14789 -6359
rect 14755 -6393 14789 -6391
rect 15013 -6289 15047 -6287
rect 15013 -6321 15047 -6289
rect 15013 -6391 15047 -6359
rect 15013 -6393 15047 -6391
rect 15271 -6289 15305 -6287
rect 15271 -6321 15305 -6289
rect 15271 -6391 15305 -6359
rect 15271 -6393 15305 -6391
rect 15529 -6289 15563 -6287
rect 15529 -6321 15563 -6289
rect 15529 -6391 15563 -6359
rect 15529 -6393 15563 -6391
rect 15723 -6289 15757 -6287
rect 15723 -6321 15757 -6289
rect 15723 -6391 15757 -6359
rect 15723 -6393 15757 -6391
rect 15981 -6289 16015 -6287
rect 15981 -6321 16015 -6289
rect 15981 -6391 16015 -6359
rect 15981 -6393 16015 -6391
rect 16239 -6289 16273 -6287
rect 16239 -6321 16273 -6289
rect 16239 -6391 16273 -6359
rect 16239 -6393 16273 -6391
rect 16497 -6289 16531 -6287
rect 16497 -6321 16531 -6289
rect 16497 -6391 16531 -6359
rect 16497 -6393 16531 -6391
rect 16691 -6289 16725 -6287
rect 16691 -6321 16725 -6289
rect 16691 -6391 16725 -6359
rect 16691 -6393 16725 -6391
rect 16949 -6289 16983 -6287
rect 16949 -6321 16983 -6289
rect 16949 -6391 16983 -6359
rect 16949 -6393 16983 -6391
rect 17207 -6289 17241 -6287
rect 17207 -6321 17241 -6289
rect 17207 -6391 17241 -6359
rect 17207 -6393 17241 -6391
rect 17465 -6289 17499 -6287
rect 17465 -6321 17499 -6289
rect 17465 -6391 17499 -6359
rect 17465 -6393 17499 -6391
rect 17723 -6289 17757 -6287
rect 17723 -6321 17757 -6289
rect 17723 -6391 17757 -6359
rect 17723 -6393 17757 -6391
rect 17917 -6289 17951 -6287
rect 17917 -6321 17951 -6289
rect 17917 -6391 17951 -6359
rect 17917 -6393 17951 -6391
rect 18175 -6289 18209 -6287
rect 18175 -6321 18209 -6289
rect 18175 -6391 18209 -6359
rect 18175 -6393 18209 -6391
rect 18290 -6260 18324 -6228
rect 18290 -6262 18324 -6260
rect 18290 -6328 18324 -6300
rect 18290 -6334 18324 -6328
rect 18290 -6396 18324 -6372
rect 18290 -6406 18324 -6396
rect 856 -6464 890 -6444
rect 856 -6478 890 -6464
rect 856 -6532 890 -6516
rect 856 -6550 890 -6532
rect 856 -6600 890 -6588
rect 856 -6622 890 -6600
rect 856 -6668 890 -6660
rect 856 -6694 890 -6668
rect 856 -6766 890 -6732
rect 5214 -6464 5248 -6444
rect 5214 -6478 5248 -6464
rect 5214 -6532 5248 -6516
rect 5214 -6550 5248 -6532
rect 5214 -6600 5248 -6588
rect 5214 -6622 5248 -6600
rect 5214 -6668 5248 -6660
rect 5214 -6694 5248 -6668
rect 5214 -6766 5248 -6732
rect 9573 -6464 9607 -6444
rect 9573 -6478 9607 -6464
rect 9573 -6532 9607 -6516
rect 9573 -6550 9607 -6532
rect 9573 -6600 9607 -6588
rect 9573 -6622 9607 -6600
rect 9573 -6668 9607 -6660
rect 9573 -6694 9607 -6668
rect 9573 -6766 9607 -6732
rect 13932 -6464 13966 -6444
rect 13932 -6478 13966 -6464
rect 13932 -6532 13966 -6516
rect 13932 -6550 13966 -6532
rect 13932 -6600 13966 -6588
rect 13932 -6622 13966 -6600
rect 13932 -6668 13966 -6660
rect 13932 -6694 13966 -6668
rect 13932 -6766 13966 -6732
rect 18290 -6464 18324 -6444
rect 18290 -6478 18324 -6464
rect 18290 -6532 18324 -6516
rect 18290 -6550 18324 -6532
rect 18290 -6600 18324 -6588
rect 18290 -6622 18324 -6600
rect 18290 -6668 18324 -6660
rect 18290 -6694 18324 -6668
rect 18290 -6766 18324 -6732
rect 856 -6838 890 -6804
rect 5214 -6838 5248 -6804
rect 9573 -6838 9607 -6804
rect 13932 -6838 13966 -6804
rect 18290 -6838 18324 -6804
rect 856 -6910 890 -6876
rect 856 -6974 890 -6948
rect 856 -6982 890 -6974
rect 856 -7042 890 -7020
rect 856 -7054 890 -7042
rect 856 -7110 890 -7092
rect 856 -7126 890 -7110
rect 856 -7178 890 -7164
rect 856 -7198 890 -7178
rect 5214 -6910 5248 -6876
rect 5214 -6974 5248 -6948
rect 5214 -6982 5248 -6974
rect 5214 -7042 5248 -7020
rect 5214 -7054 5248 -7042
rect 5214 -7110 5248 -7092
rect 5214 -7126 5248 -7110
rect 5214 -7178 5248 -7164
rect 856 -7246 890 -7236
rect 856 -7270 890 -7246
rect 856 -7314 890 -7308
rect 856 -7342 890 -7314
rect 856 -7382 890 -7380
rect 856 -7414 890 -7382
rect 971 -7246 1005 -7244
rect 971 -7278 1005 -7246
rect 971 -7348 1005 -7316
rect 971 -7350 1005 -7348
rect 1229 -7246 1263 -7244
rect 1229 -7278 1263 -7246
rect 1229 -7348 1263 -7316
rect 1229 -7350 1263 -7348
rect 1423 -7246 1457 -7244
rect 1423 -7278 1457 -7246
rect 1423 -7348 1457 -7316
rect 1423 -7350 1457 -7348
rect 1681 -7246 1715 -7244
rect 1681 -7278 1715 -7246
rect 1681 -7348 1715 -7316
rect 1681 -7350 1715 -7348
rect 1939 -7246 1973 -7244
rect 1939 -7278 1973 -7246
rect 1939 -7348 1973 -7316
rect 1939 -7350 1973 -7348
rect 2197 -7246 2231 -7244
rect 2197 -7278 2231 -7246
rect 2197 -7348 2231 -7316
rect 2197 -7350 2231 -7348
rect 2455 -7246 2489 -7244
rect 2455 -7278 2489 -7246
rect 2455 -7348 2489 -7316
rect 2455 -7350 2489 -7348
rect 2649 -7246 2683 -7244
rect 2649 -7278 2683 -7246
rect 2649 -7348 2683 -7316
rect 2649 -7350 2683 -7348
rect 2907 -7246 2941 -7244
rect 2907 -7278 2941 -7246
rect 2907 -7348 2941 -7316
rect 2907 -7350 2941 -7348
rect 3165 -7246 3199 -7244
rect 3165 -7278 3199 -7246
rect 3165 -7348 3199 -7316
rect 3165 -7350 3199 -7348
rect 3423 -7246 3457 -7244
rect 3423 -7278 3457 -7246
rect 3423 -7348 3457 -7316
rect 3423 -7350 3457 -7348
rect 3617 -7246 3651 -7244
rect 3617 -7278 3651 -7246
rect 3617 -7348 3651 -7316
rect 3617 -7350 3651 -7348
rect 3875 -7246 3909 -7244
rect 3875 -7278 3909 -7246
rect 3875 -7348 3909 -7316
rect 3875 -7350 3909 -7348
rect 4133 -7246 4167 -7244
rect 4133 -7278 4167 -7246
rect 4133 -7348 4167 -7316
rect 4133 -7350 4167 -7348
rect 4391 -7246 4425 -7244
rect 4391 -7278 4425 -7246
rect 4391 -7348 4425 -7316
rect 4391 -7350 4425 -7348
rect 4649 -7246 4683 -7244
rect 4649 -7278 4683 -7246
rect 4649 -7348 4683 -7316
rect 4649 -7350 4683 -7348
rect 4842 -7246 4876 -7244
rect 4842 -7278 4876 -7246
rect 4842 -7348 4876 -7316
rect 4842 -7350 4876 -7348
rect 5100 -7246 5134 -7244
rect 5100 -7278 5134 -7246
rect 5100 -7348 5134 -7316
rect 5100 -7350 5134 -7348
rect 5214 -7198 5248 -7178
rect 9573 -6910 9607 -6876
rect 9573 -6974 9607 -6948
rect 9573 -6982 9607 -6974
rect 9573 -7042 9607 -7020
rect 9573 -7054 9607 -7042
rect 9573 -7110 9607 -7092
rect 9573 -7126 9607 -7110
rect 9573 -7178 9607 -7164
rect 5214 -7246 5248 -7236
rect 5214 -7270 5248 -7246
rect 5214 -7314 5248 -7308
rect 5214 -7342 5248 -7314
rect 5214 -7382 5248 -7380
rect 5214 -7414 5248 -7382
rect 5328 -7246 5362 -7244
rect 5328 -7278 5362 -7246
rect 5328 -7348 5362 -7316
rect 5328 -7350 5362 -7348
rect 5586 -7246 5620 -7244
rect 5586 -7278 5620 -7246
rect 5586 -7348 5620 -7316
rect 5586 -7350 5620 -7348
rect 5780 -7246 5814 -7244
rect 5780 -7278 5814 -7246
rect 5780 -7348 5814 -7316
rect 5780 -7350 5814 -7348
rect 6038 -7246 6072 -7244
rect 6038 -7278 6072 -7246
rect 6038 -7348 6072 -7316
rect 6038 -7350 6072 -7348
rect 6296 -7246 6330 -7244
rect 6296 -7278 6330 -7246
rect 6296 -7348 6330 -7316
rect 6296 -7350 6330 -7348
rect 6554 -7246 6588 -7244
rect 6554 -7278 6588 -7246
rect 6554 -7348 6588 -7316
rect 6554 -7350 6588 -7348
rect 6812 -7246 6846 -7244
rect 6812 -7278 6846 -7246
rect 6812 -7348 6846 -7316
rect 6812 -7350 6846 -7348
rect 7006 -7246 7040 -7244
rect 7006 -7278 7040 -7246
rect 7006 -7348 7040 -7316
rect 7006 -7350 7040 -7348
rect 7264 -7246 7298 -7244
rect 7264 -7278 7298 -7246
rect 7264 -7348 7298 -7316
rect 7264 -7350 7298 -7348
rect 7522 -7246 7556 -7244
rect 7522 -7278 7556 -7246
rect 7522 -7348 7556 -7316
rect 7522 -7350 7556 -7348
rect 7780 -7246 7814 -7244
rect 7780 -7278 7814 -7246
rect 7780 -7348 7814 -7316
rect 7780 -7350 7814 -7348
rect 7974 -7246 8008 -7244
rect 7974 -7278 8008 -7246
rect 7974 -7348 8008 -7316
rect 7974 -7350 8008 -7348
rect 8232 -7246 8266 -7244
rect 8232 -7278 8266 -7246
rect 8232 -7348 8266 -7316
rect 8232 -7350 8266 -7348
rect 8490 -7246 8524 -7244
rect 8490 -7278 8524 -7246
rect 8490 -7348 8524 -7316
rect 8490 -7350 8524 -7348
rect 8748 -7246 8782 -7244
rect 8748 -7278 8782 -7246
rect 8748 -7348 8782 -7316
rect 8748 -7350 8782 -7348
rect 9006 -7246 9040 -7244
rect 9006 -7278 9040 -7246
rect 9006 -7348 9040 -7316
rect 9006 -7350 9040 -7348
rect 9200 -7246 9234 -7244
rect 9200 -7278 9234 -7246
rect 9200 -7348 9234 -7316
rect 9200 -7350 9234 -7348
rect 9458 -7246 9492 -7244
rect 9458 -7278 9492 -7246
rect 9458 -7348 9492 -7316
rect 9458 -7350 9492 -7348
rect 9573 -7198 9607 -7178
rect 13932 -6910 13966 -6876
rect 13932 -6974 13966 -6948
rect 13932 -6982 13966 -6974
rect 13932 -7042 13966 -7020
rect 13932 -7054 13966 -7042
rect 13932 -7110 13966 -7092
rect 13932 -7126 13966 -7110
rect 9573 -7246 9607 -7236
rect 9573 -7270 9607 -7246
rect 9573 -7314 9607 -7308
rect 9573 -7342 9607 -7314
rect 9573 -7382 9607 -7380
rect 856 -7484 890 -7452
rect 1064 -7478 1066 -7444
rect 1066 -7478 1098 -7444
rect 1136 -7478 1168 -7444
rect 1168 -7478 1170 -7444
rect 1516 -7478 1518 -7444
rect 1518 -7478 1550 -7444
rect 1588 -7478 1620 -7444
rect 1620 -7478 1622 -7444
rect 1774 -7478 1776 -7444
rect 1776 -7478 1808 -7444
rect 1846 -7478 1878 -7444
rect 1878 -7478 1880 -7444
rect 2032 -7478 2034 -7444
rect 2034 -7478 2066 -7444
rect 2104 -7478 2136 -7444
rect 2136 -7478 2138 -7444
rect 2290 -7478 2292 -7444
rect 2292 -7478 2324 -7444
rect 2362 -7478 2394 -7444
rect 2394 -7478 2396 -7444
rect 2742 -7478 2744 -7444
rect 2744 -7478 2776 -7444
rect 2814 -7478 2846 -7444
rect 2846 -7478 2848 -7444
rect 3000 -7478 3002 -7444
rect 3002 -7478 3034 -7444
rect 3072 -7478 3104 -7444
rect 3104 -7478 3106 -7444
rect 3258 -7478 3260 -7444
rect 3260 -7478 3292 -7444
rect 3330 -7478 3362 -7444
rect 3362 -7478 3364 -7444
rect 3710 -7478 3712 -7444
rect 3712 -7478 3744 -7444
rect 3782 -7478 3814 -7444
rect 3814 -7478 3816 -7444
rect 3968 -7478 3970 -7444
rect 3970 -7478 4002 -7444
rect 4040 -7478 4072 -7444
rect 4072 -7478 4074 -7444
rect 4226 -7478 4228 -7444
rect 4228 -7478 4260 -7444
rect 4298 -7478 4330 -7444
rect 4330 -7478 4332 -7444
rect 4484 -7478 4486 -7444
rect 4486 -7478 4518 -7444
rect 4556 -7478 4588 -7444
rect 4588 -7478 4590 -7444
rect 4935 -7478 4937 -7444
rect 4937 -7478 4969 -7444
rect 5007 -7478 5039 -7444
rect 5039 -7478 5041 -7444
rect 9573 -7414 9607 -7382
rect 9688 -7246 9722 -7244
rect 9688 -7278 9722 -7246
rect 9688 -7348 9722 -7316
rect 9688 -7350 9722 -7348
rect 9946 -7246 9980 -7244
rect 9946 -7278 9980 -7246
rect 9946 -7348 9980 -7316
rect 9946 -7350 9980 -7348
rect 10140 -7246 10174 -7244
rect 10140 -7278 10174 -7246
rect 10140 -7348 10174 -7316
rect 10140 -7350 10174 -7348
rect 10398 -7246 10432 -7244
rect 10398 -7278 10432 -7246
rect 10398 -7348 10432 -7316
rect 10398 -7350 10432 -7348
rect 10656 -7246 10690 -7244
rect 10656 -7278 10690 -7246
rect 10656 -7348 10690 -7316
rect 10656 -7350 10690 -7348
rect 10914 -7246 10948 -7244
rect 10914 -7278 10948 -7246
rect 10914 -7348 10948 -7316
rect 10914 -7350 10948 -7348
rect 11172 -7246 11206 -7244
rect 11172 -7278 11206 -7246
rect 11172 -7348 11206 -7316
rect 11172 -7350 11206 -7348
rect 11366 -7246 11400 -7244
rect 11366 -7278 11400 -7246
rect 11366 -7348 11400 -7316
rect 11366 -7350 11400 -7348
rect 11624 -7246 11658 -7244
rect 11624 -7278 11658 -7246
rect 11624 -7348 11658 -7316
rect 11624 -7350 11658 -7348
rect 11882 -7246 11916 -7244
rect 11882 -7278 11916 -7246
rect 11882 -7348 11916 -7316
rect 11882 -7350 11916 -7348
rect 12140 -7246 12174 -7244
rect 12140 -7278 12174 -7246
rect 12140 -7348 12174 -7316
rect 12140 -7350 12174 -7348
rect 12334 -7246 12368 -7244
rect 12334 -7278 12368 -7246
rect 12334 -7348 12368 -7316
rect 12334 -7350 12368 -7348
rect 12592 -7246 12626 -7244
rect 12592 -7278 12626 -7246
rect 12592 -7348 12626 -7316
rect 12592 -7350 12626 -7348
rect 12850 -7246 12884 -7244
rect 12850 -7278 12884 -7246
rect 12850 -7348 12884 -7316
rect 12850 -7350 12884 -7348
rect 13108 -7246 13142 -7244
rect 13108 -7278 13142 -7246
rect 13108 -7348 13142 -7316
rect 13108 -7350 13142 -7348
rect 13366 -7246 13400 -7244
rect 13366 -7278 13400 -7246
rect 13366 -7348 13400 -7316
rect 13366 -7350 13400 -7348
rect 13560 -7246 13594 -7244
rect 13560 -7278 13594 -7246
rect 13560 -7348 13594 -7316
rect 13560 -7350 13594 -7348
rect 13818 -7246 13852 -7244
rect 13818 -7278 13852 -7246
rect 13818 -7348 13852 -7316
rect 13818 -7350 13852 -7348
rect 13932 -7178 13966 -7164
rect 13932 -7198 13966 -7178
rect 18290 -6910 18324 -6876
rect 18290 -6974 18324 -6948
rect 18290 -6982 18324 -6974
rect 18290 -7042 18324 -7020
rect 18290 -7054 18324 -7042
rect 18290 -7110 18324 -7092
rect 18290 -7126 18324 -7110
rect 18290 -7178 18324 -7164
rect 13932 -7246 13966 -7236
rect 13932 -7270 13966 -7246
rect 13932 -7314 13966 -7308
rect 13932 -7342 13966 -7314
rect 856 -7486 890 -7484
rect 856 -7552 890 -7524
rect 856 -7558 890 -7552
rect 856 -7620 890 -7596
rect 856 -7630 890 -7620
rect 856 -7688 890 -7668
rect 856 -7702 890 -7688
rect 856 -7756 890 -7740
rect 856 -7774 890 -7756
rect 5214 -7484 5248 -7452
rect 5214 -7486 5248 -7484
rect 5421 -7478 5423 -7444
rect 5423 -7478 5455 -7444
rect 5493 -7478 5525 -7444
rect 5525 -7478 5527 -7444
rect 5873 -7478 5875 -7444
rect 5875 -7478 5907 -7444
rect 5945 -7478 5977 -7444
rect 5977 -7478 5979 -7444
rect 6131 -7478 6133 -7444
rect 6133 -7478 6165 -7444
rect 6203 -7478 6235 -7444
rect 6235 -7478 6237 -7444
rect 6389 -7478 6391 -7444
rect 6391 -7478 6423 -7444
rect 6461 -7478 6493 -7444
rect 6493 -7478 6495 -7444
rect 6647 -7478 6649 -7444
rect 6649 -7478 6681 -7444
rect 6719 -7478 6751 -7444
rect 6751 -7478 6753 -7444
rect 7099 -7478 7101 -7444
rect 7101 -7478 7133 -7444
rect 7171 -7478 7203 -7444
rect 7203 -7478 7205 -7444
rect 7357 -7478 7359 -7444
rect 7359 -7478 7391 -7444
rect 7429 -7478 7461 -7444
rect 7461 -7478 7463 -7444
rect 7615 -7478 7617 -7444
rect 7617 -7478 7649 -7444
rect 7687 -7478 7719 -7444
rect 7719 -7478 7721 -7444
rect 8067 -7478 8069 -7444
rect 8069 -7478 8101 -7444
rect 8139 -7478 8171 -7444
rect 8171 -7478 8173 -7444
rect 8325 -7478 8327 -7444
rect 8327 -7478 8359 -7444
rect 8397 -7478 8429 -7444
rect 8429 -7478 8431 -7444
rect 8583 -7478 8585 -7444
rect 8585 -7478 8617 -7444
rect 8655 -7478 8687 -7444
rect 8687 -7478 8689 -7444
rect 8841 -7478 8843 -7444
rect 8843 -7478 8875 -7444
rect 8913 -7478 8945 -7444
rect 8945 -7478 8947 -7444
rect 9293 -7478 9295 -7444
rect 9295 -7478 9327 -7444
rect 9365 -7478 9397 -7444
rect 9397 -7478 9399 -7444
rect 13932 -7382 13966 -7380
rect 13932 -7414 13966 -7382
rect 14046 -7246 14080 -7244
rect 14046 -7278 14080 -7246
rect 14046 -7348 14080 -7316
rect 14046 -7350 14080 -7348
rect 14304 -7246 14338 -7244
rect 14304 -7278 14338 -7246
rect 14304 -7348 14338 -7316
rect 14304 -7350 14338 -7348
rect 14497 -7246 14531 -7244
rect 14497 -7278 14531 -7246
rect 14497 -7348 14531 -7316
rect 14497 -7350 14531 -7348
rect 14755 -7246 14789 -7244
rect 14755 -7278 14789 -7246
rect 14755 -7348 14789 -7316
rect 14755 -7350 14789 -7348
rect 15013 -7246 15047 -7244
rect 15013 -7278 15047 -7246
rect 15013 -7348 15047 -7316
rect 15013 -7350 15047 -7348
rect 15271 -7246 15305 -7244
rect 15271 -7278 15305 -7246
rect 15271 -7348 15305 -7316
rect 15271 -7350 15305 -7348
rect 15529 -7246 15563 -7244
rect 15529 -7278 15563 -7246
rect 15529 -7348 15563 -7316
rect 15529 -7350 15563 -7348
rect 15723 -7246 15757 -7244
rect 15723 -7278 15757 -7246
rect 15723 -7348 15757 -7316
rect 15723 -7350 15757 -7348
rect 15981 -7246 16015 -7244
rect 15981 -7278 16015 -7246
rect 15981 -7348 16015 -7316
rect 15981 -7350 16015 -7348
rect 16239 -7246 16273 -7244
rect 16239 -7278 16273 -7246
rect 16239 -7348 16273 -7316
rect 16239 -7350 16273 -7348
rect 16497 -7246 16531 -7244
rect 16497 -7278 16531 -7246
rect 16497 -7348 16531 -7316
rect 16497 -7350 16531 -7348
rect 16691 -7246 16725 -7244
rect 16691 -7278 16725 -7246
rect 16691 -7348 16725 -7316
rect 16691 -7350 16725 -7348
rect 16949 -7246 16983 -7244
rect 16949 -7278 16983 -7246
rect 16949 -7348 16983 -7316
rect 16949 -7350 16983 -7348
rect 17207 -7246 17241 -7244
rect 17207 -7278 17241 -7246
rect 17207 -7348 17241 -7316
rect 17207 -7350 17241 -7348
rect 17465 -7246 17499 -7244
rect 17465 -7278 17499 -7246
rect 17465 -7348 17499 -7316
rect 17465 -7350 17499 -7348
rect 17723 -7246 17757 -7244
rect 17723 -7278 17757 -7246
rect 17723 -7348 17757 -7316
rect 17723 -7350 17757 -7348
rect 17917 -7246 17951 -7244
rect 17917 -7278 17951 -7246
rect 17917 -7348 17951 -7316
rect 17917 -7350 17951 -7348
rect 18175 -7246 18209 -7244
rect 18175 -7278 18209 -7246
rect 18175 -7348 18209 -7316
rect 18175 -7350 18209 -7348
rect 18290 -7198 18324 -7178
rect 18290 -7246 18324 -7236
rect 18290 -7270 18324 -7246
rect 18290 -7314 18324 -7308
rect 18290 -7342 18324 -7314
rect 18290 -7382 18324 -7380
rect 5214 -7552 5248 -7524
rect 5214 -7558 5248 -7552
rect 5214 -7620 5248 -7596
rect 5214 -7630 5248 -7620
rect 5214 -7688 5248 -7668
rect 5214 -7702 5248 -7688
rect 5214 -7756 5248 -7740
rect 5214 -7774 5248 -7756
rect 856 -7824 890 -7812
rect 856 -7846 890 -7824
rect 1064 -7840 1066 -7806
rect 1066 -7840 1098 -7806
rect 1136 -7840 1168 -7806
rect 1168 -7840 1170 -7806
rect 1516 -7840 1518 -7806
rect 1518 -7840 1550 -7806
rect 1588 -7840 1620 -7806
rect 1620 -7840 1622 -7806
rect 1774 -7840 1776 -7806
rect 1776 -7840 1808 -7806
rect 1846 -7840 1878 -7806
rect 1878 -7840 1880 -7806
rect 2032 -7840 2034 -7806
rect 2034 -7840 2066 -7806
rect 2104 -7840 2136 -7806
rect 2136 -7840 2138 -7806
rect 2290 -7840 2292 -7806
rect 2292 -7840 2324 -7806
rect 2362 -7840 2394 -7806
rect 2394 -7840 2396 -7806
rect 2742 -7840 2744 -7806
rect 2744 -7840 2776 -7806
rect 2814 -7840 2846 -7806
rect 2846 -7840 2848 -7806
rect 3000 -7840 3002 -7806
rect 3002 -7840 3034 -7806
rect 3072 -7840 3104 -7806
rect 3104 -7840 3106 -7806
rect 3258 -7840 3260 -7806
rect 3260 -7840 3292 -7806
rect 3330 -7840 3362 -7806
rect 3362 -7840 3364 -7806
rect 3710 -7840 3712 -7806
rect 3712 -7840 3744 -7806
rect 3782 -7840 3814 -7806
rect 3814 -7840 3816 -7806
rect 3968 -7840 3970 -7806
rect 3970 -7840 4002 -7806
rect 4040 -7840 4072 -7806
rect 4072 -7840 4074 -7806
rect 4226 -7840 4228 -7806
rect 4228 -7840 4260 -7806
rect 4298 -7840 4330 -7806
rect 4330 -7840 4332 -7806
rect 4484 -7840 4486 -7806
rect 4486 -7840 4518 -7806
rect 4556 -7840 4588 -7806
rect 4588 -7840 4590 -7806
rect 4935 -7840 4937 -7806
rect 4937 -7840 4969 -7806
rect 5007 -7840 5039 -7806
rect 5039 -7840 5041 -7806
rect 9573 -7484 9607 -7452
rect 9781 -7478 9783 -7444
rect 9783 -7478 9815 -7444
rect 9853 -7478 9885 -7444
rect 9885 -7478 9887 -7444
rect 10233 -7478 10235 -7444
rect 10235 -7478 10267 -7444
rect 10305 -7478 10337 -7444
rect 10337 -7478 10339 -7444
rect 10491 -7478 10493 -7444
rect 10493 -7478 10525 -7444
rect 10563 -7478 10595 -7444
rect 10595 -7478 10597 -7444
rect 10749 -7478 10751 -7444
rect 10751 -7478 10783 -7444
rect 10821 -7478 10853 -7444
rect 10853 -7478 10855 -7444
rect 11007 -7478 11009 -7444
rect 11009 -7478 11041 -7444
rect 11079 -7478 11111 -7444
rect 11111 -7478 11113 -7444
rect 11459 -7478 11461 -7444
rect 11461 -7478 11493 -7444
rect 11531 -7478 11563 -7444
rect 11563 -7478 11565 -7444
rect 11717 -7478 11719 -7444
rect 11719 -7478 11751 -7444
rect 11789 -7478 11821 -7444
rect 11821 -7478 11823 -7444
rect 11975 -7478 11977 -7444
rect 11977 -7478 12009 -7444
rect 12047 -7478 12079 -7444
rect 12079 -7478 12081 -7444
rect 12427 -7478 12429 -7444
rect 12429 -7478 12461 -7444
rect 12499 -7478 12531 -7444
rect 12531 -7478 12533 -7444
rect 12685 -7478 12687 -7444
rect 12687 -7478 12719 -7444
rect 12757 -7478 12789 -7444
rect 12789 -7478 12791 -7444
rect 12943 -7478 12945 -7444
rect 12945 -7478 12977 -7444
rect 13015 -7478 13047 -7444
rect 13047 -7478 13049 -7444
rect 13201 -7478 13203 -7444
rect 13203 -7478 13235 -7444
rect 13273 -7478 13305 -7444
rect 13305 -7478 13307 -7444
rect 13653 -7478 13655 -7444
rect 13655 -7478 13687 -7444
rect 13725 -7478 13757 -7444
rect 13757 -7478 13759 -7444
rect 18290 -7414 18324 -7382
rect 9573 -7486 9607 -7484
rect 9573 -7552 9607 -7524
rect 9573 -7558 9607 -7552
rect 9573 -7620 9607 -7596
rect 9573 -7630 9607 -7620
rect 9573 -7688 9607 -7668
rect 9573 -7702 9607 -7688
rect 9573 -7756 9607 -7740
rect 9573 -7774 9607 -7756
rect 5214 -7824 5248 -7812
rect 5214 -7846 5248 -7824
rect 5421 -7840 5423 -7806
rect 5423 -7840 5455 -7806
rect 5493 -7840 5525 -7806
rect 5525 -7840 5527 -7806
rect 5873 -7840 5875 -7806
rect 5875 -7840 5907 -7806
rect 5945 -7840 5977 -7806
rect 5977 -7840 5979 -7806
rect 6131 -7840 6133 -7806
rect 6133 -7840 6165 -7806
rect 6203 -7840 6235 -7806
rect 6235 -7840 6237 -7806
rect 6389 -7840 6391 -7806
rect 6391 -7840 6423 -7806
rect 6461 -7840 6493 -7806
rect 6493 -7840 6495 -7806
rect 6647 -7840 6649 -7806
rect 6649 -7840 6681 -7806
rect 6719 -7840 6751 -7806
rect 6751 -7840 6753 -7806
rect 7099 -7840 7101 -7806
rect 7101 -7840 7133 -7806
rect 7171 -7840 7203 -7806
rect 7203 -7840 7205 -7806
rect 7357 -7840 7359 -7806
rect 7359 -7840 7391 -7806
rect 7429 -7840 7461 -7806
rect 7461 -7840 7463 -7806
rect 7615 -7840 7617 -7806
rect 7617 -7840 7649 -7806
rect 7687 -7840 7719 -7806
rect 7719 -7840 7721 -7806
rect 8067 -7840 8069 -7806
rect 8069 -7840 8101 -7806
rect 8139 -7840 8171 -7806
rect 8171 -7840 8173 -7806
rect 8325 -7840 8327 -7806
rect 8327 -7840 8359 -7806
rect 8397 -7840 8429 -7806
rect 8429 -7840 8431 -7806
rect 8583 -7840 8585 -7806
rect 8585 -7840 8617 -7806
rect 8655 -7840 8687 -7806
rect 8687 -7840 8689 -7806
rect 8841 -7840 8843 -7806
rect 8843 -7840 8875 -7806
rect 8913 -7840 8945 -7806
rect 8945 -7840 8947 -7806
rect 9293 -7840 9295 -7806
rect 9295 -7840 9327 -7806
rect 9365 -7840 9397 -7806
rect 9397 -7840 9399 -7806
rect 13932 -7484 13966 -7452
rect 14139 -7478 14141 -7444
rect 14141 -7478 14173 -7444
rect 14211 -7478 14243 -7444
rect 14243 -7478 14245 -7444
rect 14590 -7478 14592 -7444
rect 14592 -7478 14624 -7444
rect 14662 -7478 14694 -7444
rect 14694 -7478 14696 -7444
rect 14848 -7478 14850 -7444
rect 14850 -7478 14882 -7444
rect 14920 -7478 14952 -7444
rect 14952 -7478 14954 -7444
rect 15106 -7478 15108 -7444
rect 15108 -7478 15140 -7444
rect 15178 -7478 15210 -7444
rect 15210 -7478 15212 -7444
rect 15364 -7478 15366 -7444
rect 15366 -7478 15398 -7444
rect 15436 -7478 15468 -7444
rect 15468 -7478 15470 -7444
rect 15816 -7478 15818 -7444
rect 15818 -7478 15850 -7444
rect 15888 -7478 15920 -7444
rect 15920 -7478 15922 -7444
rect 16074 -7478 16076 -7444
rect 16076 -7478 16108 -7444
rect 16146 -7478 16178 -7444
rect 16178 -7478 16180 -7444
rect 16332 -7478 16334 -7444
rect 16334 -7478 16366 -7444
rect 16404 -7478 16436 -7444
rect 16436 -7478 16438 -7444
rect 16784 -7478 16786 -7444
rect 16786 -7478 16818 -7444
rect 16856 -7478 16888 -7444
rect 16888 -7478 16890 -7444
rect 17042 -7478 17044 -7444
rect 17044 -7478 17076 -7444
rect 17114 -7478 17146 -7444
rect 17146 -7478 17148 -7444
rect 17300 -7478 17302 -7444
rect 17302 -7478 17334 -7444
rect 17372 -7478 17404 -7444
rect 17404 -7478 17406 -7444
rect 17558 -7478 17560 -7444
rect 17560 -7478 17592 -7444
rect 17630 -7478 17662 -7444
rect 17662 -7478 17664 -7444
rect 18010 -7478 18012 -7444
rect 18012 -7478 18044 -7444
rect 18082 -7478 18114 -7444
rect 18114 -7478 18116 -7444
rect 13932 -7486 13966 -7484
rect 13932 -7552 13966 -7524
rect 13932 -7558 13966 -7552
rect 13932 -7620 13966 -7596
rect 13932 -7630 13966 -7620
rect 13932 -7688 13966 -7668
rect 13932 -7702 13966 -7688
rect 13932 -7756 13966 -7740
rect 13932 -7774 13966 -7756
rect 9573 -7824 9607 -7812
rect 856 -7892 890 -7884
rect 856 -7918 890 -7892
rect 856 -7960 890 -7956
rect 856 -7990 890 -7960
rect 856 -8062 890 -8028
rect 971 -7936 1005 -7934
rect 971 -7968 1005 -7936
rect 971 -8038 1005 -8006
rect 971 -8040 1005 -8038
rect 1229 -7936 1263 -7934
rect 1229 -7968 1263 -7936
rect 1229 -8038 1263 -8006
rect 1229 -8040 1263 -8038
rect 1423 -7936 1457 -7934
rect 1423 -7968 1457 -7936
rect 1423 -8038 1457 -8006
rect 1423 -8040 1457 -8038
rect 1681 -7936 1715 -7934
rect 1681 -7968 1715 -7936
rect 1681 -8038 1715 -8006
rect 1681 -8040 1715 -8038
rect 1939 -7936 1973 -7934
rect 1939 -7968 1973 -7936
rect 1939 -8038 1973 -8006
rect 1939 -8040 1973 -8038
rect 2197 -7936 2231 -7934
rect 2197 -7968 2231 -7936
rect 2197 -8038 2231 -8006
rect 2197 -8040 2231 -8038
rect 2455 -7936 2489 -7934
rect 2455 -7968 2489 -7936
rect 2455 -8038 2489 -8006
rect 2455 -8040 2489 -8038
rect 2649 -7936 2683 -7934
rect 2649 -7968 2683 -7936
rect 2649 -8038 2683 -8006
rect 2649 -8040 2683 -8038
rect 2907 -7936 2941 -7934
rect 2907 -7968 2941 -7936
rect 2907 -8038 2941 -8006
rect 2907 -8040 2941 -8038
rect 3165 -7936 3199 -7934
rect 3165 -7968 3199 -7936
rect 3165 -8038 3199 -8006
rect 3165 -8040 3199 -8038
rect 3423 -7936 3457 -7934
rect 3423 -7968 3457 -7936
rect 3423 -8038 3457 -8006
rect 3423 -8040 3457 -8038
rect 3617 -7936 3651 -7934
rect 3617 -7968 3651 -7936
rect 3617 -8038 3651 -8006
rect 3617 -8040 3651 -8038
rect 3875 -7936 3909 -7934
rect 3875 -7968 3909 -7936
rect 3875 -8038 3909 -8006
rect 3875 -8040 3909 -8038
rect 4133 -7936 4167 -7934
rect 4133 -7968 4167 -7936
rect 4133 -8038 4167 -8006
rect 4133 -8040 4167 -8038
rect 4391 -7936 4425 -7934
rect 4391 -7968 4425 -7936
rect 4391 -8038 4425 -8006
rect 4391 -8040 4425 -8038
rect 4649 -7936 4683 -7934
rect 4649 -7968 4683 -7936
rect 4649 -8038 4683 -8006
rect 4649 -8040 4683 -8038
rect 4842 -7936 4876 -7934
rect 4842 -7968 4876 -7936
rect 4842 -8038 4876 -8006
rect 4842 -8040 4876 -8038
rect 5100 -7936 5134 -7934
rect 5100 -7968 5134 -7936
rect 5100 -8038 5134 -8006
rect 5100 -8040 5134 -8038
rect 9573 -7846 9607 -7824
rect 9781 -7840 9783 -7806
rect 9783 -7840 9815 -7806
rect 9853 -7840 9885 -7806
rect 9885 -7840 9887 -7806
rect 10233 -7840 10235 -7806
rect 10235 -7840 10267 -7806
rect 10305 -7840 10337 -7806
rect 10337 -7840 10339 -7806
rect 10491 -7840 10493 -7806
rect 10493 -7840 10525 -7806
rect 10563 -7840 10595 -7806
rect 10595 -7840 10597 -7806
rect 10749 -7840 10751 -7806
rect 10751 -7840 10783 -7806
rect 10821 -7840 10853 -7806
rect 10853 -7840 10855 -7806
rect 11007 -7840 11009 -7806
rect 11009 -7840 11041 -7806
rect 11079 -7840 11111 -7806
rect 11111 -7840 11113 -7806
rect 11459 -7840 11461 -7806
rect 11461 -7840 11493 -7806
rect 11531 -7840 11563 -7806
rect 11563 -7840 11565 -7806
rect 11717 -7840 11719 -7806
rect 11719 -7840 11751 -7806
rect 11789 -7840 11821 -7806
rect 11821 -7840 11823 -7806
rect 11975 -7840 11977 -7806
rect 11977 -7840 12009 -7806
rect 12047 -7840 12079 -7806
rect 12079 -7840 12081 -7806
rect 12427 -7840 12429 -7806
rect 12429 -7840 12461 -7806
rect 12499 -7840 12531 -7806
rect 12531 -7840 12533 -7806
rect 12685 -7840 12687 -7806
rect 12687 -7840 12719 -7806
rect 12757 -7840 12789 -7806
rect 12789 -7840 12791 -7806
rect 12943 -7840 12945 -7806
rect 12945 -7840 12977 -7806
rect 13015 -7840 13047 -7806
rect 13047 -7840 13049 -7806
rect 13201 -7840 13203 -7806
rect 13203 -7840 13235 -7806
rect 13273 -7840 13305 -7806
rect 13305 -7840 13307 -7806
rect 13653 -7840 13655 -7806
rect 13655 -7840 13687 -7806
rect 13725 -7840 13757 -7806
rect 13757 -7840 13759 -7806
rect 18290 -7484 18324 -7452
rect 18290 -7486 18324 -7484
rect 18290 -7552 18324 -7524
rect 18290 -7558 18324 -7552
rect 18290 -7620 18324 -7596
rect 18290 -7630 18324 -7620
rect 18290 -7688 18324 -7668
rect 18290 -7702 18324 -7688
rect 18290 -7756 18324 -7740
rect 18290 -7774 18324 -7756
rect 5214 -7892 5248 -7884
rect 5214 -7918 5248 -7892
rect 5214 -7960 5248 -7956
rect 5214 -7990 5248 -7960
rect 5214 -8062 5248 -8028
rect 856 -8130 890 -8100
rect 856 -8134 890 -8130
rect 856 -8198 890 -8172
rect 856 -8206 890 -8198
rect 856 -8266 890 -8244
rect 856 -8278 890 -8266
rect 856 -8334 890 -8316
rect 856 -8350 890 -8334
rect 856 -8402 890 -8388
rect 5328 -7936 5362 -7934
rect 5328 -7968 5362 -7936
rect 5328 -8038 5362 -8006
rect 5328 -8040 5362 -8038
rect 5586 -7936 5620 -7934
rect 5586 -7968 5620 -7936
rect 5586 -8038 5620 -8006
rect 5586 -8040 5620 -8038
rect 5780 -7936 5814 -7934
rect 5780 -7968 5814 -7936
rect 5780 -8038 5814 -8006
rect 5780 -8040 5814 -8038
rect 6038 -7936 6072 -7934
rect 6038 -7968 6072 -7936
rect 6038 -8038 6072 -8006
rect 6038 -8040 6072 -8038
rect 6296 -7936 6330 -7934
rect 6296 -7968 6330 -7936
rect 6296 -8038 6330 -8006
rect 6296 -8040 6330 -8038
rect 6554 -7936 6588 -7934
rect 6554 -7968 6588 -7936
rect 6554 -8038 6588 -8006
rect 6554 -8040 6588 -8038
rect 6812 -7936 6846 -7934
rect 6812 -7968 6846 -7936
rect 6812 -8038 6846 -8006
rect 6812 -8040 6846 -8038
rect 7006 -7936 7040 -7934
rect 7006 -7968 7040 -7936
rect 7006 -8038 7040 -8006
rect 7006 -8040 7040 -8038
rect 7264 -7936 7298 -7934
rect 7264 -7968 7298 -7936
rect 7264 -8038 7298 -8006
rect 7264 -8040 7298 -8038
rect 7522 -7936 7556 -7934
rect 7522 -7968 7556 -7936
rect 7522 -8038 7556 -8006
rect 7522 -8040 7556 -8038
rect 7780 -7936 7814 -7934
rect 7780 -7968 7814 -7936
rect 7780 -8038 7814 -8006
rect 7780 -8040 7814 -8038
rect 7974 -7936 8008 -7934
rect 7974 -7968 8008 -7936
rect 7974 -8038 8008 -8006
rect 7974 -8040 8008 -8038
rect 8232 -7936 8266 -7934
rect 8232 -7968 8266 -7936
rect 8232 -8038 8266 -8006
rect 8232 -8040 8266 -8038
rect 8490 -7936 8524 -7934
rect 8490 -7968 8524 -7936
rect 8490 -8038 8524 -8006
rect 8490 -8040 8524 -8038
rect 8748 -7936 8782 -7934
rect 8748 -7968 8782 -7936
rect 8748 -8038 8782 -8006
rect 8748 -8040 8782 -8038
rect 9006 -7936 9040 -7934
rect 9006 -7968 9040 -7936
rect 9006 -8038 9040 -8006
rect 9006 -8040 9040 -8038
rect 9200 -7936 9234 -7934
rect 9200 -7968 9234 -7936
rect 9200 -8038 9234 -8006
rect 9200 -8040 9234 -8038
rect 9458 -7936 9492 -7934
rect 9458 -7968 9492 -7936
rect 9458 -8038 9492 -8006
rect 9458 -8040 9492 -8038
rect 13932 -7824 13966 -7812
rect 13932 -7846 13966 -7824
rect 14139 -7840 14141 -7806
rect 14141 -7840 14173 -7806
rect 14211 -7840 14243 -7806
rect 14243 -7840 14245 -7806
rect 14590 -7840 14592 -7806
rect 14592 -7840 14624 -7806
rect 14662 -7840 14694 -7806
rect 14694 -7840 14696 -7806
rect 14848 -7840 14850 -7806
rect 14850 -7840 14882 -7806
rect 14920 -7840 14952 -7806
rect 14952 -7840 14954 -7806
rect 15106 -7840 15108 -7806
rect 15108 -7840 15140 -7806
rect 15178 -7840 15210 -7806
rect 15210 -7840 15212 -7806
rect 15364 -7840 15366 -7806
rect 15366 -7840 15398 -7806
rect 15436 -7840 15468 -7806
rect 15468 -7840 15470 -7806
rect 15816 -7840 15818 -7806
rect 15818 -7840 15850 -7806
rect 15888 -7840 15920 -7806
rect 15920 -7840 15922 -7806
rect 16074 -7840 16076 -7806
rect 16076 -7840 16108 -7806
rect 16146 -7840 16178 -7806
rect 16178 -7840 16180 -7806
rect 16332 -7840 16334 -7806
rect 16334 -7840 16366 -7806
rect 16404 -7840 16436 -7806
rect 16436 -7840 16438 -7806
rect 16784 -7840 16786 -7806
rect 16786 -7840 16818 -7806
rect 16856 -7840 16888 -7806
rect 16888 -7840 16890 -7806
rect 17042 -7840 17044 -7806
rect 17044 -7840 17076 -7806
rect 17114 -7840 17146 -7806
rect 17146 -7840 17148 -7806
rect 17300 -7840 17302 -7806
rect 17302 -7840 17334 -7806
rect 17372 -7840 17404 -7806
rect 17404 -7840 17406 -7806
rect 17558 -7840 17560 -7806
rect 17560 -7840 17592 -7806
rect 17630 -7840 17662 -7806
rect 17662 -7840 17664 -7806
rect 18010 -7840 18012 -7806
rect 18012 -7840 18044 -7806
rect 18082 -7840 18114 -7806
rect 18114 -7840 18116 -7806
rect 18290 -7824 18324 -7812
rect 9573 -7892 9607 -7884
rect 9573 -7918 9607 -7892
rect 9573 -7960 9607 -7956
rect 9573 -7990 9607 -7960
rect 9573 -8062 9607 -8028
rect 5214 -8130 5248 -8100
rect 5214 -8134 5248 -8130
rect 5214 -8198 5248 -8172
rect 5214 -8206 5248 -8198
rect 5214 -8266 5248 -8244
rect 5214 -8278 5248 -8266
rect 5214 -8334 5248 -8316
rect 5214 -8350 5248 -8334
rect 5214 -8402 5248 -8388
rect 9688 -7936 9722 -7934
rect 9688 -7968 9722 -7936
rect 9688 -8038 9722 -8006
rect 9688 -8040 9722 -8038
rect 9946 -7936 9980 -7934
rect 9946 -7968 9980 -7936
rect 9946 -8038 9980 -8006
rect 9946 -8040 9980 -8038
rect 10140 -7936 10174 -7934
rect 10140 -7968 10174 -7936
rect 10140 -8038 10174 -8006
rect 10140 -8040 10174 -8038
rect 10398 -7936 10432 -7934
rect 10398 -7968 10432 -7936
rect 10398 -8038 10432 -8006
rect 10398 -8040 10432 -8038
rect 10656 -7936 10690 -7934
rect 10656 -7968 10690 -7936
rect 10656 -8038 10690 -8006
rect 10656 -8040 10690 -8038
rect 10914 -7936 10948 -7934
rect 10914 -7968 10948 -7936
rect 10914 -8038 10948 -8006
rect 10914 -8040 10948 -8038
rect 11172 -7936 11206 -7934
rect 11172 -7968 11206 -7936
rect 11172 -8038 11206 -8006
rect 11172 -8040 11206 -8038
rect 11366 -7936 11400 -7934
rect 11366 -7968 11400 -7936
rect 11366 -8038 11400 -8006
rect 11366 -8040 11400 -8038
rect 11624 -7936 11658 -7934
rect 11624 -7968 11658 -7936
rect 11624 -8038 11658 -8006
rect 11624 -8040 11658 -8038
rect 11882 -7936 11916 -7934
rect 11882 -7968 11916 -7936
rect 11882 -8038 11916 -8006
rect 11882 -8040 11916 -8038
rect 12140 -7936 12174 -7934
rect 12140 -7968 12174 -7936
rect 12140 -8038 12174 -8006
rect 12140 -8040 12174 -8038
rect 12334 -7936 12368 -7934
rect 12334 -7968 12368 -7936
rect 12334 -8038 12368 -8006
rect 12334 -8040 12368 -8038
rect 12592 -7936 12626 -7934
rect 12592 -7968 12626 -7936
rect 12592 -8038 12626 -8006
rect 12592 -8040 12626 -8038
rect 12850 -7936 12884 -7934
rect 12850 -7968 12884 -7936
rect 12850 -8038 12884 -8006
rect 12850 -8040 12884 -8038
rect 13108 -7936 13142 -7934
rect 13108 -7968 13142 -7936
rect 13108 -8038 13142 -8006
rect 13108 -8040 13142 -8038
rect 13366 -7936 13400 -7934
rect 13366 -7968 13400 -7936
rect 13366 -8038 13400 -8006
rect 13366 -8040 13400 -8038
rect 13560 -7936 13594 -7934
rect 13560 -7968 13594 -7936
rect 13560 -8038 13594 -8006
rect 13560 -8040 13594 -8038
rect 13818 -7936 13852 -7934
rect 13818 -7968 13852 -7936
rect 13818 -8038 13852 -8006
rect 13818 -8040 13852 -8038
rect 18290 -7846 18324 -7824
rect 13932 -7892 13966 -7884
rect 13932 -7918 13966 -7892
rect 13932 -7960 13966 -7956
rect 13932 -7990 13966 -7960
rect 13932 -8062 13966 -8028
rect 9573 -8130 9607 -8100
rect 9573 -8134 9607 -8130
rect 9573 -8198 9607 -8172
rect 9573 -8206 9607 -8198
rect 9573 -8266 9607 -8244
rect 9573 -8278 9607 -8266
rect 9573 -8334 9607 -8316
rect 9573 -8350 9607 -8334
rect 9573 -8402 9607 -8388
rect 14046 -7936 14080 -7934
rect 14046 -7968 14080 -7936
rect 14046 -8038 14080 -8006
rect 14046 -8040 14080 -8038
rect 14304 -7936 14338 -7934
rect 14304 -7968 14338 -7936
rect 14304 -8038 14338 -8006
rect 14304 -8040 14338 -8038
rect 14497 -7936 14531 -7934
rect 14497 -7968 14531 -7936
rect 14497 -8038 14531 -8006
rect 14497 -8040 14531 -8038
rect 14755 -7936 14789 -7934
rect 14755 -7968 14789 -7936
rect 14755 -8038 14789 -8006
rect 14755 -8040 14789 -8038
rect 15013 -7936 15047 -7934
rect 15013 -7968 15047 -7936
rect 15013 -8038 15047 -8006
rect 15013 -8040 15047 -8038
rect 15271 -7936 15305 -7934
rect 15271 -7968 15305 -7936
rect 15271 -8038 15305 -8006
rect 15271 -8040 15305 -8038
rect 15529 -7936 15563 -7934
rect 15529 -7968 15563 -7936
rect 15529 -8038 15563 -8006
rect 15529 -8040 15563 -8038
rect 15723 -7936 15757 -7934
rect 15723 -7968 15757 -7936
rect 15723 -8038 15757 -8006
rect 15723 -8040 15757 -8038
rect 15981 -7936 16015 -7934
rect 15981 -7968 16015 -7936
rect 15981 -8038 16015 -8006
rect 15981 -8040 16015 -8038
rect 16239 -7936 16273 -7934
rect 16239 -7968 16273 -7936
rect 16239 -8038 16273 -8006
rect 16239 -8040 16273 -8038
rect 16497 -7936 16531 -7934
rect 16497 -7968 16531 -7936
rect 16497 -8038 16531 -8006
rect 16497 -8040 16531 -8038
rect 16691 -7936 16725 -7934
rect 16691 -7968 16725 -7936
rect 16691 -8038 16725 -8006
rect 16691 -8040 16725 -8038
rect 16949 -7936 16983 -7934
rect 16949 -7968 16983 -7936
rect 16949 -8038 16983 -8006
rect 16949 -8040 16983 -8038
rect 17207 -7936 17241 -7934
rect 17207 -7968 17241 -7936
rect 17207 -8038 17241 -8006
rect 17207 -8040 17241 -8038
rect 17465 -7936 17499 -7934
rect 17465 -7968 17499 -7936
rect 17465 -8038 17499 -8006
rect 17465 -8040 17499 -8038
rect 17723 -7936 17757 -7934
rect 17723 -7968 17757 -7936
rect 17723 -8038 17757 -8006
rect 17723 -8040 17757 -8038
rect 17917 -7936 17951 -7934
rect 17917 -7968 17951 -7936
rect 17917 -8038 17951 -8006
rect 17917 -8040 17951 -8038
rect 18175 -7936 18209 -7934
rect 18175 -7968 18209 -7936
rect 18175 -8038 18209 -8006
rect 18175 -8040 18209 -8038
rect 18290 -7892 18324 -7884
rect 18290 -7918 18324 -7892
rect 18290 -7960 18324 -7956
rect 18290 -7990 18324 -7960
rect 18290 -8062 18324 -8028
rect 13932 -8130 13966 -8100
rect 13932 -8134 13966 -8130
rect 13932 -8198 13966 -8172
rect 13932 -8206 13966 -8198
rect 13932 -8266 13966 -8244
rect 13932 -8278 13966 -8266
rect 13932 -8334 13966 -8316
rect 13932 -8350 13966 -8334
rect 13932 -8402 13966 -8388
rect 18290 -8130 18324 -8100
rect 18290 -8134 18324 -8130
rect 18290 -8198 18324 -8172
rect 18290 -8206 18324 -8198
rect 18290 -8266 18324 -8244
rect 18290 -8278 18324 -8266
rect 18290 -8334 18324 -8316
rect 18290 -8350 18324 -8334
rect 18290 -8402 18324 -8388
rect 856 -8422 890 -8402
rect 5214 -8422 5248 -8402
rect 9573 -8422 9607 -8402
rect 13932 -8422 13966 -8402
rect 18290 -8422 18324 -8402
rect 856 -8470 890 -8460
rect 856 -8494 890 -8470
rect 856 -8538 890 -8532
rect 856 -8566 890 -8538
rect 856 -8606 890 -8604
rect 856 -8638 890 -8606
rect 856 -8708 890 -8676
rect 856 -8710 890 -8708
rect 856 -8776 890 -8748
rect 856 -8782 890 -8776
rect 856 -8844 890 -8820
rect 5214 -8470 5248 -8460
rect 5214 -8494 5248 -8470
rect 5214 -8538 5248 -8532
rect 5214 -8566 5248 -8538
rect 5214 -8606 5248 -8604
rect 5214 -8638 5248 -8606
rect 5214 -8708 5248 -8676
rect 5214 -8710 5248 -8708
rect 5214 -8776 5248 -8748
rect 5214 -8782 5248 -8776
rect 856 -8854 890 -8844
rect 856 -8912 890 -8892
rect 856 -8926 890 -8912
rect 856 -8980 890 -8964
rect 856 -8998 890 -8980
rect 971 -8880 1005 -8878
rect 971 -8912 1005 -8880
rect 971 -8982 1005 -8950
rect 971 -8984 1005 -8982
rect 1229 -8880 1263 -8878
rect 1229 -8912 1263 -8880
rect 1229 -8982 1263 -8950
rect 1229 -8984 1263 -8982
rect 1423 -8880 1457 -8878
rect 1423 -8912 1457 -8880
rect 1423 -8982 1457 -8950
rect 1423 -8984 1457 -8982
rect 1681 -8880 1715 -8878
rect 1681 -8912 1715 -8880
rect 1681 -8982 1715 -8950
rect 1681 -8984 1715 -8982
rect 1939 -8880 1973 -8878
rect 1939 -8912 1973 -8880
rect 1939 -8982 1973 -8950
rect 1939 -8984 1973 -8982
rect 2197 -8880 2231 -8878
rect 2197 -8912 2231 -8880
rect 2197 -8982 2231 -8950
rect 2197 -8984 2231 -8982
rect 2455 -8880 2489 -8878
rect 2455 -8912 2489 -8880
rect 2455 -8982 2489 -8950
rect 2455 -8984 2489 -8982
rect 2649 -8880 2683 -8878
rect 2649 -8912 2683 -8880
rect 2649 -8982 2683 -8950
rect 2649 -8984 2683 -8982
rect 2907 -8880 2941 -8878
rect 2907 -8912 2941 -8880
rect 2907 -8982 2941 -8950
rect 2907 -8984 2941 -8982
rect 3165 -8880 3199 -8878
rect 3165 -8912 3199 -8880
rect 3165 -8982 3199 -8950
rect 3165 -8984 3199 -8982
rect 3423 -8880 3457 -8878
rect 3423 -8912 3457 -8880
rect 3423 -8982 3457 -8950
rect 3423 -8984 3457 -8982
rect 3617 -8880 3651 -8878
rect 3617 -8912 3651 -8880
rect 3617 -8982 3651 -8950
rect 3617 -8984 3651 -8982
rect 3875 -8880 3909 -8878
rect 3875 -8912 3909 -8880
rect 3875 -8982 3909 -8950
rect 3875 -8984 3909 -8982
rect 4133 -8880 4167 -8878
rect 4133 -8912 4167 -8880
rect 4133 -8982 4167 -8950
rect 4133 -8984 4167 -8982
rect 4391 -8880 4425 -8878
rect 4391 -8912 4425 -8880
rect 4391 -8982 4425 -8950
rect 4391 -8984 4425 -8982
rect 4649 -8880 4683 -8878
rect 4649 -8912 4683 -8880
rect 4649 -8982 4683 -8950
rect 4649 -8984 4683 -8982
rect 4842 -8880 4876 -8878
rect 4842 -8912 4876 -8880
rect 4842 -8982 4876 -8950
rect 4842 -8984 4876 -8982
rect 5100 -8880 5134 -8878
rect 5100 -8912 5134 -8880
rect 5100 -8982 5134 -8950
rect 5100 -8984 5134 -8982
rect 5214 -8844 5248 -8820
rect 5214 -8854 5248 -8844
rect 9573 -8470 9607 -8460
rect 9573 -8494 9607 -8470
rect 9573 -8538 9607 -8532
rect 9573 -8566 9607 -8538
rect 9573 -8606 9607 -8604
rect 9573 -8638 9607 -8606
rect 9573 -8708 9607 -8676
rect 9573 -8710 9607 -8708
rect 9573 -8776 9607 -8748
rect 9573 -8782 9607 -8776
rect 5214 -8912 5248 -8892
rect 5214 -8926 5248 -8912
rect 5214 -8980 5248 -8964
rect 5214 -8998 5248 -8980
rect 856 -9070 890 -9036
rect 5328 -8880 5362 -8878
rect 5328 -8912 5362 -8880
rect 5328 -8982 5362 -8950
rect 5328 -8984 5362 -8982
rect 5586 -8880 5620 -8878
rect 5586 -8912 5620 -8880
rect 5586 -8982 5620 -8950
rect 5586 -8984 5620 -8982
rect 5780 -8880 5814 -8878
rect 5780 -8912 5814 -8880
rect 5780 -8982 5814 -8950
rect 5780 -8984 5814 -8982
rect 6038 -8880 6072 -8878
rect 6038 -8912 6072 -8880
rect 6038 -8982 6072 -8950
rect 6038 -8984 6072 -8982
rect 6296 -8880 6330 -8878
rect 6296 -8912 6330 -8880
rect 6296 -8982 6330 -8950
rect 6296 -8984 6330 -8982
rect 6554 -8880 6588 -8878
rect 6554 -8912 6588 -8880
rect 6554 -8982 6588 -8950
rect 6554 -8984 6588 -8982
rect 6812 -8880 6846 -8878
rect 6812 -8912 6846 -8880
rect 6812 -8982 6846 -8950
rect 6812 -8984 6846 -8982
rect 7006 -8880 7040 -8878
rect 7006 -8912 7040 -8880
rect 7006 -8982 7040 -8950
rect 7006 -8984 7040 -8982
rect 7264 -8880 7298 -8878
rect 7264 -8912 7298 -8880
rect 7264 -8982 7298 -8950
rect 7264 -8984 7298 -8982
rect 7522 -8880 7556 -8878
rect 7522 -8912 7556 -8880
rect 7522 -8982 7556 -8950
rect 7522 -8984 7556 -8982
rect 7780 -8880 7814 -8878
rect 7780 -8912 7814 -8880
rect 7780 -8982 7814 -8950
rect 7780 -8984 7814 -8982
rect 7974 -8880 8008 -8878
rect 7974 -8912 8008 -8880
rect 7974 -8982 8008 -8950
rect 7974 -8984 8008 -8982
rect 8232 -8880 8266 -8878
rect 8232 -8912 8266 -8880
rect 8232 -8982 8266 -8950
rect 8232 -8984 8266 -8982
rect 8490 -8880 8524 -8878
rect 8490 -8912 8524 -8880
rect 8490 -8982 8524 -8950
rect 8490 -8984 8524 -8982
rect 8748 -8880 8782 -8878
rect 8748 -8912 8782 -8880
rect 8748 -8982 8782 -8950
rect 8748 -8984 8782 -8982
rect 9006 -8880 9040 -8878
rect 9006 -8912 9040 -8880
rect 9006 -8982 9040 -8950
rect 9006 -8984 9040 -8982
rect 9200 -8880 9234 -8878
rect 9200 -8912 9234 -8880
rect 9200 -8982 9234 -8950
rect 9200 -8984 9234 -8982
rect 9458 -8880 9492 -8878
rect 9458 -8912 9492 -8880
rect 9458 -8982 9492 -8950
rect 9458 -8984 9492 -8982
rect 9573 -8844 9607 -8820
rect 13932 -8470 13966 -8460
rect 13932 -8494 13966 -8470
rect 13932 -8538 13966 -8532
rect 13932 -8566 13966 -8538
rect 13932 -8606 13966 -8604
rect 13932 -8638 13966 -8606
rect 13932 -8708 13966 -8676
rect 13932 -8710 13966 -8708
rect 13932 -8776 13966 -8748
rect 13932 -8782 13966 -8776
rect 9573 -8854 9607 -8844
rect 9573 -8912 9607 -8892
rect 9573 -8926 9607 -8912
rect 9573 -8980 9607 -8964
rect 9573 -8998 9607 -8980
rect 5214 -9070 5248 -9036
rect 1064 -9112 1066 -9078
rect 1066 -9112 1098 -9078
rect 1136 -9112 1168 -9078
rect 1168 -9112 1170 -9078
rect 1516 -9112 1518 -9078
rect 1518 -9112 1550 -9078
rect 1588 -9112 1620 -9078
rect 1620 -9112 1622 -9078
rect 1774 -9112 1776 -9078
rect 1776 -9112 1808 -9078
rect 1846 -9112 1878 -9078
rect 1878 -9112 1880 -9078
rect 2032 -9112 2034 -9078
rect 2034 -9112 2066 -9078
rect 2104 -9112 2136 -9078
rect 2136 -9112 2138 -9078
rect 2290 -9112 2292 -9078
rect 2292 -9112 2324 -9078
rect 2362 -9112 2394 -9078
rect 2394 -9112 2396 -9078
rect 2742 -9112 2744 -9078
rect 2744 -9112 2776 -9078
rect 2814 -9112 2846 -9078
rect 2846 -9112 2848 -9078
rect 3000 -9112 3002 -9078
rect 3002 -9112 3034 -9078
rect 3072 -9112 3104 -9078
rect 3104 -9112 3106 -9078
rect 3258 -9112 3260 -9078
rect 3260 -9112 3292 -9078
rect 3330 -9112 3362 -9078
rect 3362 -9112 3364 -9078
rect 3710 -9112 3712 -9078
rect 3712 -9112 3744 -9078
rect 3782 -9112 3814 -9078
rect 3814 -9112 3816 -9078
rect 3968 -9112 3970 -9078
rect 3970 -9112 4002 -9078
rect 4040 -9112 4072 -9078
rect 4072 -9112 4074 -9078
rect 4226 -9112 4228 -9078
rect 4228 -9112 4260 -9078
rect 4298 -9112 4330 -9078
rect 4330 -9112 4332 -9078
rect 4484 -9112 4486 -9078
rect 4486 -9112 4518 -9078
rect 4556 -9112 4588 -9078
rect 4588 -9112 4590 -9078
rect 4935 -9112 4937 -9078
rect 4937 -9112 4969 -9078
rect 5007 -9112 5039 -9078
rect 5039 -9112 5041 -9078
rect 9688 -8880 9722 -8878
rect 9688 -8912 9722 -8880
rect 9688 -8982 9722 -8950
rect 9688 -8984 9722 -8982
rect 9946 -8880 9980 -8878
rect 9946 -8912 9980 -8880
rect 9946 -8982 9980 -8950
rect 9946 -8984 9980 -8982
rect 10140 -8880 10174 -8878
rect 10140 -8912 10174 -8880
rect 10140 -8982 10174 -8950
rect 10140 -8984 10174 -8982
rect 10398 -8880 10432 -8878
rect 10398 -8912 10432 -8880
rect 10398 -8982 10432 -8950
rect 10398 -8984 10432 -8982
rect 10656 -8880 10690 -8878
rect 10656 -8912 10690 -8880
rect 10656 -8982 10690 -8950
rect 10656 -8984 10690 -8982
rect 10914 -8880 10948 -8878
rect 10914 -8912 10948 -8880
rect 10914 -8982 10948 -8950
rect 10914 -8984 10948 -8982
rect 11172 -8880 11206 -8878
rect 11172 -8912 11206 -8880
rect 11172 -8982 11206 -8950
rect 11172 -8984 11206 -8982
rect 11366 -8880 11400 -8878
rect 11366 -8912 11400 -8880
rect 11366 -8982 11400 -8950
rect 11366 -8984 11400 -8982
rect 11624 -8880 11658 -8878
rect 11624 -8912 11658 -8880
rect 11624 -8982 11658 -8950
rect 11624 -8984 11658 -8982
rect 11882 -8880 11916 -8878
rect 11882 -8912 11916 -8880
rect 11882 -8982 11916 -8950
rect 11882 -8984 11916 -8982
rect 12140 -8880 12174 -8878
rect 12140 -8912 12174 -8880
rect 12140 -8982 12174 -8950
rect 12140 -8984 12174 -8982
rect 12334 -8880 12368 -8878
rect 12334 -8912 12368 -8880
rect 12334 -8982 12368 -8950
rect 12334 -8984 12368 -8982
rect 12592 -8880 12626 -8878
rect 12592 -8912 12626 -8880
rect 12592 -8982 12626 -8950
rect 12592 -8984 12626 -8982
rect 12850 -8880 12884 -8878
rect 12850 -8912 12884 -8880
rect 12850 -8982 12884 -8950
rect 12850 -8984 12884 -8982
rect 13108 -8880 13142 -8878
rect 13108 -8912 13142 -8880
rect 13108 -8982 13142 -8950
rect 13108 -8984 13142 -8982
rect 13366 -8880 13400 -8878
rect 13366 -8912 13400 -8880
rect 13366 -8982 13400 -8950
rect 13366 -8984 13400 -8982
rect 13560 -8880 13594 -8878
rect 13560 -8912 13594 -8880
rect 13560 -8982 13594 -8950
rect 13560 -8984 13594 -8982
rect 13818 -8880 13852 -8878
rect 13818 -8912 13852 -8880
rect 13818 -8982 13852 -8950
rect 13818 -8984 13852 -8982
rect 13932 -8844 13966 -8820
rect 18290 -8470 18324 -8460
rect 18290 -8494 18324 -8470
rect 18290 -8538 18324 -8532
rect 18290 -8566 18324 -8538
rect 18290 -8606 18324 -8604
rect 18290 -8638 18324 -8606
rect 18290 -8708 18324 -8676
rect 18290 -8710 18324 -8708
rect 18290 -8776 18324 -8748
rect 18290 -8782 18324 -8776
rect 13932 -8854 13966 -8844
rect 13932 -8912 13966 -8892
rect 13932 -8926 13966 -8912
rect 13932 -8980 13966 -8964
rect 13932 -8998 13966 -8980
rect 9573 -9070 9607 -9036
rect 5421 -9112 5423 -9078
rect 5423 -9112 5455 -9078
rect 5493 -9112 5525 -9078
rect 5525 -9112 5527 -9078
rect 5873 -9112 5875 -9078
rect 5875 -9112 5907 -9078
rect 5945 -9112 5977 -9078
rect 5977 -9112 5979 -9078
rect 6131 -9112 6133 -9078
rect 6133 -9112 6165 -9078
rect 6203 -9112 6235 -9078
rect 6235 -9112 6237 -9078
rect 6389 -9112 6391 -9078
rect 6391 -9112 6423 -9078
rect 6461 -9112 6493 -9078
rect 6493 -9112 6495 -9078
rect 6647 -9112 6649 -9078
rect 6649 -9112 6681 -9078
rect 6719 -9112 6751 -9078
rect 6751 -9112 6753 -9078
rect 7099 -9112 7101 -9078
rect 7101 -9112 7133 -9078
rect 7171 -9112 7203 -9078
rect 7203 -9112 7205 -9078
rect 7357 -9112 7359 -9078
rect 7359 -9112 7391 -9078
rect 7429 -9112 7461 -9078
rect 7461 -9112 7463 -9078
rect 7615 -9112 7617 -9078
rect 7617 -9112 7649 -9078
rect 7687 -9112 7719 -9078
rect 7719 -9112 7721 -9078
rect 8067 -9112 8069 -9078
rect 8069 -9112 8101 -9078
rect 8139 -9112 8171 -9078
rect 8171 -9112 8173 -9078
rect 8325 -9112 8327 -9078
rect 8327 -9112 8359 -9078
rect 8397 -9112 8429 -9078
rect 8429 -9112 8431 -9078
rect 8583 -9112 8585 -9078
rect 8585 -9112 8617 -9078
rect 8655 -9112 8687 -9078
rect 8687 -9112 8689 -9078
rect 8841 -9112 8843 -9078
rect 8843 -9112 8875 -9078
rect 8913 -9112 8945 -9078
rect 8945 -9112 8947 -9078
rect 9293 -9112 9295 -9078
rect 9295 -9112 9327 -9078
rect 9365 -9112 9397 -9078
rect 9397 -9112 9399 -9078
rect 14046 -8880 14080 -8878
rect 14046 -8912 14080 -8880
rect 14046 -8982 14080 -8950
rect 14046 -8984 14080 -8982
rect 14304 -8880 14338 -8878
rect 14304 -8912 14338 -8880
rect 14304 -8982 14338 -8950
rect 14304 -8984 14338 -8982
rect 14497 -8880 14531 -8878
rect 14497 -8912 14531 -8880
rect 14497 -8982 14531 -8950
rect 14497 -8984 14531 -8982
rect 14755 -8880 14789 -8878
rect 14755 -8912 14789 -8880
rect 14755 -8982 14789 -8950
rect 14755 -8984 14789 -8982
rect 15013 -8880 15047 -8878
rect 15013 -8912 15047 -8880
rect 15013 -8982 15047 -8950
rect 15013 -8984 15047 -8982
rect 15271 -8880 15305 -8878
rect 15271 -8912 15305 -8880
rect 15271 -8982 15305 -8950
rect 15271 -8984 15305 -8982
rect 15529 -8880 15563 -8878
rect 15529 -8912 15563 -8880
rect 15529 -8982 15563 -8950
rect 15529 -8984 15563 -8982
rect 15723 -8880 15757 -8878
rect 15723 -8912 15757 -8880
rect 15723 -8982 15757 -8950
rect 15723 -8984 15757 -8982
rect 15981 -8880 16015 -8878
rect 15981 -8912 16015 -8880
rect 15981 -8982 16015 -8950
rect 15981 -8984 16015 -8982
rect 16239 -8880 16273 -8878
rect 16239 -8912 16273 -8880
rect 16239 -8982 16273 -8950
rect 16239 -8984 16273 -8982
rect 16497 -8880 16531 -8878
rect 16497 -8912 16531 -8880
rect 16497 -8982 16531 -8950
rect 16497 -8984 16531 -8982
rect 16691 -8880 16725 -8878
rect 16691 -8912 16725 -8880
rect 16691 -8982 16725 -8950
rect 16691 -8984 16725 -8982
rect 16949 -8880 16983 -8878
rect 16949 -8912 16983 -8880
rect 16949 -8982 16983 -8950
rect 16949 -8984 16983 -8982
rect 17207 -8880 17241 -8878
rect 17207 -8912 17241 -8880
rect 17207 -8982 17241 -8950
rect 17207 -8984 17241 -8982
rect 17465 -8880 17499 -8878
rect 17465 -8912 17499 -8880
rect 17465 -8982 17499 -8950
rect 17465 -8984 17499 -8982
rect 17723 -8880 17757 -8878
rect 17723 -8912 17757 -8880
rect 17723 -8982 17757 -8950
rect 17723 -8984 17757 -8982
rect 17917 -8880 17951 -8878
rect 17917 -8912 17951 -8880
rect 17917 -8982 17951 -8950
rect 17917 -8984 17951 -8982
rect 18175 -8880 18209 -8878
rect 18175 -8912 18209 -8880
rect 18175 -8982 18209 -8950
rect 18175 -8984 18209 -8982
rect 18290 -8844 18324 -8820
rect 18290 -8854 18324 -8844
rect 18290 -8912 18324 -8892
rect 18290 -8926 18324 -8912
rect 18290 -8980 18324 -8964
rect 18290 -8998 18324 -8980
rect 13932 -9070 13966 -9036
rect 9781 -9112 9783 -9078
rect 9783 -9112 9815 -9078
rect 9853 -9112 9885 -9078
rect 9885 -9112 9887 -9078
rect 10233 -9112 10235 -9078
rect 10235 -9112 10267 -9078
rect 10305 -9112 10337 -9078
rect 10337 -9112 10339 -9078
rect 10491 -9112 10493 -9078
rect 10493 -9112 10525 -9078
rect 10563 -9112 10595 -9078
rect 10595 -9112 10597 -9078
rect 10749 -9112 10751 -9078
rect 10751 -9112 10783 -9078
rect 10821 -9112 10853 -9078
rect 10853 -9112 10855 -9078
rect 11007 -9112 11009 -9078
rect 11009 -9112 11041 -9078
rect 11079 -9112 11111 -9078
rect 11111 -9112 11113 -9078
rect 11459 -9112 11461 -9078
rect 11461 -9112 11493 -9078
rect 11531 -9112 11563 -9078
rect 11563 -9112 11565 -9078
rect 11717 -9112 11719 -9078
rect 11719 -9112 11751 -9078
rect 11789 -9112 11821 -9078
rect 11821 -9112 11823 -9078
rect 11975 -9112 11977 -9078
rect 11977 -9112 12009 -9078
rect 12047 -9112 12079 -9078
rect 12079 -9112 12081 -9078
rect 12427 -9112 12429 -9078
rect 12429 -9112 12461 -9078
rect 12499 -9112 12531 -9078
rect 12531 -9112 12533 -9078
rect 12685 -9112 12687 -9078
rect 12687 -9112 12719 -9078
rect 12757 -9112 12789 -9078
rect 12789 -9112 12791 -9078
rect 12943 -9112 12945 -9078
rect 12945 -9112 12977 -9078
rect 13015 -9112 13047 -9078
rect 13047 -9112 13049 -9078
rect 13201 -9112 13203 -9078
rect 13203 -9112 13235 -9078
rect 13273 -9112 13305 -9078
rect 13305 -9112 13307 -9078
rect 13653 -9112 13655 -9078
rect 13655 -9112 13687 -9078
rect 13725 -9112 13757 -9078
rect 13757 -9112 13759 -9078
rect 18290 -9070 18324 -9036
rect 14139 -9112 14141 -9078
rect 14141 -9112 14173 -9078
rect 14211 -9112 14243 -9078
rect 14243 -9112 14245 -9078
rect 14590 -9112 14592 -9078
rect 14592 -9112 14624 -9078
rect 14662 -9112 14694 -9078
rect 14694 -9112 14696 -9078
rect 14848 -9112 14850 -9078
rect 14850 -9112 14882 -9078
rect 14920 -9112 14952 -9078
rect 14952 -9112 14954 -9078
rect 15106 -9112 15108 -9078
rect 15108 -9112 15140 -9078
rect 15178 -9112 15210 -9078
rect 15210 -9112 15212 -9078
rect 15364 -9112 15366 -9078
rect 15366 -9112 15398 -9078
rect 15436 -9112 15468 -9078
rect 15468 -9112 15470 -9078
rect 15816 -9112 15818 -9078
rect 15818 -9112 15850 -9078
rect 15888 -9112 15920 -9078
rect 15920 -9112 15922 -9078
rect 16074 -9112 16076 -9078
rect 16076 -9112 16108 -9078
rect 16146 -9112 16178 -9078
rect 16178 -9112 16180 -9078
rect 16332 -9112 16334 -9078
rect 16334 -9112 16366 -9078
rect 16404 -9112 16436 -9078
rect 16436 -9112 16438 -9078
rect 16784 -9112 16786 -9078
rect 16786 -9112 16818 -9078
rect 16856 -9112 16888 -9078
rect 16888 -9112 16890 -9078
rect 17042 -9112 17044 -9078
rect 17044 -9112 17076 -9078
rect 17114 -9112 17146 -9078
rect 17146 -9112 17148 -9078
rect 17300 -9112 17302 -9078
rect 17302 -9112 17334 -9078
rect 17372 -9112 17404 -9078
rect 17404 -9112 17406 -9078
rect 17558 -9112 17560 -9078
rect 17560 -9112 17592 -9078
rect 17630 -9112 17662 -9078
rect 17662 -9112 17664 -9078
rect 18010 -9112 18012 -9078
rect 18012 -9112 18044 -9078
rect 18082 -9112 18114 -9078
rect 18114 -9112 18116 -9078
rect 930 -9226 964 -9192
rect 1002 -9226 1011 -9192
rect 1011 -9226 1036 -9192
rect 1074 -9226 1079 -9192
rect 1079 -9226 1108 -9192
rect 1146 -9226 1147 -9192
rect 1147 -9226 1180 -9192
rect 1218 -9226 1249 -9192
rect 1249 -9226 1252 -9192
rect 1290 -9226 1317 -9192
rect 1317 -9226 1324 -9192
rect 1362 -9226 1385 -9192
rect 1385 -9226 1396 -9192
rect 1434 -9226 1453 -9192
rect 1453 -9226 1468 -9192
rect 1506 -9226 1521 -9192
rect 1521 -9226 1540 -9192
rect 1578 -9226 1589 -9192
rect 1589 -9226 1612 -9192
rect 1650 -9226 1657 -9192
rect 1657 -9226 1684 -9192
rect 1722 -9226 1725 -9192
rect 1725 -9226 1756 -9192
rect 1794 -9226 1827 -9192
rect 1827 -9226 1828 -9192
rect 1866 -9226 1895 -9192
rect 1895 -9226 1900 -9192
rect 1938 -9226 1963 -9192
rect 1963 -9226 1972 -9192
rect 2010 -9226 2031 -9192
rect 2031 -9226 2044 -9192
rect 2082 -9226 2099 -9192
rect 2099 -9226 2116 -9192
rect 2154 -9226 2167 -9192
rect 2167 -9226 2188 -9192
rect 2226 -9226 2235 -9192
rect 2235 -9226 2260 -9192
rect 2298 -9226 2303 -9192
rect 2303 -9226 2332 -9192
rect 2370 -9226 2371 -9192
rect 2371 -9226 2404 -9192
rect 2442 -9226 2473 -9192
rect 2473 -9226 2476 -9192
rect 2514 -9226 2541 -9192
rect 2541 -9226 2548 -9192
rect 2586 -9226 2609 -9192
rect 2609 -9226 2620 -9192
rect 2658 -9226 2677 -9192
rect 2677 -9226 2692 -9192
rect 2730 -9226 2745 -9192
rect 2745 -9226 2764 -9192
rect 2802 -9226 2813 -9192
rect 2813 -9226 2836 -9192
rect 2874 -9226 2881 -9192
rect 2881 -9226 2908 -9192
rect 2946 -9226 2949 -9192
rect 2949 -9226 2980 -9192
rect 3018 -9226 3051 -9192
rect 3051 -9226 3052 -9192
rect 3090 -9226 3119 -9192
rect 3119 -9226 3124 -9192
rect 3162 -9226 3187 -9192
rect 3187 -9226 3196 -9192
rect 3234 -9226 3255 -9192
rect 3255 -9226 3268 -9192
rect 3306 -9226 3323 -9192
rect 3323 -9226 3340 -9192
rect 3378 -9226 3391 -9192
rect 3391 -9226 3412 -9192
rect 3450 -9226 3459 -9192
rect 3459 -9226 3484 -9192
rect 3522 -9226 3527 -9192
rect 3527 -9226 3556 -9192
rect 3594 -9226 3595 -9192
rect 3595 -9226 3628 -9192
rect 3666 -9226 3697 -9192
rect 3697 -9226 3700 -9192
rect 3738 -9226 3765 -9192
rect 3765 -9226 3772 -9192
rect 3810 -9226 3833 -9192
rect 3833 -9226 3844 -9192
rect 3882 -9226 3901 -9192
rect 3901 -9226 3916 -9192
rect 3954 -9226 3969 -9192
rect 3969 -9226 3988 -9192
rect 4026 -9226 4037 -9192
rect 4037 -9226 4060 -9192
rect 4098 -9226 4105 -9192
rect 4105 -9226 4132 -9192
rect 4170 -9226 4173 -9192
rect 4173 -9226 4204 -9192
rect 4242 -9226 4275 -9192
rect 4275 -9226 4276 -9192
rect 4314 -9226 4343 -9192
rect 4343 -9226 4348 -9192
rect 4386 -9226 4411 -9192
rect 4411 -9226 4420 -9192
rect 4458 -9226 4479 -9192
rect 4479 -9226 4492 -9192
rect 4530 -9226 4547 -9192
rect 4547 -9226 4564 -9192
rect 4602 -9226 4615 -9192
rect 4615 -9226 4636 -9192
rect 4674 -9226 4683 -9192
rect 4683 -9226 4708 -9192
rect 4746 -9226 4751 -9192
rect 4751 -9226 4780 -9192
rect 4818 -9226 4819 -9192
rect 4819 -9226 4852 -9192
rect 4890 -9226 4921 -9192
rect 4921 -9226 4924 -9192
rect 4962 -9226 4989 -9192
rect 4989 -9226 4996 -9192
rect 5034 -9226 5057 -9192
rect 5057 -9226 5068 -9192
rect 5106 -9226 5140 -9192
rect 5323 -9226 5357 -9192
rect 5395 -9226 5406 -9192
rect 5406 -9226 5429 -9192
rect 5467 -9226 5474 -9192
rect 5474 -9226 5501 -9192
rect 5539 -9226 5542 -9192
rect 5542 -9226 5573 -9192
rect 5611 -9226 5644 -9192
rect 5644 -9226 5645 -9192
rect 5683 -9226 5712 -9192
rect 5712 -9226 5717 -9192
rect 5755 -9226 5780 -9192
rect 5780 -9226 5789 -9192
rect 5827 -9226 5848 -9192
rect 5848 -9226 5861 -9192
rect 5899 -9226 5916 -9192
rect 5916 -9226 5933 -9192
rect 5971 -9226 5984 -9192
rect 5984 -9226 6005 -9192
rect 6043 -9226 6052 -9192
rect 6052 -9226 6077 -9192
rect 6115 -9226 6120 -9192
rect 6120 -9226 6149 -9192
rect 6187 -9226 6188 -9192
rect 6188 -9226 6221 -9192
rect 6259 -9226 6290 -9192
rect 6290 -9226 6293 -9192
rect 6331 -9226 6358 -9192
rect 6358 -9226 6365 -9192
rect 6403 -9226 6426 -9192
rect 6426 -9226 6437 -9192
rect 6475 -9226 6494 -9192
rect 6494 -9226 6509 -9192
rect 6547 -9226 6562 -9192
rect 6562 -9226 6581 -9192
rect 6619 -9226 6630 -9192
rect 6630 -9226 6653 -9192
rect 6691 -9226 6698 -9192
rect 6698 -9226 6725 -9192
rect 6763 -9226 6766 -9192
rect 6766 -9226 6797 -9192
rect 6835 -9226 6868 -9192
rect 6868 -9226 6869 -9192
rect 6907 -9226 6936 -9192
rect 6936 -9226 6941 -9192
rect 6979 -9226 7004 -9192
rect 7004 -9226 7013 -9192
rect 7051 -9226 7072 -9192
rect 7072 -9226 7085 -9192
rect 7123 -9226 7140 -9192
rect 7140 -9226 7157 -9192
rect 7195 -9226 7208 -9192
rect 7208 -9226 7229 -9192
rect 7267 -9226 7276 -9192
rect 7276 -9226 7301 -9192
rect 7339 -9226 7344 -9192
rect 7344 -9226 7373 -9192
rect 7411 -9226 7412 -9192
rect 7412 -9226 7445 -9192
rect 7483 -9226 7514 -9192
rect 7514 -9226 7517 -9192
rect 7555 -9226 7582 -9192
rect 7582 -9226 7589 -9192
rect 7627 -9226 7650 -9192
rect 7650 -9226 7661 -9192
rect 7699 -9226 7718 -9192
rect 7718 -9226 7733 -9192
rect 7771 -9226 7786 -9192
rect 7786 -9226 7805 -9192
rect 7843 -9226 7854 -9192
rect 7854 -9226 7877 -9192
rect 7915 -9226 7922 -9192
rect 7922 -9226 7949 -9192
rect 7987 -9226 7990 -9192
rect 7990 -9226 8021 -9192
rect 8059 -9226 8092 -9192
rect 8092 -9226 8093 -9192
rect 8131 -9226 8160 -9192
rect 8160 -9226 8165 -9192
rect 8203 -9226 8228 -9192
rect 8228 -9226 8237 -9192
rect 8275 -9226 8296 -9192
rect 8296 -9226 8309 -9192
rect 8347 -9226 8364 -9192
rect 8364 -9226 8381 -9192
rect 8419 -9226 8432 -9192
rect 8432 -9226 8453 -9192
rect 8491 -9226 8500 -9192
rect 8500 -9226 8525 -9192
rect 8563 -9226 8568 -9192
rect 8568 -9226 8597 -9192
rect 8635 -9226 8636 -9192
rect 8636 -9226 8669 -9192
rect 8707 -9226 8738 -9192
rect 8738 -9226 8741 -9192
rect 8779 -9226 8806 -9192
rect 8806 -9226 8813 -9192
rect 8851 -9226 8874 -9192
rect 8874 -9226 8885 -9192
rect 8923 -9226 8942 -9192
rect 8942 -9226 8957 -9192
rect 8995 -9226 9010 -9192
rect 9010 -9226 9029 -9192
rect 9067 -9226 9078 -9192
rect 9078 -9226 9101 -9192
rect 9139 -9226 9146 -9192
rect 9146 -9226 9173 -9192
rect 9211 -9226 9214 -9192
rect 9214 -9226 9245 -9192
rect 9283 -9226 9316 -9192
rect 9316 -9226 9317 -9192
rect 9355 -9226 9384 -9192
rect 9384 -9226 9389 -9192
rect 9427 -9226 9452 -9192
rect 9452 -9226 9461 -9192
rect 9499 -9226 9533 -9192
rect 9647 -9226 9681 -9192
rect 9719 -9226 9728 -9192
rect 9728 -9226 9753 -9192
rect 9791 -9226 9796 -9192
rect 9796 -9226 9825 -9192
rect 9863 -9226 9864 -9192
rect 9864 -9226 9897 -9192
rect 9935 -9226 9966 -9192
rect 9966 -9226 9969 -9192
rect 10007 -9226 10034 -9192
rect 10034 -9226 10041 -9192
rect 10079 -9226 10102 -9192
rect 10102 -9226 10113 -9192
rect 10151 -9226 10170 -9192
rect 10170 -9226 10185 -9192
rect 10223 -9226 10238 -9192
rect 10238 -9226 10257 -9192
rect 10295 -9226 10306 -9192
rect 10306 -9226 10329 -9192
rect 10367 -9226 10374 -9192
rect 10374 -9226 10401 -9192
rect 10439 -9226 10442 -9192
rect 10442 -9226 10473 -9192
rect 10511 -9226 10544 -9192
rect 10544 -9226 10545 -9192
rect 10583 -9226 10612 -9192
rect 10612 -9226 10617 -9192
rect 10655 -9226 10680 -9192
rect 10680 -9226 10689 -9192
rect 10727 -9226 10748 -9192
rect 10748 -9226 10761 -9192
rect 10799 -9226 10816 -9192
rect 10816 -9226 10833 -9192
rect 10871 -9226 10884 -9192
rect 10884 -9226 10905 -9192
rect 10943 -9226 10952 -9192
rect 10952 -9226 10977 -9192
rect 11015 -9226 11020 -9192
rect 11020 -9226 11049 -9192
rect 11087 -9226 11088 -9192
rect 11088 -9226 11121 -9192
rect 11159 -9226 11190 -9192
rect 11190 -9226 11193 -9192
rect 11231 -9226 11258 -9192
rect 11258 -9226 11265 -9192
rect 11303 -9226 11326 -9192
rect 11326 -9226 11337 -9192
rect 11375 -9226 11394 -9192
rect 11394 -9226 11409 -9192
rect 11447 -9226 11462 -9192
rect 11462 -9226 11481 -9192
rect 11519 -9226 11530 -9192
rect 11530 -9226 11553 -9192
rect 11591 -9226 11598 -9192
rect 11598 -9226 11625 -9192
rect 11663 -9226 11666 -9192
rect 11666 -9226 11697 -9192
rect 11735 -9226 11768 -9192
rect 11768 -9226 11769 -9192
rect 11807 -9226 11836 -9192
rect 11836 -9226 11841 -9192
rect 11879 -9226 11904 -9192
rect 11904 -9226 11913 -9192
rect 11951 -9226 11972 -9192
rect 11972 -9226 11985 -9192
rect 12023 -9226 12040 -9192
rect 12040 -9226 12057 -9192
rect 12095 -9226 12108 -9192
rect 12108 -9226 12129 -9192
rect 12167 -9226 12176 -9192
rect 12176 -9226 12201 -9192
rect 12239 -9226 12244 -9192
rect 12244 -9226 12273 -9192
rect 12311 -9226 12312 -9192
rect 12312 -9226 12345 -9192
rect 12383 -9226 12414 -9192
rect 12414 -9226 12417 -9192
rect 12455 -9226 12482 -9192
rect 12482 -9226 12489 -9192
rect 12527 -9226 12550 -9192
rect 12550 -9226 12561 -9192
rect 12599 -9226 12618 -9192
rect 12618 -9226 12633 -9192
rect 12671 -9226 12686 -9192
rect 12686 -9226 12705 -9192
rect 12743 -9226 12754 -9192
rect 12754 -9226 12777 -9192
rect 12815 -9226 12822 -9192
rect 12822 -9226 12849 -9192
rect 12887 -9226 12890 -9192
rect 12890 -9226 12921 -9192
rect 12959 -9226 12992 -9192
rect 12992 -9226 12993 -9192
rect 13031 -9226 13060 -9192
rect 13060 -9226 13065 -9192
rect 13103 -9226 13128 -9192
rect 13128 -9226 13137 -9192
rect 13175 -9226 13196 -9192
rect 13196 -9226 13209 -9192
rect 13247 -9226 13264 -9192
rect 13264 -9226 13281 -9192
rect 13319 -9226 13332 -9192
rect 13332 -9226 13353 -9192
rect 13391 -9226 13400 -9192
rect 13400 -9226 13425 -9192
rect 13463 -9226 13468 -9192
rect 13468 -9226 13497 -9192
rect 13535 -9226 13536 -9192
rect 13536 -9226 13569 -9192
rect 13607 -9226 13638 -9192
rect 13638 -9226 13641 -9192
rect 13679 -9226 13706 -9192
rect 13706 -9226 13713 -9192
rect 13751 -9226 13774 -9192
rect 13774 -9226 13785 -9192
rect 13823 -9226 13857 -9192
rect 14040 -9226 14074 -9192
rect 14112 -9226 14123 -9192
rect 14123 -9226 14146 -9192
rect 14184 -9226 14191 -9192
rect 14191 -9226 14218 -9192
rect 14256 -9226 14259 -9192
rect 14259 -9226 14290 -9192
rect 14328 -9226 14361 -9192
rect 14361 -9226 14362 -9192
rect 14400 -9226 14429 -9192
rect 14429 -9226 14434 -9192
rect 14472 -9226 14497 -9192
rect 14497 -9226 14506 -9192
rect 14544 -9226 14565 -9192
rect 14565 -9226 14578 -9192
rect 14616 -9226 14633 -9192
rect 14633 -9226 14650 -9192
rect 14688 -9226 14701 -9192
rect 14701 -9226 14722 -9192
rect 14760 -9226 14769 -9192
rect 14769 -9226 14794 -9192
rect 14832 -9226 14837 -9192
rect 14837 -9226 14866 -9192
rect 14904 -9226 14905 -9192
rect 14905 -9226 14938 -9192
rect 14976 -9226 15007 -9192
rect 15007 -9226 15010 -9192
rect 15048 -9226 15075 -9192
rect 15075 -9226 15082 -9192
rect 15120 -9226 15143 -9192
rect 15143 -9226 15154 -9192
rect 15192 -9226 15211 -9192
rect 15211 -9226 15226 -9192
rect 15264 -9226 15279 -9192
rect 15279 -9226 15298 -9192
rect 15336 -9226 15347 -9192
rect 15347 -9226 15370 -9192
rect 15408 -9226 15415 -9192
rect 15415 -9226 15442 -9192
rect 15480 -9226 15483 -9192
rect 15483 -9226 15514 -9192
rect 15552 -9226 15585 -9192
rect 15585 -9226 15586 -9192
rect 15624 -9226 15653 -9192
rect 15653 -9226 15658 -9192
rect 15696 -9226 15721 -9192
rect 15721 -9226 15730 -9192
rect 15768 -9226 15789 -9192
rect 15789 -9226 15802 -9192
rect 15840 -9226 15857 -9192
rect 15857 -9226 15874 -9192
rect 15912 -9226 15925 -9192
rect 15925 -9226 15946 -9192
rect 15984 -9226 15993 -9192
rect 15993 -9226 16018 -9192
rect 16056 -9226 16061 -9192
rect 16061 -9226 16090 -9192
rect 16128 -9226 16129 -9192
rect 16129 -9226 16162 -9192
rect 16200 -9226 16231 -9192
rect 16231 -9226 16234 -9192
rect 16272 -9226 16299 -9192
rect 16299 -9226 16306 -9192
rect 16344 -9226 16367 -9192
rect 16367 -9226 16378 -9192
rect 16416 -9226 16435 -9192
rect 16435 -9226 16450 -9192
rect 16488 -9226 16503 -9192
rect 16503 -9226 16522 -9192
rect 16560 -9226 16571 -9192
rect 16571 -9226 16594 -9192
rect 16632 -9226 16639 -9192
rect 16639 -9226 16666 -9192
rect 16704 -9226 16707 -9192
rect 16707 -9226 16738 -9192
rect 16776 -9226 16809 -9192
rect 16809 -9226 16810 -9192
rect 16848 -9226 16877 -9192
rect 16877 -9226 16882 -9192
rect 16920 -9226 16945 -9192
rect 16945 -9226 16954 -9192
rect 16992 -9226 17013 -9192
rect 17013 -9226 17026 -9192
rect 17064 -9226 17081 -9192
rect 17081 -9226 17098 -9192
rect 17136 -9226 17149 -9192
rect 17149 -9226 17170 -9192
rect 17208 -9226 17217 -9192
rect 17217 -9226 17242 -9192
rect 17280 -9226 17285 -9192
rect 17285 -9226 17314 -9192
rect 17352 -9226 17353 -9192
rect 17353 -9226 17386 -9192
rect 17424 -9226 17455 -9192
rect 17455 -9226 17458 -9192
rect 17496 -9226 17523 -9192
rect 17523 -9226 17530 -9192
rect 17568 -9226 17591 -9192
rect 17591 -9226 17602 -9192
rect 17640 -9226 17659 -9192
rect 17659 -9226 17674 -9192
rect 17712 -9226 17727 -9192
rect 17727 -9226 17746 -9192
rect 17784 -9226 17795 -9192
rect 17795 -9226 17818 -9192
rect 17856 -9226 17863 -9192
rect 17863 -9226 17890 -9192
rect 17928 -9226 17931 -9192
rect 17931 -9226 17962 -9192
rect 18000 -9226 18033 -9192
rect 18033 -9226 18034 -9192
rect 18072 -9226 18101 -9192
rect 18101 -9226 18106 -9192
rect 18144 -9226 18169 -9192
rect 18169 -9226 18178 -9192
rect 18216 -9226 18250 -9192
<< metal1 >>
rect 831 463 18349 488
rect 831 429 930 463
rect 964 429 1002 463
rect 1036 429 1074 463
rect 1108 429 1146 463
rect 1180 429 1218 463
rect 1252 429 1290 463
rect 1324 429 1362 463
rect 1396 429 1434 463
rect 1468 429 1506 463
rect 1540 429 1578 463
rect 1612 429 1650 463
rect 1684 429 1722 463
rect 1756 429 1794 463
rect 1828 429 1866 463
rect 1900 429 1938 463
rect 1972 429 2010 463
rect 2044 429 2082 463
rect 2116 429 2154 463
rect 2188 429 2226 463
rect 2260 429 2298 463
rect 2332 429 2370 463
rect 2404 429 2442 463
rect 2476 429 2514 463
rect 2548 429 2586 463
rect 2620 429 2658 463
rect 2692 429 2730 463
rect 2764 429 2802 463
rect 2836 429 2874 463
rect 2908 429 2946 463
rect 2980 429 3018 463
rect 3052 429 3090 463
rect 3124 429 3162 463
rect 3196 429 3234 463
rect 3268 429 3306 463
rect 3340 429 3378 463
rect 3412 429 3450 463
rect 3484 429 3522 463
rect 3556 429 3594 463
rect 3628 429 3666 463
rect 3700 429 3738 463
rect 3772 429 3810 463
rect 3844 429 3882 463
rect 3916 429 3954 463
rect 3988 429 4026 463
rect 4060 429 4098 463
rect 4132 429 4170 463
rect 4204 429 4242 463
rect 4276 429 4314 463
rect 4348 429 4386 463
rect 4420 429 4458 463
rect 4492 429 4530 463
rect 4564 429 4602 463
rect 4636 429 4674 463
rect 4708 429 4746 463
rect 4780 429 4818 463
rect 4852 429 4890 463
rect 4924 429 4962 463
rect 4996 429 5034 463
rect 5068 429 5106 463
rect 5140 429 5323 463
rect 5357 429 5395 463
rect 5429 429 5467 463
rect 5501 429 5539 463
rect 5573 429 5611 463
rect 5645 429 5683 463
rect 5717 429 5755 463
rect 5789 429 5827 463
rect 5861 429 5899 463
rect 5933 429 5971 463
rect 6005 429 6043 463
rect 6077 429 6115 463
rect 6149 429 6187 463
rect 6221 429 6259 463
rect 6293 429 6331 463
rect 6365 429 6403 463
rect 6437 429 6475 463
rect 6509 429 6547 463
rect 6581 429 6619 463
rect 6653 429 6691 463
rect 6725 429 6763 463
rect 6797 429 6835 463
rect 6869 429 6907 463
rect 6941 429 6979 463
rect 7013 429 7051 463
rect 7085 429 7123 463
rect 7157 429 7195 463
rect 7229 429 7267 463
rect 7301 429 7339 463
rect 7373 429 7411 463
rect 7445 429 7483 463
rect 7517 429 7555 463
rect 7589 429 7627 463
rect 7661 429 7699 463
rect 7733 429 7771 463
rect 7805 429 7843 463
rect 7877 429 7915 463
rect 7949 429 7987 463
rect 8021 429 8059 463
rect 8093 429 8131 463
rect 8165 429 8203 463
rect 8237 429 8275 463
rect 8309 429 8347 463
rect 8381 429 8419 463
rect 8453 429 8491 463
rect 8525 429 8563 463
rect 8597 429 8635 463
rect 8669 429 8707 463
rect 8741 429 8779 463
rect 8813 429 8851 463
rect 8885 429 8923 463
rect 8957 429 8995 463
rect 9029 429 9067 463
rect 9101 429 9139 463
rect 9173 429 9211 463
rect 9245 429 9283 463
rect 9317 429 9355 463
rect 9389 429 9427 463
rect 9461 429 9499 463
rect 9533 429 9647 463
rect 9681 429 9719 463
rect 9753 429 9791 463
rect 9825 429 9863 463
rect 9897 429 9935 463
rect 9969 429 10007 463
rect 10041 429 10079 463
rect 10113 429 10151 463
rect 10185 429 10223 463
rect 10257 429 10295 463
rect 10329 429 10367 463
rect 10401 429 10439 463
rect 10473 429 10511 463
rect 10545 429 10583 463
rect 10617 429 10655 463
rect 10689 429 10727 463
rect 10761 429 10799 463
rect 10833 429 10871 463
rect 10905 429 10943 463
rect 10977 429 11015 463
rect 11049 429 11087 463
rect 11121 429 11159 463
rect 11193 429 11231 463
rect 11265 429 11303 463
rect 11337 429 11375 463
rect 11409 429 11447 463
rect 11481 429 11519 463
rect 11553 429 11591 463
rect 11625 429 11663 463
rect 11697 429 11735 463
rect 11769 429 11807 463
rect 11841 429 11879 463
rect 11913 429 11951 463
rect 11985 429 12023 463
rect 12057 429 12095 463
rect 12129 429 12167 463
rect 12201 429 12239 463
rect 12273 429 12311 463
rect 12345 429 12383 463
rect 12417 429 12455 463
rect 12489 429 12527 463
rect 12561 429 12599 463
rect 12633 429 12671 463
rect 12705 429 12743 463
rect 12777 429 12815 463
rect 12849 429 12887 463
rect 12921 429 12959 463
rect 12993 429 13031 463
rect 13065 429 13103 463
rect 13137 429 13175 463
rect 13209 429 13247 463
rect 13281 429 13319 463
rect 13353 429 13391 463
rect 13425 429 13463 463
rect 13497 429 13535 463
rect 13569 429 13607 463
rect 13641 429 13679 463
rect 13713 429 13751 463
rect 13785 429 13823 463
rect 13857 429 14040 463
rect 14074 429 14112 463
rect 14146 429 14184 463
rect 14218 429 14256 463
rect 14290 429 14328 463
rect 14362 429 14400 463
rect 14434 429 14472 463
rect 14506 429 14544 463
rect 14578 429 14616 463
rect 14650 429 14688 463
rect 14722 429 14760 463
rect 14794 429 14832 463
rect 14866 429 14904 463
rect 14938 429 14976 463
rect 15010 429 15048 463
rect 15082 429 15120 463
rect 15154 429 15192 463
rect 15226 429 15264 463
rect 15298 429 15336 463
rect 15370 429 15408 463
rect 15442 429 15480 463
rect 15514 429 15552 463
rect 15586 429 15624 463
rect 15658 429 15696 463
rect 15730 429 15768 463
rect 15802 429 15840 463
rect 15874 429 15912 463
rect 15946 429 15984 463
rect 16018 429 16056 463
rect 16090 429 16128 463
rect 16162 429 16200 463
rect 16234 429 16272 463
rect 16306 429 16344 463
rect 16378 429 16416 463
rect 16450 429 16488 463
rect 16522 429 16560 463
rect 16594 429 16632 463
rect 16666 429 16704 463
rect 16738 429 16776 463
rect 16810 429 16848 463
rect 16882 429 16920 463
rect 16954 429 16992 463
rect 17026 429 17064 463
rect 17098 429 17136 463
rect 17170 429 17208 463
rect 17242 429 17280 463
rect 17314 429 17352 463
rect 17386 429 17424 463
rect 17458 429 17496 463
rect 17530 429 17568 463
rect 17602 429 17640 463
rect 17674 429 17712 463
rect 17746 429 17784 463
rect 17818 429 17856 463
rect 17890 429 17928 463
rect 17962 429 18000 463
rect 18034 429 18072 463
rect 18106 429 18144 463
rect 18178 429 18216 463
rect 18250 429 18349 463
rect 831 349 18349 429
rect 831 315 1064 349
rect 1098 315 1136 349
rect 1170 315 1516 349
rect 1550 315 1588 349
rect 1622 315 1774 349
rect 1808 315 1846 349
rect 1880 315 2032 349
rect 2066 315 2104 349
rect 2138 315 2290 349
rect 2324 315 2362 349
rect 2396 315 2742 349
rect 2776 315 2814 349
rect 2848 315 3000 349
rect 3034 315 3072 349
rect 3106 315 3258 349
rect 3292 315 3330 349
rect 3364 315 3710 349
rect 3744 315 3782 349
rect 3816 315 3968 349
rect 4002 315 4040 349
rect 4074 315 4226 349
rect 4260 315 4298 349
rect 4332 315 4484 349
rect 4518 315 4556 349
rect 4590 315 4935 349
rect 4969 315 5007 349
rect 5041 315 5421 349
rect 5455 315 5493 349
rect 5527 315 5873 349
rect 5907 315 5945 349
rect 5979 315 6131 349
rect 6165 315 6203 349
rect 6237 315 6389 349
rect 6423 315 6461 349
rect 6495 315 6647 349
rect 6681 315 6719 349
rect 6753 315 7099 349
rect 7133 315 7171 349
rect 7205 315 7357 349
rect 7391 315 7429 349
rect 7463 315 7615 349
rect 7649 315 7687 349
rect 7721 315 8067 349
rect 8101 315 8139 349
rect 8173 315 8325 349
rect 8359 315 8397 349
rect 8431 315 8583 349
rect 8617 315 8655 349
rect 8689 315 8841 349
rect 8875 315 8913 349
rect 8947 315 9293 349
rect 9327 315 9365 349
rect 9399 315 9781 349
rect 9815 315 9853 349
rect 9887 315 10233 349
rect 10267 315 10305 349
rect 10339 315 10491 349
rect 10525 315 10563 349
rect 10597 315 10749 349
rect 10783 315 10821 349
rect 10855 315 11007 349
rect 11041 315 11079 349
rect 11113 315 11459 349
rect 11493 315 11531 349
rect 11565 315 11717 349
rect 11751 315 11789 349
rect 11823 315 11975 349
rect 12009 315 12047 349
rect 12081 315 12427 349
rect 12461 315 12499 349
rect 12533 315 12685 349
rect 12719 315 12757 349
rect 12791 315 12943 349
rect 12977 315 13015 349
rect 13049 315 13201 349
rect 13235 315 13273 349
rect 13307 315 13653 349
rect 13687 315 13725 349
rect 13759 315 14139 349
rect 14173 315 14211 349
rect 14245 315 14590 349
rect 14624 315 14662 349
rect 14696 315 14848 349
rect 14882 315 14920 349
rect 14954 315 15106 349
rect 15140 315 15178 349
rect 15212 315 15364 349
rect 15398 315 15436 349
rect 15470 315 15816 349
rect 15850 315 15888 349
rect 15922 315 16074 349
rect 16108 315 16146 349
rect 16180 315 16332 349
rect 16366 315 16404 349
rect 16438 315 16784 349
rect 16818 315 16856 349
rect 16890 315 17042 349
rect 17076 315 17114 349
rect 17148 315 17300 349
rect 17334 315 17372 349
rect 17406 315 17558 349
rect 17592 315 17630 349
rect 17664 315 18010 349
rect 18044 315 18082 349
rect 18116 315 18349 349
rect 831 309 18349 315
rect 833 306 1269 309
rect 833 272 856 306
rect 890 272 1269 306
rect 833 234 1269 272
rect 833 200 856 234
rect 890 221 1269 234
rect 890 200 971 221
rect 833 187 971 200
rect 1005 187 1229 221
rect 1263 187 1269 221
rect 833 162 1269 187
rect 833 128 856 162
rect 890 149 1269 162
rect 890 128 971 149
rect 833 115 971 128
rect 1005 115 1229 149
rect 1263 115 1269 149
rect 833 90 1269 115
rect 833 56 856 90
rect 890 56 1269 90
rect 1417 221 1463 309
rect 1417 187 1423 221
rect 1457 187 1463 221
rect 1417 149 1463 187
rect 1417 115 1423 149
rect 1457 115 1463 149
rect 1417 68 1463 115
rect 1675 221 1721 309
rect 1675 187 1681 221
rect 1715 187 1721 221
rect 1675 149 1721 187
rect 1675 115 1681 149
rect 1715 115 1721 149
rect 1675 68 1721 115
rect 1933 221 1979 309
rect 1933 187 1939 221
rect 1973 187 1979 221
rect 1933 149 1979 187
rect 1933 115 1939 149
rect 1973 115 1979 149
rect 1933 68 1979 115
rect 2191 221 2237 309
rect 2191 187 2197 221
rect 2231 187 2237 221
rect 2191 149 2237 187
rect 2191 115 2197 149
rect 2231 115 2237 149
rect 2191 68 2237 115
rect 2449 221 2495 309
rect 2449 187 2455 221
rect 2489 187 2495 221
rect 2449 149 2495 187
rect 2449 115 2455 149
rect 2489 115 2495 149
rect 2449 68 2495 115
rect 2643 221 2689 309
rect 2643 187 2649 221
rect 2683 187 2689 221
rect 2643 149 2689 187
rect 2643 115 2649 149
rect 2683 115 2689 149
rect 2643 68 2689 115
rect 2901 221 2947 309
rect 2901 187 2907 221
rect 2941 187 2947 221
rect 2901 149 2947 187
rect 2901 115 2907 149
rect 2941 115 2947 149
rect 2901 68 2947 115
rect 3159 221 3205 309
rect 3159 187 3165 221
rect 3199 187 3205 221
rect 3159 149 3205 187
rect 3159 115 3165 149
rect 3199 115 3205 149
rect 3159 68 3205 115
rect 3417 221 3463 309
rect 3417 187 3423 221
rect 3457 187 3463 221
rect 3417 149 3463 187
rect 3417 115 3423 149
rect 3457 115 3463 149
rect 3417 68 3463 115
rect 3611 221 3657 309
rect 3611 187 3617 221
rect 3651 187 3657 221
rect 3611 149 3657 187
rect 3611 115 3617 149
rect 3651 115 3657 149
rect 3611 68 3657 115
rect 3869 221 3915 309
rect 3869 187 3875 221
rect 3909 187 3915 221
rect 3869 149 3915 187
rect 3869 115 3875 149
rect 3909 115 3915 149
rect 3869 68 3915 115
rect 4127 221 4173 309
rect 4127 187 4133 221
rect 4167 187 4173 221
rect 4127 149 4173 187
rect 4127 115 4133 149
rect 4167 115 4173 149
rect 4127 68 4173 115
rect 4385 221 4431 309
rect 4385 187 4391 221
rect 4425 187 4431 221
rect 4385 149 4431 187
rect 4385 115 4391 149
rect 4425 115 4431 149
rect 4385 68 4431 115
rect 4643 221 4689 309
rect 4643 187 4649 221
rect 4683 187 4689 221
rect 4643 149 4689 187
rect 4643 115 4649 149
rect 4683 115 4689 149
rect 4643 68 4689 115
rect 4836 306 5626 309
rect 4836 272 5214 306
rect 5248 272 5626 306
rect 4836 234 5626 272
rect 4836 221 5214 234
rect 4836 187 4842 221
rect 4876 187 5100 221
rect 5134 200 5214 221
rect 5248 221 5626 234
rect 5248 200 5328 221
rect 5134 187 5328 200
rect 5362 187 5586 221
rect 5620 187 5626 221
rect 4836 162 5626 187
rect 4836 149 5214 162
rect 4836 115 4842 149
rect 4876 115 5100 149
rect 5134 128 5214 149
rect 5248 149 5626 162
rect 5248 128 5328 149
rect 5134 115 5328 128
rect 5362 115 5586 149
rect 5620 115 5626 149
rect 4836 90 5626 115
rect 833 18 1269 56
rect 833 -16 856 18
rect 890 -16 1269 18
rect 4836 56 5214 90
rect 5248 56 5626 90
rect 5774 221 5820 309
rect 5774 187 5780 221
rect 5814 187 5820 221
rect 5774 149 5820 187
rect 5774 115 5780 149
rect 5814 115 5820 149
rect 5774 68 5820 115
rect 6032 221 6078 309
rect 6032 187 6038 221
rect 6072 187 6078 221
rect 6032 149 6078 187
rect 6032 115 6038 149
rect 6072 115 6078 149
rect 6032 68 6078 115
rect 6290 221 6336 309
rect 6290 187 6296 221
rect 6330 187 6336 221
rect 6290 149 6336 187
rect 6290 115 6296 149
rect 6330 115 6336 149
rect 6290 68 6336 115
rect 6548 221 6594 309
rect 6548 187 6554 221
rect 6588 187 6594 221
rect 6548 149 6594 187
rect 6548 115 6554 149
rect 6588 115 6594 149
rect 6548 68 6594 115
rect 6806 221 6852 309
rect 6806 187 6812 221
rect 6846 187 6852 221
rect 6806 149 6852 187
rect 6806 115 6812 149
rect 6846 115 6852 149
rect 6806 68 6852 115
rect 7000 221 7046 309
rect 7000 187 7006 221
rect 7040 187 7046 221
rect 7000 149 7046 187
rect 7000 115 7006 149
rect 7040 115 7046 149
rect 7000 68 7046 115
rect 7258 221 7304 309
rect 7258 187 7264 221
rect 7298 187 7304 221
rect 7258 149 7304 187
rect 7258 115 7264 149
rect 7298 115 7304 149
rect 7258 68 7304 115
rect 7516 221 7562 309
rect 7516 187 7522 221
rect 7556 187 7562 221
rect 7516 149 7562 187
rect 7516 115 7522 149
rect 7556 115 7562 149
rect 7516 68 7562 115
rect 7774 221 7820 309
rect 7774 187 7780 221
rect 7814 187 7820 221
rect 7774 149 7820 187
rect 7774 115 7780 149
rect 7814 115 7820 149
rect 7774 68 7820 115
rect 7968 221 8014 309
rect 7968 187 7974 221
rect 8008 187 8014 221
rect 7968 149 8014 187
rect 7968 115 7974 149
rect 8008 115 8014 149
rect 7968 68 8014 115
rect 8226 221 8272 309
rect 8226 187 8232 221
rect 8266 187 8272 221
rect 8226 149 8272 187
rect 8226 115 8232 149
rect 8266 115 8272 149
rect 8226 68 8272 115
rect 8484 221 8530 309
rect 8484 187 8490 221
rect 8524 187 8530 221
rect 8484 149 8530 187
rect 8484 115 8490 149
rect 8524 115 8530 149
rect 8484 68 8530 115
rect 8742 221 8788 309
rect 8742 187 8748 221
rect 8782 187 8788 221
rect 8742 149 8788 187
rect 8742 115 8748 149
rect 8782 115 8788 149
rect 8742 68 8788 115
rect 9000 221 9046 309
rect 9000 187 9006 221
rect 9040 187 9046 221
rect 9000 149 9046 187
rect 9000 115 9006 149
rect 9040 115 9046 149
rect 9000 68 9046 115
rect 9194 306 9986 309
rect 9194 272 9573 306
rect 9607 272 9986 306
rect 9194 234 9986 272
rect 9194 221 9573 234
rect 9194 187 9200 221
rect 9234 187 9458 221
rect 9492 200 9573 221
rect 9607 221 9986 234
rect 9607 200 9688 221
rect 9492 187 9688 200
rect 9722 187 9946 221
rect 9980 187 9986 221
rect 9194 162 9986 187
rect 9194 149 9573 162
rect 9194 115 9200 149
rect 9234 115 9458 149
rect 9492 128 9573 149
rect 9607 149 9986 162
rect 9607 128 9688 149
rect 9492 115 9688 128
rect 9722 115 9946 149
rect 9980 115 9986 149
rect 9194 90 9986 115
rect 4836 18 5626 56
rect 833 -54 1269 -16
rect 833 -88 856 -54
rect 890 -88 1269 -54
rect 2827 -12 3023 -4
rect 2827 -64 2834 -12
rect 2886 -64 2898 -12
rect 2950 -64 2962 -12
rect 3014 -64 3023 -12
rect 2827 -74 3023 -64
rect 3344 -12 3540 -4
rect 3344 -64 3351 -12
rect 3403 -64 3415 -12
rect 3467 -64 3479 -12
rect 3531 -64 3540 -12
rect 3344 -74 3540 -64
rect 4836 -16 5214 18
rect 5248 -16 5626 18
rect 9194 56 9573 90
rect 9607 56 9986 90
rect 10134 221 10180 309
rect 10134 187 10140 221
rect 10174 187 10180 221
rect 10134 149 10180 187
rect 10134 115 10140 149
rect 10174 115 10180 149
rect 10134 68 10180 115
rect 10392 221 10438 309
rect 10392 187 10398 221
rect 10432 187 10438 221
rect 10392 149 10438 187
rect 10392 115 10398 149
rect 10432 115 10438 149
rect 10392 68 10438 115
rect 10650 221 10696 309
rect 10650 187 10656 221
rect 10690 187 10696 221
rect 10650 149 10696 187
rect 10650 115 10656 149
rect 10690 115 10696 149
rect 10650 68 10696 115
rect 10908 221 10954 309
rect 10908 187 10914 221
rect 10948 187 10954 221
rect 10908 149 10954 187
rect 10908 115 10914 149
rect 10948 115 10954 149
rect 10908 68 10954 115
rect 11166 221 11212 309
rect 11166 187 11172 221
rect 11206 187 11212 221
rect 11166 149 11212 187
rect 11166 115 11172 149
rect 11206 115 11212 149
rect 11166 68 11212 115
rect 11360 221 11406 309
rect 11360 187 11366 221
rect 11400 187 11406 221
rect 11360 149 11406 187
rect 11360 115 11366 149
rect 11400 115 11406 149
rect 11360 68 11406 115
rect 11618 221 11664 309
rect 11618 187 11624 221
rect 11658 187 11664 221
rect 11618 149 11664 187
rect 11618 115 11624 149
rect 11658 115 11664 149
rect 11618 68 11664 115
rect 11876 221 11922 309
rect 11876 187 11882 221
rect 11916 187 11922 221
rect 11876 149 11922 187
rect 11876 115 11882 149
rect 11916 115 11922 149
rect 11876 68 11922 115
rect 12134 221 12180 309
rect 12134 187 12140 221
rect 12174 187 12180 221
rect 12134 149 12180 187
rect 12134 115 12140 149
rect 12174 115 12180 149
rect 12134 68 12180 115
rect 12328 221 12374 309
rect 12328 187 12334 221
rect 12368 187 12374 221
rect 12328 149 12374 187
rect 12328 115 12334 149
rect 12368 115 12374 149
rect 12328 68 12374 115
rect 12586 221 12632 309
rect 12586 187 12592 221
rect 12626 187 12632 221
rect 12586 149 12632 187
rect 12586 115 12592 149
rect 12626 115 12632 149
rect 12586 68 12632 115
rect 12844 221 12890 309
rect 12844 187 12850 221
rect 12884 187 12890 221
rect 12844 149 12890 187
rect 12844 115 12850 149
rect 12884 115 12890 149
rect 12844 68 12890 115
rect 13102 221 13148 309
rect 13102 187 13108 221
rect 13142 187 13148 221
rect 13102 149 13148 187
rect 13102 115 13108 149
rect 13142 115 13148 149
rect 13102 68 13148 115
rect 13360 221 13406 309
rect 13360 187 13366 221
rect 13400 187 13406 221
rect 13360 149 13406 187
rect 13360 115 13366 149
rect 13400 115 13406 149
rect 13360 68 13406 115
rect 13554 306 14344 309
rect 13554 272 13932 306
rect 13966 272 14344 306
rect 13554 234 14344 272
rect 13554 221 13932 234
rect 13554 187 13560 221
rect 13594 187 13818 221
rect 13852 200 13932 221
rect 13966 221 14344 234
rect 13966 200 14046 221
rect 13852 187 14046 200
rect 14080 187 14304 221
rect 14338 187 14344 221
rect 13554 162 14344 187
rect 13554 149 13932 162
rect 13554 115 13560 149
rect 13594 115 13818 149
rect 13852 128 13932 149
rect 13966 149 14344 162
rect 13966 128 14046 149
rect 13852 115 14046 128
rect 14080 115 14304 149
rect 14338 115 14344 149
rect 13554 90 14344 115
rect 9194 18 9986 56
rect 4836 -54 5626 -16
rect 833 -126 1269 -88
rect 833 -160 856 -126
rect 890 -160 1269 -126
rect 833 -198 1269 -160
rect 833 -232 856 -198
rect 890 -232 1269 -198
rect 833 -270 1269 -232
rect 1339 -181 1535 -173
rect 1339 -233 1348 -181
rect 1400 -233 1412 -181
rect 1464 -233 1476 -181
rect 1528 -233 1535 -181
rect 1339 -243 1535 -233
rect 1856 -181 2052 -173
rect 1856 -233 1865 -181
rect 1917 -233 1929 -181
rect 1981 -233 1993 -181
rect 2045 -233 2052 -181
rect 1856 -243 2052 -233
rect 2373 -181 2569 -173
rect 2373 -233 2382 -181
rect 2434 -233 2446 -181
rect 2498 -233 2510 -181
rect 2562 -233 2569 -181
rect 2373 -243 2569 -233
rect 833 -304 856 -270
rect 890 -304 1269 -270
rect 833 -342 1269 -304
rect 833 -376 856 -342
rect 890 -376 1269 -342
rect 833 -414 1269 -376
rect 833 -448 856 -414
rect 890 -448 1269 -414
rect 833 -486 1269 -448
rect 833 -520 856 -486
rect 890 -520 1269 -486
rect 833 -558 1269 -520
rect 833 -592 856 -558
rect 890 -592 1269 -558
rect 833 -630 1269 -592
rect 833 -664 856 -630
rect 890 -664 1269 -630
rect 833 -702 1269 -664
rect 833 -736 856 -702
rect 890 -723 1269 -702
rect 890 -736 971 -723
rect 833 -757 971 -736
rect 1005 -757 1229 -723
rect 1263 -757 1269 -723
rect 833 -774 1269 -757
rect 833 -808 856 -774
rect 890 -795 1269 -774
rect 890 -808 971 -795
rect 833 -829 971 -808
rect 1005 -829 1229 -795
rect 1263 -829 1269 -795
rect 833 -846 1269 -829
rect 833 -880 856 -846
rect 890 -880 1269 -846
rect 1417 -723 1463 -243
rect 1598 -512 1794 -504
rect 1598 -564 1607 -512
rect 1659 -564 1671 -512
rect 1723 -564 1735 -512
rect 1787 -564 1794 -512
rect 1598 -574 1794 -564
rect 1417 -757 1423 -723
rect 1457 -757 1463 -723
rect 1417 -795 1463 -757
rect 1417 -829 1423 -795
rect 1457 -829 1463 -795
rect 1417 -876 1463 -829
rect 1675 -723 1721 -574
rect 1675 -757 1681 -723
rect 1715 -757 1721 -723
rect 1675 -795 1721 -757
rect 1675 -829 1681 -795
rect 1715 -829 1721 -795
rect 1675 -876 1721 -829
rect 1933 -723 1979 -243
rect 2116 -512 2312 -504
rect 2116 -564 2125 -512
rect 2177 -564 2189 -512
rect 2241 -564 2253 -512
rect 2305 -564 2312 -512
rect 2116 -574 2312 -564
rect 1933 -757 1939 -723
rect 1973 -757 1979 -723
rect 1933 -795 1979 -757
rect 1933 -829 1939 -795
rect 1973 -829 1979 -795
rect 1933 -876 1979 -829
rect 2191 -723 2237 -574
rect 2191 -757 2197 -723
rect 2231 -757 2237 -723
rect 2191 -795 2237 -757
rect 2191 -829 2197 -795
rect 2231 -829 2237 -795
rect 2191 -876 2237 -829
rect 2449 -723 2495 -243
rect 2570 -344 2766 -336
rect 2570 -396 2577 -344
rect 2629 -396 2641 -344
rect 2693 -396 2705 -344
rect 2757 -396 2766 -344
rect 2570 -406 2766 -396
rect 2449 -757 2455 -723
rect 2489 -757 2495 -723
rect 2449 -795 2495 -757
rect 2449 -829 2455 -795
rect 2489 -829 2495 -795
rect 2449 -876 2495 -829
rect 2643 -723 2689 -406
rect 2643 -757 2649 -723
rect 2683 -757 2689 -723
rect 2643 -795 2689 -757
rect 2643 -829 2649 -795
rect 2683 -829 2689 -795
rect 2643 -876 2689 -829
rect 2901 -723 2947 -74
rect 3087 -344 3283 -336
rect 3087 -396 3094 -344
rect 3146 -396 3158 -344
rect 3210 -396 3222 -344
rect 3274 -396 3283 -344
rect 3087 -406 3283 -396
rect 2901 -757 2907 -723
rect 2941 -757 2947 -723
rect 2901 -795 2947 -757
rect 2901 -829 2907 -795
rect 2941 -829 2947 -795
rect 2901 -876 2947 -829
rect 3159 -723 3205 -406
rect 3159 -757 3165 -723
rect 3199 -757 3205 -723
rect 3159 -795 3205 -757
rect 3159 -829 3165 -795
rect 3199 -829 3205 -795
rect 3159 -876 3205 -829
rect 3417 -723 3463 -74
rect 4836 -88 5214 -54
rect 5248 -88 5626 -54
rect 6922 -12 7118 -4
rect 6922 -64 6931 -12
rect 6983 -64 6995 -12
rect 7047 -64 7059 -12
rect 7111 -64 7118 -12
rect 6922 -74 7118 -64
rect 7440 -12 7636 -4
rect 7440 -64 7449 -12
rect 7501 -64 7513 -12
rect 7565 -64 7577 -12
rect 7629 -64 7636 -12
rect 7440 -74 7636 -64
rect 9194 -16 9573 18
rect 9607 -16 9986 18
rect 13554 56 13932 90
rect 13966 56 14344 90
rect 14491 221 14537 309
rect 14491 187 14497 221
rect 14531 187 14537 221
rect 14491 149 14537 187
rect 14491 115 14497 149
rect 14531 115 14537 149
rect 14491 68 14537 115
rect 14749 221 14795 309
rect 14749 187 14755 221
rect 14789 187 14795 221
rect 14749 149 14795 187
rect 14749 115 14755 149
rect 14789 115 14795 149
rect 14749 68 14795 115
rect 15007 221 15053 309
rect 15007 187 15013 221
rect 15047 187 15053 221
rect 15007 149 15053 187
rect 15007 115 15013 149
rect 15047 115 15053 149
rect 15007 68 15053 115
rect 15265 221 15311 309
rect 15265 187 15271 221
rect 15305 187 15311 221
rect 15265 149 15311 187
rect 15265 115 15271 149
rect 15305 115 15311 149
rect 15265 68 15311 115
rect 15523 221 15569 309
rect 15523 187 15529 221
rect 15563 187 15569 221
rect 15523 149 15569 187
rect 15523 115 15529 149
rect 15563 115 15569 149
rect 15523 68 15569 115
rect 15717 221 15763 309
rect 15717 187 15723 221
rect 15757 187 15763 221
rect 15717 149 15763 187
rect 15717 115 15723 149
rect 15757 115 15763 149
rect 15717 68 15763 115
rect 15975 221 16021 309
rect 15975 187 15981 221
rect 16015 187 16021 221
rect 15975 149 16021 187
rect 15975 115 15981 149
rect 16015 115 16021 149
rect 15975 68 16021 115
rect 16233 221 16279 309
rect 16233 187 16239 221
rect 16273 187 16279 221
rect 16233 149 16279 187
rect 16233 115 16239 149
rect 16273 115 16279 149
rect 16233 68 16279 115
rect 16491 221 16537 309
rect 16491 187 16497 221
rect 16531 187 16537 221
rect 16491 149 16537 187
rect 16491 115 16497 149
rect 16531 115 16537 149
rect 16491 68 16537 115
rect 16685 221 16731 309
rect 16685 187 16691 221
rect 16725 187 16731 221
rect 16685 149 16731 187
rect 16685 115 16691 149
rect 16725 115 16731 149
rect 16685 68 16731 115
rect 16943 221 16989 309
rect 16943 187 16949 221
rect 16983 187 16989 221
rect 16943 149 16989 187
rect 16943 115 16949 149
rect 16983 115 16989 149
rect 16943 68 16989 115
rect 17201 221 17247 309
rect 17201 187 17207 221
rect 17241 187 17247 221
rect 17201 149 17247 187
rect 17201 115 17207 149
rect 17241 115 17247 149
rect 17201 68 17247 115
rect 17459 221 17505 309
rect 17459 187 17465 221
rect 17499 187 17505 221
rect 17459 149 17505 187
rect 17459 115 17465 149
rect 17499 115 17505 149
rect 17459 68 17505 115
rect 17717 221 17763 309
rect 17717 187 17723 221
rect 17757 187 17763 221
rect 17717 149 17763 187
rect 17717 115 17723 149
rect 17757 115 17763 149
rect 17717 68 17763 115
rect 17911 306 18347 309
rect 17911 272 18290 306
rect 18324 272 18347 306
rect 17911 234 18347 272
rect 17911 221 18290 234
rect 17911 187 17917 221
rect 17951 187 18175 221
rect 18209 200 18290 221
rect 18324 200 18347 234
rect 18209 187 18347 200
rect 17911 162 18347 187
rect 17911 149 18290 162
rect 17911 115 17917 149
rect 17951 115 18175 149
rect 18209 128 18290 149
rect 18324 128 18347 162
rect 18209 115 18347 128
rect 17911 90 18347 115
rect 13554 18 14344 56
rect 9194 -54 9986 -16
rect 4836 -126 5626 -88
rect 4836 -160 5214 -126
rect 5248 -160 5626 -126
rect 3534 -181 3730 -173
rect 3534 -233 3543 -181
rect 3595 -233 3607 -181
rect 3659 -233 3671 -181
rect 3723 -233 3730 -181
rect 3534 -243 3730 -233
rect 4051 -181 4247 -173
rect 4051 -233 4060 -181
rect 4112 -233 4124 -181
rect 4176 -233 4188 -181
rect 4240 -233 4247 -181
rect 4051 -243 4247 -233
rect 4566 -181 4762 -173
rect 4566 -233 4575 -181
rect 4627 -233 4639 -181
rect 4691 -233 4703 -181
rect 4755 -233 4762 -181
rect 4566 -243 4762 -233
rect 4836 -198 5626 -160
rect 4836 -232 5214 -198
rect 5248 -232 5626 -198
rect 3417 -757 3423 -723
rect 3457 -757 3463 -723
rect 3417 -795 3463 -757
rect 3417 -829 3423 -795
rect 3457 -829 3463 -795
rect 3417 -876 3463 -829
rect 3611 -723 3657 -243
rect 3793 -512 3989 -504
rect 3793 -564 3802 -512
rect 3854 -564 3866 -512
rect 3918 -564 3930 -512
rect 3982 -564 3989 -512
rect 3793 -574 3989 -564
rect 3611 -757 3617 -723
rect 3651 -757 3657 -723
rect 3611 -795 3657 -757
rect 3611 -829 3617 -795
rect 3651 -829 3657 -795
rect 3611 -876 3657 -829
rect 3869 -723 3915 -574
rect 3869 -757 3875 -723
rect 3909 -757 3915 -723
rect 3869 -795 3915 -757
rect 3869 -829 3875 -795
rect 3909 -829 3915 -795
rect 3869 -876 3915 -829
rect 4127 -723 4173 -243
rect 4310 -512 4506 -504
rect 4310 -564 4319 -512
rect 4371 -564 4383 -512
rect 4435 -564 4447 -512
rect 4499 -564 4506 -512
rect 4310 -574 4506 -564
rect 4127 -757 4133 -723
rect 4167 -757 4173 -723
rect 4127 -795 4173 -757
rect 4127 -829 4133 -795
rect 4167 -829 4173 -795
rect 4127 -876 4173 -829
rect 4385 -723 4431 -574
rect 4385 -757 4391 -723
rect 4425 -757 4431 -723
rect 4385 -795 4431 -757
rect 4385 -829 4391 -795
rect 4425 -829 4431 -795
rect 4385 -876 4431 -829
rect 4643 -723 4689 -243
rect 4643 -757 4649 -723
rect 4683 -757 4689 -723
rect 4643 -795 4689 -757
rect 4643 -829 4649 -795
rect 4683 -829 4689 -795
rect 4643 -876 4689 -829
rect 4836 -270 5626 -232
rect 5701 -181 5897 -173
rect 5701 -233 5708 -181
rect 5760 -233 5772 -181
rect 5824 -233 5836 -181
rect 5888 -233 5897 -181
rect 5701 -243 5897 -233
rect 6216 -181 6412 -173
rect 6216 -233 6223 -181
rect 6275 -233 6287 -181
rect 6339 -233 6351 -181
rect 6403 -233 6412 -181
rect 6216 -243 6412 -233
rect 6733 -181 6929 -173
rect 6733 -233 6740 -181
rect 6792 -233 6804 -181
rect 6856 -233 6868 -181
rect 6920 -233 6929 -181
rect 6733 -243 6929 -233
rect 4836 -304 5214 -270
rect 5248 -304 5626 -270
rect 4836 -342 5626 -304
rect 4836 -376 5214 -342
rect 5248 -376 5626 -342
rect 4836 -414 5626 -376
rect 4836 -448 5214 -414
rect 5248 -448 5626 -414
rect 4836 -486 5626 -448
rect 4836 -520 5214 -486
rect 5248 -520 5626 -486
rect 4836 -558 5626 -520
rect 4836 -592 5214 -558
rect 5248 -592 5626 -558
rect 4836 -630 5626 -592
rect 4836 -664 5214 -630
rect 5248 -664 5626 -630
rect 4836 -702 5626 -664
rect 4836 -723 5214 -702
rect 4836 -757 4842 -723
rect 4876 -757 5100 -723
rect 5134 -736 5214 -723
rect 5248 -723 5626 -702
rect 5248 -736 5328 -723
rect 5134 -757 5328 -736
rect 5362 -757 5586 -723
rect 5620 -757 5626 -723
rect 4836 -774 5626 -757
rect 4836 -795 5214 -774
rect 4836 -829 4842 -795
rect 4876 -829 5100 -795
rect 5134 -808 5214 -795
rect 5248 -795 5626 -774
rect 5248 -808 5328 -795
rect 5134 -829 5328 -808
rect 5362 -829 5586 -795
rect 5620 -829 5626 -795
rect 4836 -846 5626 -829
rect 833 -918 1269 -880
rect 4836 -880 5214 -846
rect 5248 -880 5626 -846
rect 5774 -723 5820 -243
rect 5957 -512 6153 -504
rect 5957 -564 5964 -512
rect 6016 -564 6028 -512
rect 6080 -564 6092 -512
rect 6144 -564 6153 -512
rect 5957 -574 6153 -564
rect 5774 -757 5780 -723
rect 5814 -757 5820 -723
rect 5774 -795 5820 -757
rect 5774 -829 5780 -795
rect 5814 -829 5820 -795
rect 5774 -876 5820 -829
rect 6032 -723 6078 -574
rect 6032 -757 6038 -723
rect 6072 -757 6078 -723
rect 6032 -795 6078 -757
rect 6032 -829 6038 -795
rect 6072 -829 6078 -795
rect 6032 -876 6078 -829
rect 6290 -723 6336 -243
rect 6474 -512 6670 -504
rect 6474 -564 6481 -512
rect 6533 -564 6545 -512
rect 6597 -564 6609 -512
rect 6661 -564 6670 -512
rect 6474 -574 6670 -564
rect 6290 -757 6296 -723
rect 6330 -757 6336 -723
rect 6290 -795 6336 -757
rect 6290 -829 6296 -795
rect 6330 -829 6336 -795
rect 6290 -876 6336 -829
rect 6548 -723 6594 -574
rect 6548 -757 6554 -723
rect 6588 -757 6594 -723
rect 6548 -795 6594 -757
rect 6548 -829 6554 -795
rect 6588 -829 6594 -795
rect 6548 -876 6594 -829
rect 6806 -723 6852 -243
rect 6806 -757 6812 -723
rect 6846 -757 6852 -723
rect 6806 -795 6852 -757
rect 6806 -829 6812 -795
rect 6846 -829 6852 -795
rect 6806 -876 6852 -829
rect 7000 -723 7046 -74
rect 7180 -344 7376 -336
rect 7180 -396 7189 -344
rect 7241 -396 7253 -344
rect 7305 -396 7317 -344
rect 7369 -396 7376 -344
rect 7180 -406 7376 -396
rect 7000 -757 7006 -723
rect 7040 -757 7046 -723
rect 7000 -795 7046 -757
rect 7000 -829 7006 -795
rect 7040 -829 7046 -795
rect 7000 -876 7046 -829
rect 7258 -723 7304 -406
rect 7258 -757 7264 -723
rect 7298 -757 7304 -723
rect 7258 -795 7304 -757
rect 7258 -829 7264 -795
rect 7298 -829 7304 -795
rect 7258 -876 7304 -829
rect 7516 -723 7562 -74
rect 9194 -88 9573 -54
rect 9607 -88 9986 -54
rect 11544 -12 11740 -4
rect 11544 -64 11551 -12
rect 11603 -64 11615 -12
rect 11667 -64 11679 -12
rect 11731 -64 11740 -12
rect 11544 -74 11740 -64
rect 12062 -12 12258 -4
rect 12062 -64 12069 -12
rect 12121 -64 12133 -12
rect 12185 -64 12197 -12
rect 12249 -64 12258 -12
rect 12062 -74 12258 -64
rect 13554 -16 13932 18
rect 13966 -16 14344 18
rect 17911 56 18290 90
rect 18324 56 18347 90
rect 17911 18 18347 56
rect 13554 -54 14344 -16
rect 9194 -126 9986 -88
rect 9194 -160 9573 -126
rect 9607 -160 9986 -126
rect 7894 -181 8090 -173
rect 7894 -233 7901 -181
rect 7953 -233 7965 -181
rect 8017 -233 8029 -181
rect 8081 -233 8090 -181
rect 7894 -243 8090 -233
rect 8410 -181 8606 -173
rect 8410 -233 8417 -181
rect 8469 -233 8481 -181
rect 8533 -233 8545 -181
rect 8597 -233 8606 -181
rect 8410 -243 8606 -233
rect 8928 -181 9124 -173
rect 8928 -233 8935 -181
rect 8987 -233 8999 -181
rect 9051 -233 9063 -181
rect 9115 -233 9124 -181
rect 8928 -243 9124 -233
rect 9194 -198 9986 -160
rect 9194 -232 9573 -198
rect 9607 -232 9986 -198
rect 7697 -344 7893 -336
rect 7697 -396 7706 -344
rect 7758 -396 7770 -344
rect 7822 -396 7834 -344
rect 7886 -396 7893 -344
rect 7697 -406 7893 -396
rect 7516 -757 7522 -723
rect 7556 -757 7562 -723
rect 7516 -795 7562 -757
rect 7516 -829 7522 -795
rect 7556 -829 7562 -795
rect 7516 -876 7562 -829
rect 7774 -723 7820 -406
rect 7774 -757 7780 -723
rect 7814 -757 7820 -723
rect 7774 -795 7820 -757
rect 7774 -829 7780 -795
rect 7814 -829 7820 -795
rect 7774 -876 7820 -829
rect 7968 -723 8014 -243
rect 8151 -512 8347 -504
rect 8151 -564 8158 -512
rect 8210 -564 8222 -512
rect 8274 -564 8286 -512
rect 8338 -564 8347 -512
rect 8151 -574 8347 -564
rect 7968 -757 7974 -723
rect 8008 -757 8014 -723
rect 7968 -795 8014 -757
rect 7968 -829 7974 -795
rect 8008 -829 8014 -795
rect 7968 -876 8014 -829
rect 8226 -723 8272 -574
rect 8226 -757 8232 -723
rect 8266 -757 8272 -723
rect 8226 -795 8272 -757
rect 8226 -829 8232 -795
rect 8266 -829 8272 -795
rect 8226 -876 8272 -829
rect 8484 -723 8530 -243
rect 8668 -512 8864 -504
rect 8668 -564 8675 -512
rect 8727 -564 8739 -512
rect 8791 -564 8803 -512
rect 8855 -564 8864 -512
rect 8668 -574 8864 -564
rect 8484 -757 8490 -723
rect 8524 -757 8530 -723
rect 8484 -795 8530 -757
rect 8484 -829 8490 -795
rect 8524 -829 8530 -795
rect 8484 -876 8530 -829
rect 8742 -723 8788 -574
rect 8742 -757 8748 -723
rect 8782 -757 8788 -723
rect 8742 -795 8788 -757
rect 8742 -829 8748 -795
rect 8782 -829 8788 -795
rect 8742 -876 8788 -829
rect 9000 -723 9046 -243
rect 9000 -757 9006 -723
rect 9040 -757 9046 -723
rect 9000 -795 9046 -757
rect 9000 -829 9006 -795
rect 9040 -829 9046 -795
rect 9000 -876 9046 -829
rect 9194 -270 9986 -232
rect 10056 -181 10252 -173
rect 10056 -233 10065 -181
rect 10117 -233 10129 -181
rect 10181 -233 10193 -181
rect 10245 -233 10252 -181
rect 10056 -243 10252 -233
rect 10574 -181 10770 -173
rect 10574 -233 10583 -181
rect 10635 -233 10647 -181
rect 10699 -233 10711 -181
rect 10763 -233 10770 -181
rect 10574 -243 10770 -233
rect 11090 -181 11286 -173
rect 11090 -233 11099 -181
rect 11151 -233 11163 -181
rect 11215 -233 11227 -181
rect 11279 -233 11286 -181
rect 11090 -243 11286 -233
rect 9194 -304 9573 -270
rect 9607 -304 9986 -270
rect 9194 -342 9986 -304
rect 9194 -376 9573 -342
rect 9607 -376 9986 -342
rect 9194 -414 9986 -376
rect 9194 -448 9573 -414
rect 9607 -448 9986 -414
rect 9194 -486 9986 -448
rect 9194 -520 9573 -486
rect 9607 -520 9986 -486
rect 9194 -558 9986 -520
rect 9194 -592 9573 -558
rect 9607 -592 9986 -558
rect 9194 -630 9986 -592
rect 9194 -664 9573 -630
rect 9607 -664 9986 -630
rect 9194 -702 9986 -664
rect 9194 -723 9573 -702
rect 9194 -757 9200 -723
rect 9234 -757 9458 -723
rect 9492 -736 9573 -723
rect 9607 -723 9986 -702
rect 9607 -736 9688 -723
rect 9492 -757 9688 -736
rect 9722 -757 9946 -723
rect 9980 -757 9986 -723
rect 9194 -774 9986 -757
rect 9194 -795 9573 -774
rect 9194 -829 9200 -795
rect 9234 -829 9458 -795
rect 9492 -808 9573 -795
rect 9607 -795 9986 -774
rect 9607 -808 9688 -795
rect 9492 -829 9688 -808
rect 9722 -829 9946 -795
rect 9980 -829 9986 -795
rect 9194 -846 9986 -829
rect 833 -952 856 -918
rect 890 -923 1269 -918
rect 890 -952 1064 -923
rect 833 -957 1064 -952
rect 1098 -957 1136 -923
rect 1170 -957 1269 -923
rect 833 -990 1269 -957
rect 833 -1024 856 -990
rect 890 -1024 1269 -990
rect 1473 -923 2577 -917
rect 1473 -957 1516 -923
rect 1550 -936 1588 -923
rect 1622 -936 1774 -923
rect 1808 -936 1846 -923
rect 1880 -936 2032 -923
rect 2066 -936 2104 -923
rect 2138 -936 2290 -923
rect 2324 -936 2362 -923
rect 1473 -988 1523 -957
rect 1575 -988 1587 -936
rect 1639 -988 1651 -936
rect 1703 -988 1719 -936
rect 1771 -957 1774 -936
rect 1835 -957 1846 -936
rect 1771 -988 1783 -957
rect 1835 -988 1847 -957
rect 1899 -988 2009 -936
rect 2066 -957 2073 -936
rect 2061 -988 2073 -957
rect 2125 -988 2137 -957
rect 2189 -988 2205 -936
rect 2257 -988 2269 -936
rect 2324 -957 2333 -936
rect 2396 -957 2577 -923
rect 2321 -988 2333 -957
rect 2385 -988 2577 -957
rect 1473 -1006 2577 -988
rect 833 -1062 1269 -1024
rect 833 -1096 856 -1062
rect 890 -1096 1269 -1062
rect 833 -1134 1269 -1096
rect 833 -1168 856 -1134
rect 890 -1168 1269 -1134
rect 833 -1206 1269 -1168
rect 833 -1240 856 -1206
rect 890 -1240 1269 -1206
rect 833 -1278 1269 -1240
rect 833 -1312 856 -1278
rect 890 -1286 1269 -1278
rect 890 -1312 1064 -1286
rect 833 -1320 1064 -1312
rect 1098 -1320 1136 -1286
rect 1170 -1320 1269 -1286
rect 833 -1350 1269 -1320
rect 1473 -1074 2439 -1056
rect 1473 -1126 1523 -1074
rect 1575 -1126 1587 -1074
rect 1639 -1126 1651 -1074
rect 1703 -1126 1719 -1074
rect 1771 -1126 1783 -1074
rect 1835 -1126 1847 -1074
rect 1899 -1126 2009 -1074
rect 2061 -1126 2073 -1074
rect 2125 -1126 2137 -1074
rect 2189 -1126 2205 -1074
rect 2257 -1126 2269 -1074
rect 2321 -1126 2333 -1074
rect 2385 -1126 2439 -1074
rect 1473 -1252 2439 -1126
rect 1473 -1286 1523 -1252
rect 1473 -1320 1516 -1286
rect 1575 -1304 1587 -1252
rect 1639 -1304 1651 -1252
rect 1703 -1304 1719 -1252
rect 1771 -1286 1783 -1252
rect 1835 -1286 1847 -1252
rect 1771 -1304 1774 -1286
rect 1835 -1304 1846 -1286
rect 1899 -1304 2009 -1252
rect 2061 -1286 2073 -1252
rect 2125 -1286 2137 -1252
rect 2066 -1304 2073 -1286
rect 2189 -1304 2205 -1252
rect 2257 -1304 2269 -1252
rect 2321 -1286 2333 -1252
rect 2385 -1286 2439 -1252
rect 2324 -1304 2333 -1286
rect 1550 -1320 1588 -1304
rect 1622 -1320 1774 -1304
rect 1808 -1320 1846 -1304
rect 1880 -1320 2032 -1304
rect 2066 -1320 2104 -1304
rect 2138 -1320 2290 -1304
rect 2324 -1320 2362 -1304
rect 2396 -1320 2439 -1286
rect 1473 -1326 2439 -1320
rect 2516 -1238 2577 -1006
rect 2699 -923 3407 -917
rect 2699 -957 2742 -923
rect 2776 -957 2814 -923
rect 2848 -957 3000 -923
rect 3034 -957 3072 -923
rect 3106 -957 3258 -923
rect 3292 -957 3330 -923
rect 3364 -957 3407 -923
rect 2699 -1074 3407 -957
rect 2699 -1126 2733 -1074
rect 2785 -1126 2797 -1074
rect 2849 -1126 2861 -1074
rect 2913 -1126 2929 -1074
rect 2981 -1126 2993 -1074
rect 3045 -1126 3057 -1074
rect 3109 -1126 3121 -1074
rect 3173 -1126 3189 -1074
rect 3241 -1126 3253 -1074
rect 3305 -1126 3317 -1074
rect 3369 -1126 3407 -1074
rect 2699 -1144 3407 -1126
rect 3529 -923 4633 -917
rect 3529 -957 3710 -923
rect 3744 -936 3782 -923
rect 3816 -936 3968 -923
rect 4002 -936 4040 -923
rect 4074 -936 4226 -923
rect 4260 -936 4298 -923
rect 4332 -936 4484 -923
rect 4518 -936 4556 -923
rect 3773 -957 3782 -936
rect 3529 -988 3721 -957
rect 3773 -988 3785 -957
rect 3837 -988 3849 -936
rect 3901 -988 3917 -936
rect 4033 -957 4040 -936
rect 3969 -988 3981 -957
rect 4033 -988 4045 -957
rect 4097 -988 4207 -936
rect 4260 -957 4271 -936
rect 4332 -957 4335 -936
rect 4259 -988 4271 -957
rect 4323 -988 4335 -957
rect 4387 -988 4403 -936
rect 4455 -988 4467 -936
rect 4519 -988 4531 -936
rect 4590 -957 4633 -923
rect 4583 -988 4633 -957
rect 3529 -1006 4633 -988
rect 4836 -918 5626 -880
rect 9194 -880 9573 -846
rect 9607 -880 9986 -846
rect 10134 -723 10180 -243
rect 10316 -512 10512 -504
rect 10316 -564 10325 -512
rect 10377 -564 10389 -512
rect 10441 -564 10453 -512
rect 10505 -564 10512 -512
rect 10316 -574 10512 -564
rect 10134 -757 10140 -723
rect 10174 -757 10180 -723
rect 10134 -795 10180 -757
rect 10134 -829 10140 -795
rect 10174 -829 10180 -795
rect 10134 -876 10180 -829
rect 10392 -723 10438 -574
rect 10392 -757 10398 -723
rect 10432 -757 10438 -723
rect 10392 -795 10438 -757
rect 10392 -829 10398 -795
rect 10432 -829 10438 -795
rect 10392 -876 10438 -829
rect 10650 -723 10696 -243
rect 10833 -512 11029 -504
rect 10833 -564 10842 -512
rect 10894 -564 10906 -512
rect 10958 -564 10970 -512
rect 11022 -564 11029 -512
rect 10833 -574 11029 -564
rect 10650 -757 10656 -723
rect 10690 -757 10696 -723
rect 10650 -795 10696 -757
rect 10650 -829 10656 -795
rect 10690 -829 10696 -795
rect 10650 -876 10696 -829
rect 10908 -723 10954 -574
rect 10908 -757 10914 -723
rect 10948 -757 10954 -723
rect 10908 -795 10954 -757
rect 10908 -829 10914 -795
rect 10948 -829 10954 -795
rect 10908 -876 10954 -829
rect 11166 -723 11212 -243
rect 11287 -344 11483 -336
rect 11287 -396 11294 -344
rect 11346 -396 11358 -344
rect 11410 -396 11422 -344
rect 11474 -396 11483 -344
rect 11287 -406 11483 -396
rect 11166 -757 11172 -723
rect 11206 -757 11212 -723
rect 11166 -795 11212 -757
rect 11166 -829 11172 -795
rect 11206 -829 11212 -795
rect 11166 -876 11212 -829
rect 11360 -723 11406 -406
rect 11360 -757 11366 -723
rect 11400 -757 11406 -723
rect 11360 -795 11406 -757
rect 11360 -829 11366 -795
rect 11400 -829 11406 -795
rect 11360 -876 11406 -829
rect 11618 -723 11664 -74
rect 11804 -344 12000 -336
rect 11804 -396 11811 -344
rect 11863 -396 11875 -344
rect 11927 -396 11939 -344
rect 11991 -396 12000 -344
rect 11804 -406 12000 -396
rect 11618 -757 11624 -723
rect 11658 -757 11664 -723
rect 11618 -795 11664 -757
rect 11618 -829 11624 -795
rect 11658 -829 11664 -795
rect 11618 -876 11664 -829
rect 11876 -723 11922 -406
rect 11876 -757 11882 -723
rect 11916 -757 11922 -723
rect 11876 -795 11922 -757
rect 11876 -829 11882 -795
rect 11916 -829 11922 -795
rect 11876 -876 11922 -829
rect 12134 -723 12180 -74
rect 13554 -88 13932 -54
rect 13966 -88 14344 -54
rect 15640 -12 15836 -4
rect 15640 -64 15649 -12
rect 15701 -64 15713 -12
rect 15765 -64 15777 -12
rect 15829 -64 15836 -12
rect 15640 -74 15836 -64
rect 16157 -12 16353 -4
rect 16157 -64 16166 -12
rect 16218 -64 16230 -12
rect 16282 -64 16294 -12
rect 16346 -64 16353 -12
rect 16157 -74 16353 -64
rect 17911 -16 18290 18
rect 18324 -16 18347 18
rect 17911 -54 18347 -16
rect 13554 -126 14344 -88
rect 13554 -160 13932 -126
rect 13966 -160 14344 -126
rect 12251 -181 12447 -173
rect 12251 -233 12260 -181
rect 12312 -233 12324 -181
rect 12376 -233 12388 -181
rect 12440 -233 12447 -181
rect 12251 -243 12447 -233
rect 12768 -181 12964 -173
rect 12768 -233 12777 -181
rect 12829 -233 12841 -181
rect 12893 -233 12905 -181
rect 12957 -233 12964 -181
rect 12768 -243 12964 -233
rect 13283 -181 13479 -173
rect 13283 -233 13292 -181
rect 13344 -233 13356 -181
rect 13408 -233 13420 -181
rect 13472 -233 13479 -181
rect 13283 -243 13479 -233
rect 13554 -198 14344 -160
rect 13554 -232 13932 -198
rect 13966 -232 14344 -198
rect 12134 -757 12140 -723
rect 12174 -757 12180 -723
rect 12134 -795 12180 -757
rect 12134 -829 12140 -795
rect 12174 -829 12180 -795
rect 12134 -876 12180 -829
rect 12328 -723 12374 -243
rect 12510 -512 12706 -504
rect 12510 -564 12519 -512
rect 12571 -564 12583 -512
rect 12635 -564 12647 -512
rect 12699 -564 12706 -512
rect 12510 -574 12706 -564
rect 12328 -757 12334 -723
rect 12368 -757 12374 -723
rect 12328 -795 12374 -757
rect 12328 -829 12334 -795
rect 12368 -829 12374 -795
rect 12328 -876 12374 -829
rect 12586 -723 12632 -574
rect 12586 -757 12592 -723
rect 12626 -757 12632 -723
rect 12586 -795 12632 -757
rect 12586 -829 12592 -795
rect 12626 -829 12632 -795
rect 12586 -876 12632 -829
rect 12844 -723 12890 -243
rect 13027 -512 13223 -504
rect 13027 -564 13036 -512
rect 13088 -564 13100 -512
rect 13152 -564 13164 -512
rect 13216 -564 13223 -512
rect 13027 -574 13223 -564
rect 12844 -757 12850 -723
rect 12884 -757 12890 -723
rect 12844 -795 12890 -757
rect 12844 -829 12850 -795
rect 12884 -829 12890 -795
rect 12844 -876 12890 -829
rect 13102 -723 13148 -574
rect 13102 -757 13108 -723
rect 13142 -757 13148 -723
rect 13102 -795 13148 -757
rect 13102 -829 13108 -795
rect 13142 -829 13148 -795
rect 13102 -876 13148 -829
rect 13360 -723 13406 -243
rect 13360 -757 13366 -723
rect 13400 -757 13406 -723
rect 13360 -795 13406 -757
rect 13360 -829 13366 -795
rect 13400 -829 13406 -795
rect 13360 -876 13406 -829
rect 13554 -270 14344 -232
rect 14418 -181 14614 -173
rect 14418 -233 14425 -181
rect 14477 -233 14489 -181
rect 14541 -233 14553 -181
rect 14605 -233 14614 -181
rect 14418 -243 14614 -233
rect 14933 -181 15129 -173
rect 14933 -233 14940 -181
rect 14992 -233 15004 -181
rect 15056 -233 15068 -181
rect 15120 -233 15129 -181
rect 14933 -243 15129 -233
rect 15450 -181 15646 -173
rect 15450 -233 15457 -181
rect 15509 -233 15521 -181
rect 15573 -233 15585 -181
rect 15637 -233 15646 -181
rect 15450 -243 15646 -233
rect 13554 -304 13932 -270
rect 13966 -304 14344 -270
rect 13554 -342 14344 -304
rect 13554 -376 13932 -342
rect 13966 -376 14344 -342
rect 13554 -414 14344 -376
rect 13554 -448 13932 -414
rect 13966 -448 14344 -414
rect 13554 -486 14344 -448
rect 13554 -520 13932 -486
rect 13966 -520 14344 -486
rect 13554 -558 14344 -520
rect 13554 -592 13932 -558
rect 13966 -592 14344 -558
rect 13554 -630 14344 -592
rect 13554 -664 13932 -630
rect 13966 -664 14344 -630
rect 13554 -702 14344 -664
rect 13554 -723 13932 -702
rect 13554 -757 13560 -723
rect 13594 -757 13818 -723
rect 13852 -736 13932 -723
rect 13966 -723 14344 -702
rect 13966 -736 14046 -723
rect 13852 -757 14046 -736
rect 14080 -757 14304 -723
rect 14338 -757 14344 -723
rect 13554 -774 14344 -757
rect 13554 -795 13932 -774
rect 13554 -829 13560 -795
rect 13594 -829 13818 -795
rect 13852 -808 13932 -795
rect 13966 -795 14344 -774
rect 13966 -808 14046 -795
rect 13852 -829 14046 -808
rect 14080 -829 14304 -795
rect 14338 -829 14344 -795
rect 13554 -846 14344 -829
rect 4836 -923 5214 -918
rect 4836 -957 4935 -923
rect 4969 -957 5007 -923
rect 5041 -952 5214 -923
rect 5248 -923 5626 -918
rect 5248 -952 5421 -923
rect 5041 -957 5421 -952
rect 5455 -957 5493 -923
rect 5527 -957 5626 -923
rect 4836 -990 5626 -957
rect 3529 -1238 3590 -1006
rect 4836 -1024 5214 -990
rect 5248 -1024 5626 -990
rect 5830 -923 6934 -917
rect 5830 -957 5873 -923
rect 5907 -936 5945 -923
rect 5979 -936 6131 -923
rect 6165 -936 6203 -923
rect 6237 -936 6389 -923
rect 6423 -936 6461 -923
rect 6495 -936 6647 -923
rect 6681 -936 6719 -923
rect 5830 -988 5880 -957
rect 5932 -988 5944 -936
rect 5996 -988 6008 -936
rect 6060 -988 6076 -936
rect 6128 -957 6131 -936
rect 6192 -957 6203 -936
rect 6128 -988 6140 -957
rect 6192 -988 6204 -957
rect 6256 -988 6366 -936
rect 6423 -957 6430 -936
rect 6418 -988 6430 -957
rect 6482 -988 6494 -957
rect 6546 -988 6562 -936
rect 6614 -988 6626 -936
rect 6681 -957 6690 -936
rect 6753 -957 6934 -923
rect 6678 -988 6690 -957
rect 6742 -988 6934 -957
rect 5830 -1006 6934 -988
rect 2516 -1286 3590 -1238
rect 2516 -1320 2742 -1286
rect 2776 -1320 2814 -1286
rect 2848 -1320 3000 -1286
rect 3034 -1320 3072 -1286
rect 3106 -1320 3258 -1286
rect 3292 -1320 3330 -1286
rect 3364 -1320 3590 -1286
rect 2516 -1326 3590 -1320
rect 3667 -1074 4633 -1056
rect 3667 -1126 3721 -1074
rect 3773 -1126 3785 -1074
rect 3837 -1126 3849 -1074
rect 3901 -1126 3917 -1074
rect 3969 -1126 3981 -1074
rect 4033 -1126 4045 -1074
rect 4097 -1126 4207 -1074
rect 4259 -1126 4271 -1074
rect 4323 -1126 4335 -1074
rect 4387 -1126 4403 -1074
rect 4455 -1126 4467 -1074
rect 4519 -1126 4531 -1074
rect 4583 -1126 4633 -1074
rect 3667 -1252 4633 -1126
rect 3667 -1286 3721 -1252
rect 3773 -1286 3785 -1252
rect 3667 -1320 3710 -1286
rect 3773 -1304 3782 -1286
rect 3837 -1304 3849 -1252
rect 3901 -1304 3917 -1252
rect 3969 -1286 3981 -1252
rect 4033 -1286 4045 -1252
rect 4033 -1304 4040 -1286
rect 4097 -1304 4207 -1252
rect 4259 -1286 4271 -1252
rect 4323 -1286 4335 -1252
rect 4260 -1304 4271 -1286
rect 4332 -1304 4335 -1286
rect 4387 -1304 4403 -1252
rect 4455 -1304 4467 -1252
rect 4519 -1304 4531 -1252
rect 4583 -1286 4633 -1252
rect 3744 -1320 3782 -1304
rect 3816 -1320 3968 -1304
rect 4002 -1320 4040 -1304
rect 4074 -1320 4226 -1304
rect 4260 -1320 4298 -1304
rect 4332 -1320 4484 -1304
rect 4518 -1320 4556 -1304
rect 4590 -1320 4633 -1286
rect 3667 -1326 4633 -1320
rect 4836 -1062 5626 -1024
rect 4836 -1096 5214 -1062
rect 5248 -1096 5626 -1062
rect 4836 -1134 5626 -1096
rect 4836 -1168 5214 -1134
rect 5248 -1168 5626 -1134
rect 4836 -1206 5626 -1168
rect 4836 -1240 5214 -1206
rect 5248 -1240 5626 -1206
rect 4836 -1278 5626 -1240
rect 4836 -1286 5214 -1278
rect 4836 -1320 4935 -1286
rect 4969 -1320 5007 -1286
rect 5041 -1312 5214 -1286
rect 5248 -1286 5626 -1278
rect 5248 -1312 5421 -1286
rect 5041 -1320 5421 -1312
rect 5455 -1320 5493 -1286
rect 5527 -1320 5626 -1286
rect 833 -1384 856 -1350
rect 890 -1384 1269 -1350
rect 4836 -1350 5626 -1320
rect 5830 -1074 6796 -1056
rect 5830 -1126 5880 -1074
rect 5932 -1126 5944 -1074
rect 5996 -1126 6008 -1074
rect 6060 -1126 6076 -1074
rect 6128 -1126 6140 -1074
rect 6192 -1126 6204 -1074
rect 6256 -1126 6366 -1074
rect 6418 -1126 6430 -1074
rect 6482 -1126 6494 -1074
rect 6546 -1126 6562 -1074
rect 6614 -1126 6626 -1074
rect 6678 -1126 6690 -1074
rect 6742 -1126 6796 -1074
rect 5830 -1252 6796 -1126
rect 5830 -1286 5880 -1252
rect 5830 -1320 5873 -1286
rect 5932 -1304 5944 -1252
rect 5996 -1304 6008 -1252
rect 6060 -1304 6076 -1252
rect 6128 -1286 6140 -1252
rect 6192 -1286 6204 -1252
rect 6128 -1304 6131 -1286
rect 6192 -1304 6203 -1286
rect 6256 -1304 6366 -1252
rect 6418 -1286 6430 -1252
rect 6482 -1286 6494 -1252
rect 6423 -1304 6430 -1286
rect 6546 -1304 6562 -1252
rect 6614 -1304 6626 -1252
rect 6678 -1286 6690 -1252
rect 6742 -1286 6796 -1252
rect 6681 -1304 6690 -1286
rect 5907 -1320 5945 -1304
rect 5979 -1320 6131 -1304
rect 6165 -1320 6203 -1304
rect 6237 -1320 6389 -1304
rect 6423 -1320 6461 -1304
rect 6495 -1320 6647 -1304
rect 6681 -1320 6719 -1304
rect 6753 -1320 6796 -1286
rect 5830 -1326 6796 -1320
rect 6873 -1238 6934 -1006
rect 7056 -923 7764 -917
rect 7056 -957 7099 -923
rect 7133 -957 7171 -923
rect 7205 -957 7357 -923
rect 7391 -957 7429 -923
rect 7463 -957 7615 -923
rect 7649 -957 7687 -923
rect 7721 -957 7764 -923
rect 7056 -1074 7764 -957
rect 7056 -1126 7094 -1074
rect 7146 -1126 7158 -1074
rect 7210 -1126 7222 -1074
rect 7274 -1126 7290 -1074
rect 7342 -1126 7354 -1074
rect 7406 -1126 7418 -1074
rect 7470 -1126 7482 -1074
rect 7534 -1126 7550 -1074
rect 7602 -1126 7614 -1074
rect 7666 -1126 7678 -1074
rect 7730 -1126 7764 -1074
rect 7056 -1144 7764 -1126
rect 7886 -923 8990 -917
rect 7886 -957 8067 -923
rect 8101 -936 8139 -923
rect 8173 -936 8325 -923
rect 8359 -936 8397 -923
rect 8431 -936 8583 -923
rect 8617 -936 8655 -923
rect 8689 -936 8841 -923
rect 8875 -936 8913 -923
rect 8130 -957 8139 -936
rect 7886 -988 8078 -957
rect 8130 -988 8142 -957
rect 8194 -988 8206 -936
rect 8258 -988 8274 -936
rect 8390 -957 8397 -936
rect 8326 -988 8338 -957
rect 8390 -988 8402 -957
rect 8454 -988 8564 -936
rect 8617 -957 8628 -936
rect 8689 -957 8692 -936
rect 8616 -988 8628 -957
rect 8680 -988 8692 -957
rect 8744 -988 8760 -936
rect 8812 -988 8824 -936
rect 8876 -988 8888 -936
rect 8947 -957 8990 -923
rect 8940 -988 8990 -957
rect 7886 -1006 8990 -988
rect 9194 -918 9986 -880
rect 13554 -880 13932 -846
rect 13966 -880 14344 -846
rect 14491 -723 14537 -243
rect 14674 -512 14870 -504
rect 14674 -564 14681 -512
rect 14733 -564 14745 -512
rect 14797 -564 14809 -512
rect 14861 -564 14870 -512
rect 14674 -574 14870 -564
rect 14491 -757 14497 -723
rect 14531 -757 14537 -723
rect 14491 -795 14537 -757
rect 14491 -829 14497 -795
rect 14531 -829 14537 -795
rect 14491 -876 14537 -829
rect 14749 -723 14795 -574
rect 14749 -757 14755 -723
rect 14789 -757 14795 -723
rect 14749 -795 14795 -757
rect 14749 -829 14755 -795
rect 14789 -829 14795 -795
rect 14749 -876 14795 -829
rect 15007 -723 15053 -243
rect 15191 -512 15387 -504
rect 15191 -564 15198 -512
rect 15250 -564 15262 -512
rect 15314 -564 15326 -512
rect 15378 -564 15387 -512
rect 15191 -574 15387 -564
rect 15007 -757 15013 -723
rect 15047 -757 15053 -723
rect 15007 -795 15053 -757
rect 15007 -829 15013 -795
rect 15047 -829 15053 -795
rect 15007 -876 15053 -829
rect 15265 -723 15311 -574
rect 15265 -757 15271 -723
rect 15305 -757 15311 -723
rect 15265 -795 15311 -757
rect 15265 -829 15271 -795
rect 15305 -829 15311 -795
rect 15265 -876 15311 -829
rect 15523 -723 15569 -243
rect 15523 -757 15529 -723
rect 15563 -757 15569 -723
rect 15523 -795 15569 -757
rect 15523 -829 15529 -795
rect 15563 -829 15569 -795
rect 15523 -876 15569 -829
rect 15717 -723 15763 -74
rect 15897 -344 16093 -336
rect 15897 -396 15906 -344
rect 15958 -396 15970 -344
rect 16022 -396 16034 -344
rect 16086 -396 16093 -344
rect 15897 -406 16093 -396
rect 15717 -757 15723 -723
rect 15757 -757 15763 -723
rect 15717 -795 15763 -757
rect 15717 -829 15723 -795
rect 15757 -829 15763 -795
rect 15717 -876 15763 -829
rect 15975 -723 16021 -406
rect 15975 -757 15981 -723
rect 16015 -757 16021 -723
rect 15975 -795 16021 -757
rect 15975 -829 15981 -795
rect 16015 -829 16021 -795
rect 15975 -876 16021 -829
rect 16233 -723 16279 -74
rect 17911 -88 18290 -54
rect 18324 -88 18347 -54
rect 17911 -126 18347 -88
rect 17911 -160 18290 -126
rect 18324 -160 18347 -126
rect 16611 -181 16807 -173
rect 16611 -233 16618 -181
rect 16670 -233 16682 -181
rect 16734 -233 16746 -181
rect 16798 -233 16807 -181
rect 16611 -243 16807 -233
rect 17128 -181 17324 -173
rect 17128 -233 17135 -181
rect 17187 -233 17199 -181
rect 17251 -233 17263 -181
rect 17315 -233 17324 -181
rect 17128 -243 17324 -233
rect 17645 -181 17841 -173
rect 17645 -233 17652 -181
rect 17704 -233 17716 -181
rect 17768 -233 17780 -181
rect 17832 -233 17841 -181
rect 17645 -243 17841 -233
rect 17911 -198 18347 -160
rect 17911 -232 18290 -198
rect 18324 -232 18347 -198
rect 16414 -344 16610 -336
rect 16414 -396 16423 -344
rect 16475 -396 16487 -344
rect 16539 -396 16551 -344
rect 16603 -396 16610 -344
rect 16414 -406 16610 -396
rect 16233 -757 16239 -723
rect 16273 -757 16279 -723
rect 16233 -795 16279 -757
rect 16233 -829 16239 -795
rect 16273 -829 16279 -795
rect 16233 -876 16279 -829
rect 16491 -723 16537 -406
rect 16491 -757 16497 -723
rect 16531 -757 16537 -723
rect 16491 -795 16537 -757
rect 16491 -829 16497 -795
rect 16531 -829 16537 -795
rect 16491 -876 16537 -829
rect 16685 -723 16731 -243
rect 16868 -512 17064 -504
rect 16868 -564 16875 -512
rect 16927 -564 16939 -512
rect 16991 -564 17003 -512
rect 17055 -564 17064 -512
rect 16868 -574 17064 -564
rect 16685 -757 16691 -723
rect 16725 -757 16731 -723
rect 16685 -795 16731 -757
rect 16685 -829 16691 -795
rect 16725 -829 16731 -795
rect 16685 -876 16731 -829
rect 16943 -723 16989 -574
rect 16943 -757 16949 -723
rect 16983 -757 16989 -723
rect 16943 -795 16989 -757
rect 16943 -829 16949 -795
rect 16983 -829 16989 -795
rect 16943 -876 16989 -829
rect 17201 -723 17247 -243
rect 17386 -512 17582 -504
rect 17386 -564 17393 -512
rect 17445 -564 17457 -512
rect 17509 -564 17521 -512
rect 17573 -564 17582 -512
rect 17386 -574 17582 -564
rect 17201 -757 17207 -723
rect 17241 -757 17247 -723
rect 17201 -795 17247 -757
rect 17201 -829 17207 -795
rect 17241 -829 17247 -795
rect 17201 -876 17247 -829
rect 17459 -723 17505 -574
rect 17459 -757 17465 -723
rect 17499 -757 17505 -723
rect 17459 -795 17505 -757
rect 17459 -829 17465 -795
rect 17499 -829 17505 -795
rect 17459 -876 17505 -829
rect 17717 -723 17763 -243
rect 17717 -757 17723 -723
rect 17757 -757 17763 -723
rect 17717 -795 17763 -757
rect 17717 -829 17723 -795
rect 17757 -829 17763 -795
rect 17717 -876 17763 -829
rect 17911 -270 18347 -232
rect 17911 -304 18290 -270
rect 18324 -304 18347 -270
rect 17911 -342 18347 -304
rect 17911 -376 18290 -342
rect 18324 -376 18347 -342
rect 17911 -414 18347 -376
rect 17911 -448 18290 -414
rect 18324 -448 18347 -414
rect 17911 -486 18347 -448
rect 17911 -520 18290 -486
rect 18324 -520 18347 -486
rect 17911 -558 18347 -520
rect 17911 -592 18290 -558
rect 18324 -592 18347 -558
rect 17911 -630 18347 -592
rect 17911 -664 18290 -630
rect 18324 -664 18347 -630
rect 17911 -702 18347 -664
rect 17911 -723 18290 -702
rect 17911 -757 17917 -723
rect 17951 -757 18175 -723
rect 18209 -736 18290 -723
rect 18324 -736 18347 -702
rect 18209 -757 18347 -736
rect 17911 -774 18347 -757
rect 17911 -795 18290 -774
rect 17911 -829 17917 -795
rect 17951 -829 18175 -795
rect 18209 -808 18290 -795
rect 18324 -808 18347 -774
rect 18209 -829 18347 -808
rect 17911 -846 18347 -829
rect 9194 -923 9573 -918
rect 9194 -957 9293 -923
rect 9327 -957 9365 -923
rect 9399 -952 9573 -923
rect 9607 -923 9986 -918
rect 9607 -952 9781 -923
rect 9399 -957 9781 -952
rect 9815 -957 9853 -923
rect 9887 -957 9986 -923
rect 9194 -990 9986 -957
rect 7886 -1238 7947 -1006
rect 9194 -1024 9573 -990
rect 9607 -1024 9986 -990
rect 10190 -923 11294 -917
rect 10190 -957 10233 -923
rect 10267 -936 10305 -923
rect 10339 -936 10491 -923
rect 10525 -936 10563 -923
rect 10597 -936 10749 -923
rect 10783 -936 10821 -923
rect 10855 -936 11007 -923
rect 11041 -936 11079 -923
rect 10190 -988 10240 -957
rect 10292 -988 10304 -936
rect 10356 -988 10368 -936
rect 10420 -988 10436 -936
rect 10488 -957 10491 -936
rect 10552 -957 10563 -936
rect 10488 -988 10500 -957
rect 10552 -988 10564 -957
rect 10616 -988 10726 -936
rect 10783 -957 10790 -936
rect 10778 -988 10790 -957
rect 10842 -988 10854 -957
rect 10906 -988 10922 -936
rect 10974 -988 10986 -936
rect 11041 -957 11050 -936
rect 11113 -957 11294 -923
rect 11038 -988 11050 -957
rect 11102 -988 11294 -957
rect 10190 -1006 11294 -988
rect 6873 -1286 7947 -1238
rect 6873 -1320 7099 -1286
rect 7133 -1320 7171 -1286
rect 7205 -1320 7357 -1286
rect 7391 -1320 7429 -1286
rect 7463 -1320 7615 -1286
rect 7649 -1320 7687 -1286
rect 7721 -1320 7947 -1286
rect 6873 -1326 7947 -1320
rect 8024 -1074 8990 -1056
rect 8024 -1126 8078 -1074
rect 8130 -1126 8142 -1074
rect 8194 -1126 8206 -1074
rect 8258 -1126 8274 -1074
rect 8326 -1126 8338 -1074
rect 8390 -1126 8402 -1074
rect 8454 -1126 8564 -1074
rect 8616 -1126 8628 -1074
rect 8680 -1126 8692 -1074
rect 8744 -1126 8760 -1074
rect 8812 -1126 8824 -1074
rect 8876 -1126 8888 -1074
rect 8940 -1126 8990 -1074
rect 8024 -1252 8990 -1126
rect 8024 -1286 8078 -1252
rect 8130 -1286 8142 -1252
rect 8024 -1320 8067 -1286
rect 8130 -1304 8139 -1286
rect 8194 -1304 8206 -1252
rect 8258 -1304 8274 -1252
rect 8326 -1286 8338 -1252
rect 8390 -1286 8402 -1252
rect 8390 -1304 8397 -1286
rect 8454 -1304 8564 -1252
rect 8616 -1286 8628 -1252
rect 8680 -1286 8692 -1252
rect 8617 -1304 8628 -1286
rect 8689 -1304 8692 -1286
rect 8744 -1304 8760 -1252
rect 8812 -1304 8824 -1252
rect 8876 -1304 8888 -1252
rect 8940 -1286 8990 -1252
rect 8101 -1320 8139 -1304
rect 8173 -1320 8325 -1304
rect 8359 -1320 8397 -1304
rect 8431 -1320 8583 -1304
rect 8617 -1320 8655 -1304
rect 8689 -1320 8841 -1304
rect 8875 -1320 8913 -1304
rect 8947 -1320 8990 -1286
rect 8024 -1326 8990 -1320
rect 9194 -1062 9986 -1024
rect 9194 -1096 9573 -1062
rect 9607 -1096 9986 -1062
rect 9194 -1134 9986 -1096
rect 9194 -1168 9573 -1134
rect 9607 -1168 9986 -1134
rect 9194 -1206 9986 -1168
rect 9194 -1240 9573 -1206
rect 9607 -1240 9986 -1206
rect 9194 -1278 9986 -1240
rect 9194 -1286 9573 -1278
rect 9194 -1320 9293 -1286
rect 9327 -1320 9365 -1286
rect 9399 -1312 9573 -1286
rect 9607 -1286 9986 -1278
rect 9607 -1312 9781 -1286
rect 9399 -1320 9781 -1312
rect 9815 -1320 9853 -1286
rect 9887 -1320 9986 -1286
rect 833 -1414 1269 -1384
rect 833 -1422 971 -1414
rect 833 -1456 856 -1422
rect 890 -1448 971 -1422
rect 1005 -1448 1229 -1414
rect 1263 -1448 1269 -1414
rect 890 -1456 1269 -1448
rect 833 -1486 1269 -1456
rect 833 -1494 971 -1486
rect 833 -1528 856 -1494
rect 890 -1520 971 -1494
rect 1005 -1520 1229 -1486
rect 1263 -1520 1269 -1486
rect 890 -1528 1269 -1520
rect 833 -1566 1269 -1528
rect 833 -1600 856 -1566
rect 890 -1600 1269 -1566
rect 833 -1638 1269 -1600
rect 833 -1672 856 -1638
rect 890 -1672 1269 -1638
rect 833 -1710 1269 -1672
rect 1417 -1414 1463 -1367
rect 1417 -1448 1423 -1414
rect 1457 -1448 1463 -1414
rect 1417 -1486 1463 -1448
rect 1417 -1520 1423 -1486
rect 1457 -1520 1463 -1486
rect 1417 -1694 1463 -1520
rect 1675 -1414 1721 -1367
rect 1675 -1448 1681 -1414
rect 1715 -1448 1721 -1414
rect 1675 -1486 1721 -1448
rect 1675 -1520 1681 -1486
rect 1715 -1520 1721 -1486
rect 833 -1744 856 -1710
rect 890 -1744 1269 -1710
rect 833 -1782 1269 -1744
rect 1343 -1702 1539 -1694
rect 1343 -1754 1350 -1702
rect 1402 -1754 1414 -1702
rect 1466 -1754 1478 -1702
rect 1530 -1754 1539 -1702
rect 1343 -1764 1539 -1754
rect 833 -1816 856 -1782
rect 890 -1816 1269 -1782
rect 833 -1854 1269 -1816
rect 833 -1888 856 -1854
rect 890 -1888 1269 -1854
rect 833 -1926 1269 -1888
rect 833 -1960 856 -1926
rect 890 -1960 1269 -1926
rect 833 -1998 1269 -1960
rect 833 -2032 856 -1998
rect 890 -2032 1269 -1998
rect 833 -2070 1269 -2032
rect 833 -2104 856 -2070
rect 890 -2104 1269 -2070
rect 833 -2142 1269 -2104
rect 833 -2176 856 -2142
rect 890 -2176 1269 -2142
rect 833 -2214 1269 -2176
rect 833 -2248 856 -2214
rect 890 -2248 1269 -2214
rect 833 -2286 1269 -2248
rect 833 -2320 856 -2286
rect 890 -2320 1269 -2286
rect 833 -2358 1269 -2320
rect 833 -2392 856 -2358
rect 890 -2370 1269 -2358
rect 890 -2392 971 -2370
rect 833 -2404 971 -2392
rect 1005 -2404 1229 -2370
rect 1263 -2404 1269 -2370
rect 833 -2430 1269 -2404
rect 833 -2464 856 -2430
rect 890 -2442 1269 -2430
rect 890 -2464 971 -2442
rect 833 -2476 971 -2464
rect 1005 -2476 1229 -2442
rect 1263 -2476 1269 -2442
rect 833 -2502 1269 -2476
rect 833 -2536 856 -2502
rect 890 -2536 1269 -2502
rect 1417 -2370 1463 -1764
rect 1675 -1995 1721 -1520
rect 1933 -1414 1979 -1367
rect 1933 -1448 1939 -1414
rect 1973 -1448 1979 -1414
rect 1933 -1486 1979 -1448
rect 1933 -1520 1939 -1486
rect 1973 -1520 1979 -1486
rect 1933 -1694 1979 -1520
rect 2191 -1414 2237 -1367
rect 2191 -1448 2197 -1414
rect 2231 -1448 2237 -1414
rect 2191 -1486 2237 -1448
rect 2191 -1520 2197 -1486
rect 2231 -1520 2237 -1486
rect 1858 -1702 2054 -1694
rect 1858 -1754 1865 -1702
rect 1917 -1754 1929 -1702
rect 1981 -1754 1993 -1702
rect 2045 -1754 2054 -1702
rect 1858 -1764 2054 -1754
rect 1601 -2003 1797 -1995
rect 1601 -2055 1608 -2003
rect 1660 -2055 1672 -2003
rect 1724 -2055 1736 -2003
rect 1788 -2055 1797 -2003
rect 1601 -2065 1797 -2055
rect 1417 -2404 1423 -2370
rect 1457 -2404 1463 -2370
rect 1417 -2442 1463 -2404
rect 1417 -2476 1423 -2442
rect 1457 -2476 1463 -2442
rect 1417 -2523 1463 -2476
rect 1675 -2370 1721 -2065
rect 1675 -2404 1681 -2370
rect 1715 -2404 1721 -2370
rect 1675 -2442 1721 -2404
rect 1675 -2476 1681 -2442
rect 1715 -2476 1721 -2442
rect 1675 -2523 1721 -2476
rect 1933 -2370 1979 -1764
rect 2191 -1995 2237 -1520
rect 2449 -1414 2495 -1367
rect 2449 -1448 2455 -1414
rect 2489 -1448 2495 -1414
rect 2449 -1486 2495 -1448
rect 2449 -1520 2455 -1486
rect 2489 -1520 2495 -1486
rect 2449 -1694 2495 -1520
rect 2643 -1414 2689 -1367
rect 2643 -1448 2649 -1414
rect 2683 -1448 2689 -1414
rect 2643 -1486 2689 -1448
rect 2643 -1520 2649 -1486
rect 2683 -1520 2689 -1486
rect 2376 -1702 2572 -1694
rect 2376 -1754 2383 -1702
rect 2435 -1754 2447 -1702
rect 2499 -1754 2511 -1702
rect 2563 -1754 2572 -1702
rect 2376 -1764 2572 -1754
rect 2119 -2003 2315 -1995
rect 2119 -2055 2126 -2003
rect 2178 -2055 2190 -2003
rect 2242 -2055 2254 -2003
rect 2306 -2055 2315 -2003
rect 2119 -2065 2315 -2055
rect 1933 -2404 1939 -2370
rect 1973 -2404 1979 -2370
rect 1933 -2442 1979 -2404
rect 1933 -2476 1939 -2442
rect 1973 -2476 1979 -2442
rect 1933 -2523 1979 -2476
rect 2191 -2370 2237 -2065
rect 2191 -2404 2197 -2370
rect 2231 -2404 2237 -2370
rect 2191 -2442 2237 -2404
rect 2191 -2476 2197 -2442
rect 2231 -2476 2237 -2442
rect 2191 -2523 2237 -2476
rect 2449 -2370 2495 -1764
rect 2643 -2139 2689 -1520
rect 2901 -1414 2947 -1367
rect 2901 -1448 2907 -1414
rect 2941 -1448 2947 -1414
rect 2901 -1486 2947 -1448
rect 2901 -1520 2907 -1486
rect 2941 -1520 2947 -1486
rect 2901 -1834 2947 -1520
rect 3159 -1414 3205 -1367
rect 3159 -1448 3165 -1414
rect 3199 -1448 3205 -1414
rect 3159 -1486 3205 -1448
rect 3159 -1520 3165 -1486
rect 3199 -1520 3205 -1486
rect 2824 -1842 3020 -1834
rect 2824 -1894 2833 -1842
rect 2885 -1894 2897 -1842
rect 2949 -1894 2961 -1842
rect 3013 -1894 3020 -1842
rect 2824 -1904 3020 -1894
rect 2566 -2147 2762 -2139
rect 2566 -2199 2575 -2147
rect 2627 -2199 2639 -2147
rect 2691 -2199 2703 -2147
rect 2755 -2199 2762 -2147
rect 2566 -2209 2762 -2199
rect 2449 -2404 2455 -2370
rect 2489 -2404 2495 -2370
rect 2449 -2442 2495 -2404
rect 2449 -2476 2455 -2442
rect 2489 -2476 2495 -2442
rect 2449 -2523 2495 -2476
rect 2643 -2370 2689 -2209
rect 2643 -2404 2649 -2370
rect 2683 -2404 2689 -2370
rect 2643 -2442 2689 -2404
rect 2643 -2476 2649 -2442
rect 2683 -2476 2689 -2442
rect 2643 -2523 2689 -2476
rect 2901 -2370 2947 -1904
rect 3159 -2139 3205 -1520
rect 3417 -1414 3463 -1367
rect 3417 -1448 3423 -1414
rect 3457 -1448 3463 -1414
rect 3417 -1486 3463 -1448
rect 3417 -1520 3423 -1486
rect 3457 -1520 3463 -1486
rect 3417 -1834 3463 -1520
rect 3611 -1414 3657 -1367
rect 3611 -1448 3617 -1414
rect 3651 -1448 3657 -1414
rect 3611 -1486 3657 -1448
rect 3611 -1520 3617 -1486
rect 3651 -1520 3657 -1486
rect 3611 -1694 3657 -1520
rect 3869 -1414 3915 -1367
rect 3869 -1448 3875 -1414
rect 3909 -1448 3915 -1414
rect 3869 -1486 3915 -1448
rect 3869 -1520 3875 -1486
rect 3909 -1520 3915 -1486
rect 3536 -1702 3732 -1694
rect 3536 -1754 3543 -1702
rect 3595 -1754 3607 -1702
rect 3659 -1754 3671 -1702
rect 3723 -1754 3732 -1702
rect 3536 -1764 3732 -1754
rect 3341 -1842 3537 -1834
rect 3341 -1894 3350 -1842
rect 3402 -1894 3414 -1842
rect 3466 -1894 3478 -1842
rect 3530 -1894 3537 -1842
rect 3341 -1904 3537 -1894
rect 3083 -2147 3279 -2139
rect 3083 -2199 3092 -2147
rect 3144 -2199 3156 -2147
rect 3208 -2199 3220 -2147
rect 3272 -2199 3279 -2147
rect 3083 -2209 3279 -2199
rect 2901 -2404 2907 -2370
rect 2941 -2404 2947 -2370
rect 2901 -2442 2947 -2404
rect 2901 -2476 2907 -2442
rect 2941 -2476 2947 -2442
rect 2901 -2523 2947 -2476
rect 3159 -2370 3205 -2209
rect 3159 -2404 3165 -2370
rect 3199 -2404 3205 -2370
rect 3159 -2442 3205 -2404
rect 3159 -2476 3165 -2442
rect 3199 -2476 3205 -2442
rect 3159 -2523 3205 -2476
rect 3417 -2370 3463 -1904
rect 3417 -2404 3423 -2370
rect 3457 -2404 3463 -2370
rect 3417 -2442 3463 -2404
rect 3417 -2476 3423 -2442
rect 3457 -2476 3463 -2442
rect 3417 -2523 3463 -2476
rect 3611 -2370 3657 -1764
rect 3869 -1995 3915 -1520
rect 4127 -1414 4173 -1367
rect 4127 -1448 4133 -1414
rect 4167 -1448 4173 -1414
rect 4127 -1486 4173 -1448
rect 4127 -1520 4133 -1486
rect 4167 -1520 4173 -1486
rect 4127 -1694 4173 -1520
rect 4385 -1414 4431 -1367
rect 4385 -1448 4391 -1414
rect 4425 -1448 4431 -1414
rect 4385 -1486 4431 -1448
rect 4385 -1520 4391 -1486
rect 4425 -1520 4431 -1486
rect 4053 -1702 4249 -1694
rect 4053 -1754 4060 -1702
rect 4112 -1754 4124 -1702
rect 4176 -1754 4188 -1702
rect 4240 -1754 4249 -1702
rect 4053 -1764 4249 -1754
rect 3796 -2003 3992 -1995
rect 3796 -2055 3803 -2003
rect 3855 -2055 3867 -2003
rect 3919 -2055 3931 -2003
rect 3983 -2055 3992 -2003
rect 3796 -2065 3992 -2055
rect 3611 -2404 3617 -2370
rect 3651 -2404 3657 -2370
rect 3611 -2442 3657 -2404
rect 3611 -2476 3617 -2442
rect 3651 -2476 3657 -2442
rect 3611 -2523 3657 -2476
rect 3869 -2370 3915 -2065
rect 3869 -2404 3875 -2370
rect 3909 -2404 3915 -2370
rect 3869 -2442 3915 -2404
rect 3869 -2476 3875 -2442
rect 3909 -2476 3915 -2442
rect 3869 -2523 3915 -2476
rect 4127 -2370 4173 -1764
rect 4385 -1995 4431 -1520
rect 4643 -1414 4689 -1367
rect 4643 -1448 4649 -1414
rect 4683 -1448 4689 -1414
rect 4643 -1486 4689 -1448
rect 4643 -1520 4649 -1486
rect 4683 -1520 4689 -1486
rect 4643 -1694 4689 -1520
rect 4836 -1384 5214 -1350
rect 5248 -1384 5626 -1350
rect 9194 -1350 9986 -1320
rect 10190 -1074 11156 -1056
rect 10190 -1126 10240 -1074
rect 10292 -1126 10304 -1074
rect 10356 -1126 10368 -1074
rect 10420 -1126 10436 -1074
rect 10488 -1126 10500 -1074
rect 10552 -1126 10564 -1074
rect 10616 -1126 10726 -1074
rect 10778 -1126 10790 -1074
rect 10842 -1126 10854 -1074
rect 10906 -1126 10922 -1074
rect 10974 -1126 10986 -1074
rect 11038 -1126 11050 -1074
rect 11102 -1126 11156 -1074
rect 10190 -1252 11156 -1126
rect 10190 -1286 10240 -1252
rect 10190 -1320 10233 -1286
rect 10292 -1304 10304 -1252
rect 10356 -1304 10368 -1252
rect 10420 -1304 10436 -1252
rect 10488 -1286 10500 -1252
rect 10552 -1286 10564 -1252
rect 10488 -1304 10491 -1286
rect 10552 -1304 10563 -1286
rect 10616 -1304 10726 -1252
rect 10778 -1286 10790 -1252
rect 10842 -1286 10854 -1252
rect 10783 -1304 10790 -1286
rect 10906 -1304 10922 -1252
rect 10974 -1304 10986 -1252
rect 11038 -1286 11050 -1252
rect 11102 -1286 11156 -1252
rect 11041 -1304 11050 -1286
rect 10267 -1320 10305 -1304
rect 10339 -1320 10491 -1304
rect 10525 -1320 10563 -1304
rect 10597 -1320 10749 -1304
rect 10783 -1320 10821 -1304
rect 10855 -1320 11007 -1304
rect 11041 -1320 11079 -1304
rect 11113 -1320 11156 -1286
rect 10190 -1326 11156 -1320
rect 11233 -1238 11294 -1006
rect 11416 -923 12124 -917
rect 11416 -957 11459 -923
rect 11493 -957 11531 -923
rect 11565 -957 11717 -923
rect 11751 -957 11789 -923
rect 11823 -957 11975 -923
rect 12009 -957 12047 -923
rect 12081 -957 12124 -923
rect 11416 -1074 12124 -957
rect 11416 -1126 11450 -1074
rect 11502 -1126 11514 -1074
rect 11566 -1126 11578 -1074
rect 11630 -1126 11646 -1074
rect 11698 -1126 11710 -1074
rect 11762 -1126 11774 -1074
rect 11826 -1126 11838 -1074
rect 11890 -1126 11906 -1074
rect 11958 -1126 11970 -1074
rect 12022 -1126 12034 -1074
rect 12086 -1126 12124 -1074
rect 11416 -1144 12124 -1126
rect 12246 -923 13350 -917
rect 12246 -957 12427 -923
rect 12461 -936 12499 -923
rect 12533 -936 12685 -923
rect 12719 -936 12757 -923
rect 12791 -936 12943 -923
rect 12977 -936 13015 -923
rect 13049 -936 13201 -923
rect 13235 -936 13273 -923
rect 12490 -957 12499 -936
rect 12246 -988 12438 -957
rect 12490 -988 12502 -957
rect 12554 -988 12566 -936
rect 12618 -988 12634 -936
rect 12750 -957 12757 -936
rect 12686 -988 12698 -957
rect 12750 -988 12762 -957
rect 12814 -988 12924 -936
rect 12977 -957 12988 -936
rect 13049 -957 13052 -936
rect 12976 -988 12988 -957
rect 13040 -988 13052 -957
rect 13104 -988 13120 -936
rect 13172 -988 13184 -936
rect 13236 -988 13248 -936
rect 13307 -957 13350 -923
rect 13300 -988 13350 -957
rect 12246 -1006 13350 -988
rect 13554 -918 14344 -880
rect 17911 -880 18290 -846
rect 18324 -880 18347 -846
rect 13554 -923 13932 -918
rect 13554 -957 13653 -923
rect 13687 -957 13725 -923
rect 13759 -952 13932 -923
rect 13966 -923 14344 -918
rect 13966 -952 14139 -923
rect 13759 -957 14139 -952
rect 14173 -957 14211 -923
rect 14245 -957 14344 -923
rect 13554 -990 14344 -957
rect 12246 -1238 12307 -1006
rect 13554 -1024 13932 -990
rect 13966 -1024 14344 -990
rect 14547 -923 15651 -917
rect 14547 -957 14590 -923
rect 14624 -936 14662 -923
rect 14696 -936 14848 -923
rect 14882 -936 14920 -923
rect 14954 -936 15106 -923
rect 15140 -936 15178 -923
rect 15212 -936 15364 -923
rect 15398 -936 15436 -923
rect 14547 -988 14597 -957
rect 14649 -988 14661 -936
rect 14713 -988 14725 -936
rect 14777 -988 14793 -936
rect 14845 -957 14848 -936
rect 14909 -957 14920 -936
rect 14845 -988 14857 -957
rect 14909 -988 14921 -957
rect 14973 -988 15083 -936
rect 15140 -957 15147 -936
rect 15135 -988 15147 -957
rect 15199 -988 15211 -957
rect 15263 -988 15279 -936
rect 15331 -988 15343 -936
rect 15398 -957 15407 -936
rect 15470 -957 15651 -923
rect 15395 -988 15407 -957
rect 15459 -988 15651 -957
rect 14547 -1006 15651 -988
rect 11233 -1286 12307 -1238
rect 11233 -1320 11459 -1286
rect 11493 -1320 11531 -1286
rect 11565 -1320 11717 -1286
rect 11751 -1320 11789 -1286
rect 11823 -1320 11975 -1286
rect 12009 -1320 12047 -1286
rect 12081 -1320 12307 -1286
rect 11233 -1326 12307 -1320
rect 12384 -1074 13350 -1056
rect 12384 -1126 12438 -1074
rect 12490 -1126 12502 -1074
rect 12554 -1126 12566 -1074
rect 12618 -1126 12634 -1074
rect 12686 -1126 12698 -1074
rect 12750 -1126 12762 -1074
rect 12814 -1126 12924 -1074
rect 12976 -1126 12988 -1074
rect 13040 -1126 13052 -1074
rect 13104 -1126 13120 -1074
rect 13172 -1126 13184 -1074
rect 13236 -1126 13248 -1074
rect 13300 -1126 13350 -1074
rect 12384 -1252 13350 -1126
rect 12384 -1286 12438 -1252
rect 12490 -1286 12502 -1252
rect 12384 -1320 12427 -1286
rect 12490 -1304 12499 -1286
rect 12554 -1304 12566 -1252
rect 12618 -1304 12634 -1252
rect 12686 -1286 12698 -1252
rect 12750 -1286 12762 -1252
rect 12750 -1304 12757 -1286
rect 12814 -1304 12924 -1252
rect 12976 -1286 12988 -1252
rect 13040 -1286 13052 -1252
rect 12977 -1304 12988 -1286
rect 13049 -1304 13052 -1286
rect 13104 -1304 13120 -1252
rect 13172 -1304 13184 -1252
rect 13236 -1304 13248 -1252
rect 13300 -1286 13350 -1252
rect 12461 -1320 12499 -1304
rect 12533 -1320 12685 -1304
rect 12719 -1320 12757 -1304
rect 12791 -1320 12943 -1304
rect 12977 -1320 13015 -1304
rect 13049 -1320 13201 -1304
rect 13235 -1320 13273 -1304
rect 13307 -1320 13350 -1286
rect 12384 -1326 13350 -1320
rect 13554 -1062 14344 -1024
rect 13554 -1096 13932 -1062
rect 13966 -1096 14344 -1062
rect 13554 -1134 14344 -1096
rect 13554 -1168 13932 -1134
rect 13966 -1168 14344 -1134
rect 13554 -1206 14344 -1168
rect 13554 -1240 13932 -1206
rect 13966 -1240 14344 -1206
rect 13554 -1278 14344 -1240
rect 13554 -1286 13932 -1278
rect 13554 -1320 13653 -1286
rect 13687 -1320 13725 -1286
rect 13759 -1312 13932 -1286
rect 13966 -1286 14344 -1278
rect 13966 -1312 14139 -1286
rect 13759 -1320 14139 -1312
rect 14173 -1320 14211 -1286
rect 14245 -1320 14344 -1286
rect 4836 -1414 5626 -1384
rect 4836 -1448 4842 -1414
rect 4876 -1448 5100 -1414
rect 5134 -1422 5328 -1414
rect 5134 -1448 5214 -1422
rect 4836 -1456 5214 -1448
rect 5248 -1448 5328 -1422
rect 5362 -1448 5586 -1414
rect 5620 -1448 5626 -1414
rect 5248 -1456 5626 -1448
rect 4836 -1486 5626 -1456
rect 4836 -1520 4842 -1486
rect 4876 -1520 5100 -1486
rect 5134 -1494 5328 -1486
rect 5134 -1520 5214 -1494
rect 4836 -1528 5214 -1520
rect 5248 -1520 5328 -1494
rect 5362 -1520 5586 -1486
rect 5620 -1520 5626 -1486
rect 5248 -1528 5626 -1520
rect 4836 -1566 5626 -1528
rect 4836 -1600 5214 -1566
rect 5248 -1600 5626 -1566
rect 4836 -1638 5626 -1600
rect 4836 -1672 5214 -1638
rect 5248 -1672 5626 -1638
rect 4570 -1702 4766 -1694
rect 4570 -1754 4577 -1702
rect 4629 -1754 4641 -1702
rect 4693 -1754 4705 -1702
rect 4757 -1754 4766 -1702
rect 4570 -1764 4766 -1754
rect 4836 -1710 5626 -1672
rect 5774 -1414 5820 -1367
rect 5774 -1448 5780 -1414
rect 5814 -1448 5820 -1414
rect 5774 -1486 5820 -1448
rect 5774 -1520 5780 -1486
rect 5814 -1520 5820 -1486
rect 5774 -1694 5820 -1520
rect 6032 -1414 6078 -1367
rect 6032 -1448 6038 -1414
rect 6072 -1448 6078 -1414
rect 6032 -1486 6078 -1448
rect 6032 -1520 6038 -1486
rect 6072 -1520 6078 -1486
rect 4836 -1744 5214 -1710
rect 5248 -1744 5626 -1710
rect 4313 -2003 4509 -1995
rect 4313 -2055 4320 -2003
rect 4372 -2055 4384 -2003
rect 4436 -2055 4448 -2003
rect 4500 -2055 4509 -2003
rect 4313 -2065 4509 -2055
rect 4127 -2404 4133 -2370
rect 4167 -2404 4173 -2370
rect 4127 -2442 4173 -2404
rect 4127 -2476 4133 -2442
rect 4167 -2476 4173 -2442
rect 4127 -2523 4173 -2476
rect 4385 -2370 4431 -2065
rect 4385 -2404 4391 -2370
rect 4425 -2404 4431 -2370
rect 4385 -2442 4431 -2404
rect 4385 -2476 4391 -2442
rect 4425 -2476 4431 -2442
rect 4385 -2523 4431 -2476
rect 4643 -2370 4689 -1764
rect 4643 -2404 4649 -2370
rect 4683 -2404 4689 -2370
rect 4643 -2442 4689 -2404
rect 4643 -2476 4649 -2442
rect 4683 -2476 4689 -2442
rect 4643 -2523 4689 -2476
rect 4836 -1782 5626 -1744
rect 5697 -1702 5893 -1694
rect 5697 -1754 5706 -1702
rect 5758 -1754 5770 -1702
rect 5822 -1754 5834 -1702
rect 5886 -1754 5893 -1702
rect 5697 -1764 5893 -1754
rect 4836 -1816 5214 -1782
rect 5248 -1816 5626 -1782
rect 4836 -1854 5626 -1816
rect 4836 -1888 5214 -1854
rect 5248 -1888 5626 -1854
rect 4836 -1926 5626 -1888
rect 4836 -1960 5214 -1926
rect 5248 -1960 5626 -1926
rect 4836 -1998 5626 -1960
rect 4836 -2032 5214 -1998
rect 5248 -2032 5626 -1998
rect 4836 -2070 5626 -2032
rect 4836 -2104 5214 -2070
rect 5248 -2104 5626 -2070
rect 4836 -2142 5626 -2104
rect 4836 -2176 5214 -2142
rect 5248 -2176 5626 -2142
rect 4836 -2214 5626 -2176
rect 4836 -2248 5214 -2214
rect 5248 -2248 5626 -2214
rect 4836 -2286 5626 -2248
rect 4836 -2320 5214 -2286
rect 5248 -2320 5626 -2286
rect 4836 -2358 5626 -2320
rect 4836 -2370 5214 -2358
rect 4836 -2404 4842 -2370
rect 4876 -2404 5100 -2370
rect 5134 -2392 5214 -2370
rect 5248 -2370 5626 -2358
rect 5248 -2392 5328 -2370
rect 5134 -2404 5328 -2392
rect 5362 -2404 5586 -2370
rect 5620 -2404 5626 -2370
rect 4836 -2430 5626 -2404
rect 4836 -2442 5214 -2430
rect 4836 -2476 4842 -2442
rect 4876 -2476 5100 -2442
rect 5134 -2464 5214 -2442
rect 5248 -2442 5626 -2430
rect 5248 -2464 5328 -2442
rect 5134 -2476 5328 -2464
rect 5362 -2476 5586 -2442
rect 5620 -2476 5626 -2442
rect 4836 -2502 5626 -2476
rect 833 -2570 1269 -2536
rect 4836 -2536 5214 -2502
rect 5248 -2536 5626 -2502
rect 5774 -2370 5820 -1764
rect 6032 -1995 6078 -1520
rect 6290 -1414 6336 -1367
rect 6290 -1448 6296 -1414
rect 6330 -1448 6336 -1414
rect 6290 -1486 6336 -1448
rect 6290 -1520 6296 -1486
rect 6330 -1520 6336 -1486
rect 6290 -1694 6336 -1520
rect 6548 -1414 6594 -1367
rect 6548 -1448 6554 -1414
rect 6588 -1448 6594 -1414
rect 6548 -1486 6594 -1448
rect 6548 -1520 6554 -1486
rect 6588 -1520 6594 -1486
rect 6214 -1702 6410 -1694
rect 6214 -1754 6223 -1702
rect 6275 -1754 6287 -1702
rect 6339 -1754 6351 -1702
rect 6403 -1754 6410 -1702
rect 6214 -1764 6410 -1754
rect 5954 -2003 6150 -1995
rect 5954 -2055 5963 -2003
rect 6015 -2055 6027 -2003
rect 6079 -2055 6091 -2003
rect 6143 -2055 6150 -2003
rect 5954 -2065 6150 -2055
rect 5774 -2404 5780 -2370
rect 5814 -2404 5820 -2370
rect 5774 -2442 5820 -2404
rect 5774 -2476 5780 -2442
rect 5814 -2476 5820 -2442
rect 5774 -2523 5820 -2476
rect 6032 -2370 6078 -2065
rect 6032 -2404 6038 -2370
rect 6072 -2404 6078 -2370
rect 6032 -2442 6078 -2404
rect 6032 -2476 6038 -2442
rect 6072 -2476 6078 -2442
rect 6032 -2523 6078 -2476
rect 6290 -2370 6336 -1764
rect 6548 -1995 6594 -1520
rect 6806 -1414 6852 -1367
rect 6806 -1448 6812 -1414
rect 6846 -1448 6852 -1414
rect 6806 -1486 6852 -1448
rect 6806 -1520 6812 -1486
rect 6846 -1520 6852 -1486
rect 6806 -1694 6852 -1520
rect 7000 -1414 7046 -1367
rect 7000 -1448 7006 -1414
rect 7040 -1448 7046 -1414
rect 7000 -1486 7046 -1448
rect 7000 -1520 7006 -1486
rect 7040 -1520 7046 -1486
rect 6731 -1702 6927 -1694
rect 6731 -1754 6740 -1702
rect 6792 -1754 6804 -1702
rect 6856 -1754 6868 -1702
rect 6920 -1754 6927 -1702
rect 6731 -1764 6927 -1754
rect 6471 -2003 6667 -1995
rect 6471 -2055 6480 -2003
rect 6532 -2055 6544 -2003
rect 6596 -2055 6608 -2003
rect 6660 -2055 6667 -2003
rect 6471 -2065 6667 -2055
rect 6290 -2404 6296 -2370
rect 6330 -2404 6336 -2370
rect 6290 -2442 6336 -2404
rect 6290 -2476 6296 -2442
rect 6330 -2476 6336 -2442
rect 6290 -2523 6336 -2476
rect 6548 -2370 6594 -2065
rect 6548 -2404 6554 -2370
rect 6588 -2404 6594 -2370
rect 6548 -2442 6594 -2404
rect 6548 -2476 6554 -2442
rect 6588 -2476 6594 -2442
rect 6548 -2523 6594 -2476
rect 6806 -2370 6852 -1764
rect 7000 -1834 7046 -1520
rect 7258 -1414 7304 -1367
rect 7258 -1448 7264 -1414
rect 7298 -1448 7304 -1414
rect 7258 -1486 7304 -1448
rect 7258 -1520 7264 -1486
rect 7298 -1520 7304 -1486
rect 6926 -1842 7122 -1834
rect 6926 -1894 6933 -1842
rect 6985 -1894 6997 -1842
rect 7049 -1894 7061 -1842
rect 7113 -1894 7122 -1842
rect 6926 -1904 7122 -1894
rect 6806 -2404 6812 -2370
rect 6846 -2404 6852 -2370
rect 6806 -2442 6852 -2404
rect 6806 -2476 6812 -2442
rect 6846 -2476 6852 -2442
rect 6806 -2523 6852 -2476
rect 7000 -2370 7046 -1904
rect 7258 -2139 7304 -1520
rect 7516 -1414 7562 -1367
rect 7516 -1448 7522 -1414
rect 7556 -1448 7562 -1414
rect 7516 -1486 7562 -1448
rect 7516 -1520 7522 -1486
rect 7556 -1520 7562 -1486
rect 7516 -1834 7562 -1520
rect 7774 -1414 7820 -1367
rect 7774 -1448 7780 -1414
rect 7814 -1448 7820 -1414
rect 7774 -1486 7820 -1448
rect 7774 -1520 7780 -1486
rect 7814 -1520 7820 -1486
rect 7443 -1842 7639 -1834
rect 7443 -1894 7450 -1842
rect 7502 -1894 7514 -1842
rect 7566 -1894 7578 -1842
rect 7630 -1894 7639 -1842
rect 7443 -1904 7639 -1894
rect 7184 -2147 7380 -2139
rect 7184 -2199 7191 -2147
rect 7243 -2199 7255 -2147
rect 7307 -2199 7319 -2147
rect 7371 -2199 7380 -2147
rect 7184 -2209 7380 -2199
rect 7000 -2404 7006 -2370
rect 7040 -2404 7046 -2370
rect 7000 -2442 7046 -2404
rect 7000 -2476 7006 -2442
rect 7040 -2476 7046 -2442
rect 7000 -2523 7046 -2476
rect 7258 -2370 7304 -2209
rect 7258 -2404 7264 -2370
rect 7298 -2404 7304 -2370
rect 7258 -2442 7304 -2404
rect 7258 -2476 7264 -2442
rect 7298 -2476 7304 -2442
rect 7258 -2523 7304 -2476
rect 7516 -2370 7562 -1904
rect 7774 -2139 7820 -1520
rect 7968 -1414 8014 -1367
rect 7968 -1448 7974 -1414
rect 8008 -1448 8014 -1414
rect 7968 -1486 8014 -1448
rect 7968 -1520 7974 -1486
rect 8008 -1520 8014 -1486
rect 7968 -1694 8014 -1520
rect 8226 -1414 8272 -1367
rect 8226 -1448 8232 -1414
rect 8266 -1448 8272 -1414
rect 8226 -1486 8272 -1448
rect 8226 -1520 8232 -1486
rect 8266 -1520 8272 -1486
rect 7891 -1702 8087 -1694
rect 7891 -1754 7900 -1702
rect 7952 -1754 7964 -1702
rect 8016 -1754 8028 -1702
rect 8080 -1754 8087 -1702
rect 7891 -1764 8087 -1754
rect 7701 -2147 7897 -2139
rect 7701 -2199 7708 -2147
rect 7760 -2199 7772 -2147
rect 7824 -2199 7836 -2147
rect 7888 -2199 7897 -2147
rect 7701 -2209 7897 -2199
rect 7516 -2404 7522 -2370
rect 7556 -2404 7562 -2370
rect 7516 -2442 7562 -2404
rect 7516 -2476 7522 -2442
rect 7556 -2476 7562 -2442
rect 7516 -2523 7562 -2476
rect 7774 -2370 7820 -2209
rect 7774 -2404 7780 -2370
rect 7814 -2404 7820 -2370
rect 7774 -2442 7820 -2404
rect 7774 -2476 7780 -2442
rect 7814 -2476 7820 -2442
rect 7774 -2523 7820 -2476
rect 7968 -2370 8014 -1764
rect 8226 -1995 8272 -1520
rect 8484 -1414 8530 -1367
rect 8484 -1448 8490 -1414
rect 8524 -1448 8530 -1414
rect 8484 -1486 8530 -1448
rect 8484 -1520 8490 -1486
rect 8524 -1520 8530 -1486
rect 8484 -1694 8530 -1520
rect 8742 -1414 8788 -1367
rect 8742 -1448 8748 -1414
rect 8782 -1448 8788 -1414
rect 8742 -1486 8788 -1448
rect 8742 -1520 8748 -1486
rect 8782 -1520 8788 -1486
rect 8408 -1702 8604 -1694
rect 8408 -1754 8417 -1702
rect 8469 -1754 8481 -1702
rect 8533 -1754 8545 -1702
rect 8597 -1754 8604 -1702
rect 8408 -1764 8604 -1754
rect 8148 -2003 8344 -1995
rect 8148 -2055 8157 -2003
rect 8209 -2055 8221 -2003
rect 8273 -2055 8285 -2003
rect 8337 -2055 8344 -2003
rect 8148 -2065 8344 -2055
rect 7968 -2404 7974 -2370
rect 8008 -2404 8014 -2370
rect 7968 -2442 8014 -2404
rect 7968 -2476 7974 -2442
rect 8008 -2476 8014 -2442
rect 7968 -2523 8014 -2476
rect 8226 -2370 8272 -2065
rect 8226 -2404 8232 -2370
rect 8266 -2404 8272 -2370
rect 8226 -2442 8272 -2404
rect 8226 -2476 8232 -2442
rect 8266 -2476 8272 -2442
rect 8226 -2523 8272 -2476
rect 8484 -2370 8530 -1764
rect 8742 -1995 8788 -1520
rect 9000 -1414 9046 -1367
rect 9000 -1448 9006 -1414
rect 9040 -1448 9046 -1414
rect 9000 -1486 9046 -1448
rect 9000 -1520 9006 -1486
rect 9040 -1520 9046 -1486
rect 9000 -1694 9046 -1520
rect 9194 -1384 9573 -1350
rect 9607 -1384 9986 -1350
rect 13554 -1350 14344 -1320
rect 14547 -1074 15513 -1056
rect 14547 -1126 14597 -1074
rect 14649 -1126 14661 -1074
rect 14713 -1126 14725 -1074
rect 14777 -1126 14793 -1074
rect 14845 -1126 14857 -1074
rect 14909 -1126 14921 -1074
rect 14973 -1126 15083 -1074
rect 15135 -1126 15147 -1074
rect 15199 -1126 15211 -1074
rect 15263 -1126 15279 -1074
rect 15331 -1126 15343 -1074
rect 15395 -1126 15407 -1074
rect 15459 -1126 15513 -1074
rect 14547 -1252 15513 -1126
rect 14547 -1286 14597 -1252
rect 14547 -1320 14590 -1286
rect 14649 -1304 14661 -1252
rect 14713 -1304 14725 -1252
rect 14777 -1304 14793 -1252
rect 14845 -1286 14857 -1252
rect 14909 -1286 14921 -1252
rect 14845 -1304 14848 -1286
rect 14909 -1304 14920 -1286
rect 14973 -1304 15083 -1252
rect 15135 -1286 15147 -1252
rect 15199 -1286 15211 -1252
rect 15140 -1304 15147 -1286
rect 15263 -1304 15279 -1252
rect 15331 -1304 15343 -1252
rect 15395 -1286 15407 -1252
rect 15459 -1286 15513 -1252
rect 15398 -1304 15407 -1286
rect 14624 -1320 14662 -1304
rect 14696 -1320 14848 -1304
rect 14882 -1320 14920 -1304
rect 14954 -1320 15106 -1304
rect 15140 -1320 15178 -1304
rect 15212 -1320 15364 -1304
rect 15398 -1320 15436 -1304
rect 15470 -1320 15513 -1286
rect 14547 -1326 15513 -1320
rect 15590 -1238 15651 -1006
rect 15773 -923 16481 -917
rect 15773 -957 15816 -923
rect 15850 -957 15888 -923
rect 15922 -957 16074 -923
rect 16108 -957 16146 -923
rect 16180 -957 16332 -923
rect 16366 -957 16404 -923
rect 16438 -957 16481 -923
rect 15773 -1074 16481 -957
rect 15773 -1126 15811 -1074
rect 15863 -1126 15875 -1074
rect 15927 -1126 15939 -1074
rect 15991 -1126 16007 -1074
rect 16059 -1126 16071 -1074
rect 16123 -1126 16135 -1074
rect 16187 -1126 16199 -1074
rect 16251 -1126 16267 -1074
rect 16319 -1126 16331 -1074
rect 16383 -1126 16395 -1074
rect 16447 -1126 16481 -1074
rect 15773 -1144 16481 -1126
rect 16603 -923 17707 -917
rect 16603 -957 16784 -923
rect 16818 -936 16856 -923
rect 16890 -936 17042 -923
rect 17076 -936 17114 -923
rect 17148 -936 17300 -923
rect 17334 -936 17372 -923
rect 17406 -936 17558 -923
rect 17592 -936 17630 -923
rect 16847 -957 16856 -936
rect 16603 -988 16795 -957
rect 16847 -988 16859 -957
rect 16911 -988 16923 -936
rect 16975 -988 16991 -936
rect 17107 -957 17114 -936
rect 17043 -988 17055 -957
rect 17107 -988 17119 -957
rect 17171 -988 17281 -936
rect 17334 -957 17345 -936
rect 17406 -957 17409 -936
rect 17333 -988 17345 -957
rect 17397 -988 17409 -957
rect 17461 -988 17477 -936
rect 17529 -988 17541 -936
rect 17593 -988 17605 -936
rect 17664 -957 17707 -923
rect 17657 -988 17707 -957
rect 16603 -1006 17707 -988
rect 17911 -918 18347 -880
rect 17911 -923 18290 -918
rect 17911 -957 18010 -923
rect 18044 -957 18082 -923
rect 18116 -952 18290 -923
rect 18324 -952 18347 -918
rect 18116 -957 18347 -952
rect 17911 -990 18347 -957
rect 16603 -1238 16664 -1006
rect 17911 -1024 18290 -990
rect 18324 -1024 18347 -990
rect 15590 -1286 16664 -1238
rect 15590 -1320 15816 -1286
rect 15850 -1320 15888 -1286
rect 15922 -1320 16074 -1286
rect 16108 -1320 16146 -1286
rect 16180 -1320 16332 -1286
rect 16366 -1320 16404 -1286
rect 16438 -1320 16664 -1286
rect 15590 -1326 16664 -1320
rect 16741 -1074 17707 -1056
rect 16741 -1126 16795 -1074
rect 16847 -1126 16859 -1074
rect 16911 -1126 16923 -1074
rect 16975 -1126 16991 -1074
rect 17043 -1126 17055 -1074
rect 17107 -1126 17119 -1074
rect 17171 -1126 17281 -1074
rect 17333 -1126 17345 -1074
rect 17397 -1126 17409 -1074
rect 17461 -1126 17477 -1074
rect 17529 -1126 17541 -1074
rect 17593 -1126 17605 -1074
rect 17657 -1126 17707 -1074
rect 16741 -1252 17707 -1126
rect 16741 -1286 16795 -1252
rect 16847 -1286 16859 -1252
rect 16741 -1320 16784 -1286
rect 16847 -1304 16856 -1286
rect 16911 -1304 16923 -1252
rect 16975 -1304 16991 -1252
rect 17043 -1286 17055 -1252
rect 17107 -1286 17119 -1252
rect 17107 -1304 17114 -1286
rect 17171 -1304 17281 -1252
rect 17333 -1286 17345 -1252
rect 17397 -1286 17409 -1252
rect 17334 -1304 17345 -1286
rect 17406 -1304 17409 -1286
rect 17461 -1304 17477 -1252
rect 17529 -1304 17541 -1252
rect 17593 -1304 17605 -1252
rect 17657 -1286 17707 -1252
rect 16818 -1320 16856 -1304
rect 16890 -1320 17042 -1304
rect 17076 -1320 17114 -1304
rect 17148 -1320 17300 -1304
rect 17334 -1320 17372 -1304
rect 17406 -1320 17558 -1304
rect 17592 -1320 17630 -1304
rect 17664 -1320 17707 -1286
rect 16741 -1326 17707 -1320
rect 17911 -1062 18347 -1024
rect 17911 -1096 18290 -1062
rect 18324 -1096 18347 -1062
rect 17911 -1134 18347 -1096
rect 17911 -1168 18290 -1134
rect 18324 -1168 18347 -1134
rect 17911 -1206 18347 -1168
rect 17911 -1240 18290 -1206
rect 18324 -1240 18347 -1206
rect 17911 -1278 18347 -1240
rect 17911 -1286 18290 -1278
rect 17911 -1320 18010 -1286
rect 18044 -1320 18082 -1286
rect 18116 -1312 18290 -1286
rect 18324 -1312 18347 -1278
rect 18116 -1320 18347 -1312
rect 9194 -1414 9986 -1384
rect 9194 -1448 9200 -1414
rect 9234 -1448 9458 -1414
rect 9492 -1422 9688 -1414
rect 9492 -1448 9573 -1422
rect 9194 -1456 9573 -1448
rect 9607 -1448 9688 -1422
rect 9722 -1448 9946 -1414
rect 9980 -1448 9986 -1414
rect 9607 -1456 9986 -1448
rect 9194 -1486 9986 -1456
rect 9194 -1520 9200 -1486
rect 9234 -1520 9458 -1486
rect 9492 -1494 9688 -1486
rect 9492 -1520 9573 -1494
rect 9194 -1528 9573 -1520
rect 9607 -1520 9688 -1494
rect 9722 -1520 9946 -1486
rect 9980 -1520 9986 -1486
rect 9607 -1528 9986 -1520
rect 9194 -1566 9986 -1528
rect 9194 -1600 9573 -1566
rect 9607 -1600 9986 -1566
rect 9194 -1638 9986 -1600
rect 9194 -1672 9573 -1638
rect 9607 -1672 9986 -1638
rect 8923 -1702 9119 -1694
rect 8923 -1754 8932 -1702
rect 8984 -1754 8996 -1702
rect 9048 -1754 9060 -1702
rect 9112 -1754 9119 -1702
rect 8923 -1764 9119 -1754
rect 9194 -1710 9986 -1672
rect 10134 -1414 10180 -1367
rect 10134 -1448 10140 -1414
rect 10174 -1448 10180 -1414
rect 10134 -1486 10180 -1448
rect 10134 -1520 10140 -1486
rect 10174 -1520 10180 -1486
rect 10134 -1694 10180 -1520
rect 10392 -1414 10438 -1367
rect 10392 -1448 10398 -1414
rect 10432 -1448 10438 -1414
rect 10392 -1486 10438 -1448
rect 10392 -1520 10398 -1486
rect 10432 -1520 10438 -1486
rect 9194 -1744 9573 -1710
rect 9607 -1744 9986 -1710
rect 8665 -2003 8861 -1995
rect 8665 -2055 8674 -2003
rect 8726 -2055 8738 -2003
rect 8790 -2055 8802 -2003
rect 8854 -2055 8861 -2003
rect 8665 -2065 8861 -2055
rect 8484 -2404 8490 -2370
rect 8524 -2404 8530 -2370
rect 8484 -2442 8530 -2404
rect 8484 -2476 8490 -2442
rect 8524 -2476 8530 -2442
rect 8484 -2523 8530 -2476
rect 8742 -2370 8788 -2065
rect 8742 -2404 8748 -2370
rect 8782 -2404 8788 -2370
rect 8742 -2442 8788 -2404
rect 8742 -2476 8748 -2442
rect 8782 -2476 8788 -2442
rect 8742 -2523 8788 -2476
rect 9000 -2370 9046 -1764
rect 9000 -2404 9006 -2370
rect 9040 -2404 9046 -2370
rect 9000 -2442 9046 -2404
rect 9000 -2476 9006 -2442
rect 9040 -2476 9046 -2442
rect 9000 -2523 9046 -2476
rect 9194 -1782 9986 -1744
rect 10061 -1702 10257 -1694
rect 10061 -1754 10068 -1702
rect 10120 -1754 10132 -1702
rect 10184 -1754 10196 -1702
rect 10248 -1754 10257 -1702
rect 10061 -1764 10257 -1754
rect 9194 -1816 9573 -1782
rect 9607 -1816 9986 -1782
rect 9194 -1854 9986 -1816
rect 9194 -1888 9573 -1854
rect 9607 -1888 9986 -1854
rect 9194 -1926 9986 -1888
rect 9194 -1960 9573 -1926
rect 9607 -1960 9986 -1926
rect 9194 -1998 9986 -1960
rect 9194 -2032 9573 -1998
rect 9607 -2032 9986 -1998
rect 9194 -2070 9986 -2032
rect 9194 -2104 9573 -2070
rect 9607 -2104 9986 -2070
rect 9194 -2142 9986 -2104
rect 9194 -2176 9573 -2142
rect 9607 -2176 9986 -2142
rect 9194 -2214 9986 -2176
rect 9194 -2248 9573 -2214
rect 9607 -2248 9986 -2214
rect 9194 -2286 9986 -2248
rect 9194 -2320 9573 -2286
rect 9607 -2320 9986 -2286
rect 9194 -2358 9986 -2320
rect 9194 -2370 9573 -2358
rect 9194 -2404 9200 -2370
rect 9234 -2404 9458 -2370
rect 9492 -2392 9573 -2370
rect 9607 -2370 9986 -2358
rect 9607 -2392 9688 -2370
rect 9492 -2404 9688 -2392
rect 9722 -2404 9946 -2370
rect 9980 -2404 9986 -2370
rect 9194 -2430 9986 -2404
rect 9194 -2442 9573 -2430
rect 9194 -2476 9200 -2442
rect 9234 -2476 9458 -2442
rect 9492 -2464 9573 -2442
rect 9607 -2442 9986 -2430
rect 9607 -2464 9688 -2442
rect 9492 -2476 9688 -2464
rect 9722 -2476 9946 -2442
rect 9980 -2476 9986 -2442
rect 9194 -2502 9986 -2476
rect 833 -2574 1064 -2570
rect 833 -2608 856 -2574
rect 890 -2604 1064 -2574
rect 1098 -2604 1136 -2570
rect 1170 -2604 1269 -2570
rect 890 -2608 1269 -2604
rect 833 -2646 1269 -2608
rect 833 -2680 856 -2646
rect 890 -2680 1269 -2646
rect 1473 -2570 2577 -2564
rect 1473 -2604 1516 -2570
rect 1550 -2583 1588 -2570
rect 1622 -2583 1774 -2570
rect 1808 -2583 1846 -2570
rect 1880 -2583 2032 -2570
rect 2066 -2583 2104 -2570
rect 2138 -2583 2290 -2570
rect 2324 -2583 2362 -2570
rect 1473 -2635 1523 -2604
rect 1575 -2635 1587 -2583
rect 1639 -2635 1651 -2583
rect 1703 -2635 1719 -2583
rect 1771 -2604 1774 -2583
rect 1835 -2604 1846 -2583
rect 1771 -2635 1783 -2604
rect 1835 -2635 1847 -2604
rect 1899 -2635 2009 -2583
rect 2066 -2604 2073 -2583
rect 2061 -2635 2073 -2604
rect 2125 -2635 2137 -2604
rect 2189 -2635 2205 -2583
rect 2257 -2635 2269 -2583
rect 2324 -2604 2333 -2583
rect 2396 -2604 2577 -2570
rect 2321 -2635 2333 -2604
rect 2385 -2635 2577 -2604
rect 1473 -2653 2577 -2635
rect 833 -2718 1269 -2680
rect 833 -2752 856 -2718
rect 890 -2752 1269 -2718
rect 833 -2790 1269 -2752
rect 833 -2824 856 -2790
rect 890 -2824 1269 -2790
rect 833 -2862 1269 -2824
rect 833 -2896 856 -2862
rect 890 -2896 1269 -2862
rect 833 -2933 1269 -2896
rect 833 -2934 1064 -2933
rect 833 -2968 856 -2934
rect 890 -2967 1064 -2934
rect 1098 -2967 1136 -2933
rect 1170 -2967 1269 -2933
rect 890 -2968 1269 -2967
rect 833 -3006 1269 -2968
rect 1473 -2721 2439 -2703
rect 1473 -2773 1523 -2721
rect 1575 -2773 1587 -2721
rect 1639 -2773 1651 -2721
rect 1703 -2773 1719 -2721
rect 1771 -2773 1783 -2721
rect 1835 -2773 1847 -2721
rect 1899 -2773 2009 -2721
rect 2061 -2773 2073 -2721
rect 2125 -2773 2137 -2721
rect 2189 -2773 2205 -2721
rect 2257 -2773 2269 -2721
rect 2321 -2773 2333 -2721
rect 2385 -2773 2439 -2721
rect 1473 -2899 2439 -2773
rect 1473 -2933 1523 -2899
rect 1473 -2967 1516 -2933
rect 1575 -2951 1587 -2899
rect 1639 -2951 1651 -2899
rect 1703 -2951 1719 -2899
rect 1771 -2933 1783 -2899
rect 1835 -2933 1847 -2899
rect 1771 -2951 1774 -2933
rect 1835 -2951 1846 -2933
rect 1899 -2951 2009 -2899
rect 2061 -2933 2073 -2899
rect 2125 -2933 2137 -2899
rect 2066 -2951 2073 -2933
rect 2189 -2951 2205 -2899
rect 2257 -2951 2269 -2899
rect 2321 -2933 2333 -2899
rect 2385 -2933 2439 -2899
rect 2324 -2951 2333 -2933
rect 1550 -2967 1588 -2951
rect 1622 -2967 1774 -2951
rect 1808 -2967 1846 -2951
rect 1880 -2967 2032 -2951
rect 2066 -2967 2104 -2951
rect 2138 -2967 2290 -2951
rect 2324 -2967 2362 -2951
rect 2396 -2967 2439 -2933
rect 1473 -2973 2439 -2967
rect 2516 -2885 2577 -2653
rect 2699 -2570 3407 -2564
rect 2699 -2604 2742 -2570
rect 2776 -2604 2814 -2570
rect 2848 -2604 3000 -2570
rect 3034 -2604 3072 -2570
rect 3106 -2604 3258 -2570
rect 3292 -2604 3330 -2570
rect 3364 -2604 3407 -2570
rect 2699 -2721 3407 -2604
rect 2699 -2773 2733 -2721
rect 2785 -2773 2797 -2721
rect 2849 -2773 2861 -2721
rect 2913 -2773 2929 -2721
rect 2981 -2773 2993 -2721
rect 3045 -2773 3057 -2721
rect 3109 -2773 3121 -2721
rect 3173 -2773 3189 -2721
rect 3241 -2773 3253 -2721
rect 3305 -2773 3317 -2721
rect 3369 -2773 3407 -2721
rect 2699 -2791 3407 -2773
rect 3529 -2570 4633 -2564
rect 3529 -2604 3710 -2570
rect 3744 -2583 3782 -2570
rect 3816 -2583 3968 -2570
rect 4002 -2583 4040 -2570
rect 4074 -2583 4226 -2570
rect 4260 -2583 4298 -2570
rect 4332 -2583 4484 -2570
rect 4518 -2583 4556 -2570
rect 3773 -2604 3782 -2583
rect 3529 -2635 3721 -2604
rect 3773 -2635 3785 -2604
rect 3837 -2635 3849 -2583
rect 3901 -2635 3917 -2583
rect 4033 -2604 4040 -2583
rect 3969 -2635 3981 -2604
rect 4033 -2635 4045 -2604
rect 4097 -2635 4207 -2583
rect 4260 -2604 4271 -2583
rect 4332 -2604 4335 -2583
rect 4259 -2635 4271 -2604
rect 4323 -2635 4335 -2604
rect 4387 -2635 4403 -2583
rect 4455 -2635 4467 -2583
rect 4519 -2635 4531 -2583
rect 4590 -2604 4633 -2570
rect 4583 -2635 4633 -2604
rect 3529 -2653 4633 -2635
rect 4836 -2570 5626 -2536
rect 9194 -2536 9573 -2502
rect 9607 -2536 9986 -2502
rect 10134 -2370 10180 -1764
rect 10392 -1995 10438 -1520
rect 10650 -1414 10696 -1367
rect 10650 -1448 10656 -1414
rect 10690 -1448 10696 -1414
rect 10650 -1486 10696 -1448
rect 10650 -1520 10656 -1486
rect 10690 -1520 10696 -1486
rect 10650 -1694 10696 -1520
rect 10908 -1414 10954 -1367
rect 10908 -1448 10914 -1414
rect 10948 -1448 10954 -1414
rect 10908 -1486 10954 -1448
rect 10908 -1520 10914 -1486
rect 10948 -1520 10954 -1486
rect 10576 -1702 10772 -1694
rect 10576 -1754 10583 -1702
rect 10635 -1754 10647 -1702
rect 10699 -1754 10711 -1702
rect 10763 -1754 10772 -1702
rect 10576 -1764 10772 -1754
rect 10319 -2003 10515 -1995
rect 10319 -2055 10326 -2003
rect 10378 -2055 10390 -2003
rect 10442 -2055 10454 -2003
rect 10506 -2055 10515 -2003
rect 10319 -2065 10515 -2055
rect 10134 -2404 10140 -2370
rect 10174 -2404 10180 -2370
rect 10134 -2442 10180 -2404
rect 10134 -2476 10140 -2442
rect 10174 -2476 10180 -2442
rect 10134 -2523 10180 -2476
rect 10392 -2370 10438 -2065
rect 10392 -2404 10398 -2370
rect 10432 -2404 10438 -2370
rect 10392 -2442 10438 -2404
rect 10392 -2476 10398 -2442
rect 10432 -2476 10438 -2442
rect 10392 -2523 10438 -2476
rect 10650 -2370 10696 -1764
rect 10908 -1995 10954 -1520
rect 11166 -1414 11212 -1367
rect 11166 -1448 11172 -1414
rect 11206 -1448 11212 -1414
rect 11166 -1486 11212 -1448
rect 11166 -1520 11172 -1486
rect 11206 -1520 11212 -1486
rect 11166 -1694 11212 -1520
rect 11360 -1414 11406 -1367
rect 11360 -1448 11366 -1414
rect 11400 -1448 11406 -1414
rect 11360 -1486 11406 -1448
rect 11360 -1520 11366 -1486
rect 11400 -1520 11406 -1486
rect 11093 -1702 11289 -1694
rect 11093 -1754 11100 -1702
rect 11152 -1754 11164 -1702
rect 11216 -1754 11228 -1702
rect 11280 -1754 11289 -1702
rect 11093 -1764 11289 -1754
rect 10836 -2003 11032 -1995
rect 10836 -2055 10843 -2003
rect 10895 -2055 10907 -2003
rect 10959 -2055 10971 -2003
rect 11023 -2055 11032 -2003
rect 10836 -2065 11032 -2055
rect 10650 -2404 10656 -2370
rect 10690 -2404 10696 -2370
rect 10650 -2442 10696 -2404
rect 10650 -2476 10656 -2442
rect 10690 -2476 10696 -2442
rect 10650 -2523 10696 -2476
rect 10908 -2370 10954 -2065
rect 10908 -2404 10914 -2370
rect 10948 -2404 10954 -2370
rect 10908 -2442 10954 -2404
rect 10908 -2476 10914 -2442
rect 10948 -2476 10954 -2442
rect 10908 -2523 10954 -2476
rect 11166 -2370 11212 -1764
rect 11360 -2139 11406 -1520
rect 11618 -1414 11664 -1367
rect 11618 -1448 11624 -1414
rect 11658 -1448 11664 -1414
rect 11618 -1486 11664 -1448
rect 11618 -1520 11624 -1486
rect 11658 -1520 11664 -1486
rect 11618 -1834 11664 -1520
rect 11876 -1414 11922 -1367
rect 11876 -1448 11882 -1414
rect 11916 -1448 11922 -1414
rect 11876 -1486 11922 -1448
rect 11876 -1520 11882 -1486
rect 11916 -1520 11922 -1486
rect 11541 -1842 11737 -1834
rect 11541 -1894 11550 -1842
rect 11602 -1894 11614 -1842
rect 11666 -1894 11678 -1842
rect 11730 -1894 11737 -1842
rect 11541 -1904 11737 -1894
rect 11283 -2147 11479 -2139
rect 11283 -2199 11292 -2147
rect 11344 -2199 11356 -2147
rect 11408 -2199 11420 -2147
rect 11472 -2199 11479 -2147
rect 11283 -2209 11479 -2199
rect 11166 -2404 11172 -2370
rect 11206 -2404 11212 -2370
rect 11166 -2442 11212 -2404
rect 11166 -2476 11172 -2442
rect 11206 -2476 11212 -2442
rect 11166 -2523 11212 -2476
rect 11360 -2370 11406 -2209
rect 11360 -2404 11366 -2370
rect 11400 -2404 11406 -2370
rect 11360 -2442 11406 -2404
rect 11360 -2476 11366 -2442
rect 11400 -2476 11406 -2442
rect 11360 -2523 11406 -2476
rect 11618 -2370 11664 -1904
rect 11876 -2139 11922 -1520
rect 12134 -1414 12180 -1367
rect 12134 -1448 12140 -1414
rect 12174 -1448 12180 -1414
rect 12134 -1486 12180 -1448
rect 12134 -1520 12140 -1486
rect 12174 -1520 12180 -1486
rect 12134 -1834 12180 -1520
rect 12328 -1414 12374 -1367
rect 12328 -1448 12334 -1414
rect 12368 -1448 12374 -1414
rect 12328 -1486 12374 -1448
rect 12328 -1520 12334 -1486
rect 12368 -1520 12374 -1486
rect 12328 -1694 12374 -1520
rect 12586 -1414 12632 -1367
rect 12586 -1448 12592 -1414
rect 12626 -1448 12632 -1414
rect 12586 -1486 12632 -1448
rect 12586 -1520 12592 -1486
rect 12626 -1520 12632 -1486
rect 12253 -1702 12449 -1694
rect 12253 -1754 12260 -1702
rect 12312 -1754 12324 -1702
rect 12376 -1754 12388 -1702
rect 12440 -1754 12449 -1702
rect 12253 -1764 12449 -1754
rect 12058 -1842 12254 -1834
rect 12058 -1894 12067 -1842
rect 12119 -1894 12131 -1842
rect 12183 -1894 12195 -1842
rect 12247 -1894 12254 -1842
rect 12058 -1904 12254 -1894
rect 11800 -2147 11996 -2139
rect 11800 -2199 11809 -2147
rect 11861 -2199 11873 -2147
rect 11925 -2199 11937 -2147
rect 11989 -2199 11996 -2147
rect 11800 -2209 11996 -2199
rect 11618 -2404 11624 -2370
rect 11658 -2404 11664 -2370
rect 11618 -2442 11664 -2404
rect 11618 -2476 11624 -2442
rect 11658 -2476 11664 -2442
rect 11618 -2523 11664 -2476
rect 11876 -2370 11922 -2209
rect 11876 -2404 11882 -2370
rect 11916 -2404 11922 -2370
rect 11876 -2442 11922 -2404
rect 11876 -2476 11882 -2442
rect 11916 -2476 11922 -2442
rect 11876 -2523 11922 -2476
rect 12134 -2370 12180 -1904
rect 12134 -2404 12140 -2370
rect 12174 -2404 12180 -2370
rect 12134 -2442 12180 -2404
rect 12134 -2476 12140 -2442
rect 12174 -2476 12180 -2442
rect 12134 -2523 12180 -2476
rect 12328 -2370 12374 -1764
rect 12586 -1995 12632 -1520
rect 12844 -1414 12890 -1367
rect 12844 -1448 12850 -1414
rect 12884 -1448 12890 -1414
rect 12844 -1486 12890 -1448
rect 12844 -1520 12850 -1486
rect 12884 -1520 12890 -1486
rect 12844 -1694 12890 -1520
rect 13102 -1414 13148 -1367
rect 13102 -1448 13108 -1414
rect 13142 -1448 13148 -1414
rect 13102 -1486 13148 -1448
rect 13102 -1520 13108 -1486
rect 13142 -1520 13148 -1486
rect 12770 -1702 12966 -1694
rect 12770 -1754 12777 -1702
rect 12829 -1754 12841 -1702
rect 12893 -1754 12905 -1702
rect 12957 -1754 12966 -1702
rect 12770 -1764 12966 -1754
rect 12513 -2003 12709 -1995
rect 12513 -2055 12520 -2003
rect 12572 -2055 12584 -2003
rect 12636 -2055 12648 -2003
rect 12700 -2055 12709 -2003
rect 12513 -2065 12709 -2055
rect 12328 -2404 12334 -2370
rect 12368 -2404 12374 -2370
rect 12328 -2442 12374 -2404
rect 12328 -2476 12334 -2442
rect 12368 -2476 12374 -2442
rect 12328 -2523 12374 -2476
rect 12586 -2370 12632 -2065
rect 12586 -2404 12592 -2370
rect 12626 -2404 12632 -2370
rect 12586 -2442 12632 -2404
rect 12586 -2476 12592 -2442
rect 12626 -2476 12632 -2442
rect 12586 -2523 12632 -2476
rect 12844 -2370 12890 -1764
rect 13102 -1995 13148 -1520
rect 13360 -1414 13406 -1367
rect 13360 -1448 13366 -1414
rect 13400 -1448 13406 -1414
rect 13360 -1486 13406 -1448
rect 13360 -1520 13366 -1486
rect 13400 -1520 13406 -1486
rect 13360 -1694 13406 -1520
rect 13554 -1384 13932 -1350
rect 13966 -1384 14344 -1350
rect 17911 -1350 18347 -1320
rect 13554 -1414 14344 -1384
rect 13554 -1448 13560 -1414
rect 13594 -1448 13818 -1414
rect 13852 -1422 14046 -1414
rect 13852 -1448 13932 -1422
rect 13554 -1456 13932 -1448
rect 13966 -1448 14046 -1422
rect 14080 -1448 14304 -1414
rect 14338 -1448 14344 -1414
rect 13966 -1456 14344 -1448
rect 13554 -1486 14344 -1456
rect 13554 -1520 13560 -1486
rect 13594 -1520 13818 -1486
rect 13852 -1494 14046 -1486
rect 13852 -1520 13932 -1494
rect 13554 -1528 13932 -1520
rect 13966 -1520 14046 -1494
rect 14080 -1520 14304 -1486
rect 14338 -1520 14344 -1486
rect 13966 -1528 14344 -1520
rect 13554 -1566 14344 -1528
rect 13554 -1600 13932 -1566
rect 13966 -1600 14344 -1566
rect 13554 -1638 14344 -1600
rect 13554 -1672 13932 -1638
rect 13966 -1672 14344 -1638
rect 13287 -1702 13483 -1694
rect 13287 -1754 13294 -1702
rect 13346 -1754 13358 -1702
rect 13410 -1754 13422 -1702
rect 13474 -1754 13483 -1702
rect 13287 -1764 13483 -1754
rect 13554 -1710 14344 -1672
rect 14491 -1414 14537 -1367
rect 14491 -1448 14497 -1414
rect 14531 -1448 14537 -1414
rect 14491 -1486 14537 -1448
rect 14491 -1520 14497 -1486
rect 14531 -1520 14537 -1486
rect 14491 -1694 14537 -1520
rect 14749 -1414 14795 -1367
rect 14749 -1448 14755 -1414
rect 14789 -1448 14795 -1414
rect 14749 -1486 14795 -1448
rect 14749 -1520 14755 -1486
rect 14789 -1520 14795 -1486
rect 13554 -1744 13932 -1710
rect 13966 -1744 14344 -1710
rect 13030 -2003 13226 -1995
rect 13030 -2055 13037 -2003
rect 13089 -2055 13101 -2003
rect 13153 -2055 13165 -2003
rect 13217 -2055 13226 -2003
rect 13030 -2065 13226 -2055
rect 12844 -2404 12850 -2370
rect 12884 -2404 12890 -2370
rect 12844 -2442 12890 -2404
rect 12844 -2476 12850 -2442
rect 12884 -2476 12890 -2442
rect 12844 -2523 12890 -2476
rect 13102 -2370 13148 -2065
rect 13102 -2404 13108 -2370
rect 13142 -2404 13148 -2370
rect 13102 -2442 13148 -2404
rect 13102 -2476 13108 -2442
rect 13142 -2476 13148 -2442
rect 13102 -2523 13148 -2476
rect 13360 -2370 13406 -1764
rect 13360 -2404 13366 -2370
rect 13400 -2404 13406 -2370
rect 13360 -2442 13406 -2404
rect 13360 -2476 13366 -2442
rect 13400 -2476 13406 -2442
rect 13360 -2523 13406 -2476
rect 13554 -1782 14344 -1744
rect 14414 -1702 14610 -1694
rect 14414 -1754 14423 -1702
rect 14475 -1754 14487 -1702
rect 14539 -1754 14551 -1702
rect 14603 -1754 14610 -1702
rect 14414 -1764 14610 -1754
rect 13554 -1816 13932 -1782
rect 13966 -1816 14344 -1782
rect 13554 -1854 14344 -1816
rect 13554 -1888 13932 -1854
rect 13966 -1888 14344 -1854
rect 13554 -1926 14344 -1888
rect 13554 -1960 13932 -1926
rect 13966 -1960 14344 -1926
rect 13554 -1998 14344 -1960
rect 13554 -2032 13932 -1998
rect 13966 -2032 14344 -1998
rect 13554 -2070 14344 -2032
rect 13554 -2104 13932 -2070
rect 13966 -2104 14344 -2070
rect 13554 -2142 14344 -2104
rect 13554 -2176 13932 -2142
rect 13966 -2176 14344 -2142
rect 13554 -2214 14344 -2176
rect 13554 -2248 13932 -2214
rect 13966 -2248 14344 -2214
rect 13554 -2286 14344 -2248
rect 13554 -2320 13932 -2286
rect 13966 -2320 14344 -2286
rect 13554 -2358 14344 -2320
rect 13554 -2370 13932 -2358
rect 13554 -2404 13560 -2370
rect 13594 -2404 13818 -2370
rect 13852 -2392 13932 -2370
rect 13966 -2370 14344 -2358
rect 13966 -2392 14046 -2370
rect 13852 -2404 14046 -2392
rect 14080 -2404 14304 -2370
rect 14338 -2404 14344 -2370
rect 13554 -2430 14344 -2404
rect 13554 -2442 13932 -2430
rect 13554 -2476 13560 -2442
rect 13594 -2476 13818 -2442
rect 13852 -2464 13932 -2442
rect 13966 -2442 14344 -2430
rect 13966 -2464 14046 -2442
rect 13852 -2476 14046 -2464
rect 14080 -2476 14304 -2442
rect 14338 -2476 14344 -2442
rect 13554 -2502 14344 -2476
rect 4836 -2604 4935 -2570
rect 4969 -2604 5007 -2570
rect 5041 -2574 5421 -2570
rect 5041 -2604 5214 -2574
rect 4836 -2608 5214 -2604
rect 5248 -2604 5421 -2574
rect 5455 -2604 5493 -2570
rect 5527 -2604 5626 -2570
rect 5248 -2608 5626 -2604
rect 4836 -2646 5626 -2608
rect 3529 -2885 3590 -2653
rect 4836 -2680 5214 -2646
rect 5248 -2680 5626 -2646
rect 5830 -2570 6934 -2564
rect 5830 -2604 5873 -2570
rect 5907 -2583 5945 -2570
rect 5979 -2583 6131 -2570
rect 6165 -2583 6203 -2570
rect 6237 -2583 6389 -2570
rect 6423 -2583 6461 -2570
rect 6495 -2583 6647 -2570
rect 6681 -2583 6719 -2570
rect 5830 -2635 5880 -2604
rect 5932 -2635 5944 -2583
rect 5996 -2635 6008 -2583
rect 6060 -2635 6076 -2583
rect 6128 -2604 6131 -2583
rect 6192 -2604 6203 -2583
rect 6128 -2635 6140 -2604
rect 6192 -2635 6204 -2604
rect 6256 -2635 6366 -2583
rect 6423 -2604 6430 -2583
rect 6418 -2635 6430 -2604
rect 6482 -2635 6494 -2604
rect 6546 -2635 6562 -2583
rect 6614 -2635 6626 -2583
rect 6681 -2604 6690 -2583
rect 6753 -2604 6934 -2570
rect 6678 -2635 6690 -2604
rect 6742 -2635 6934 -2604
rect 5830 -2653 6934 -2635
rect 2516 -2933 3590 -2885
rect 2516 -2967 2742 -2933
rect 2776 -2967 2814 -2933
rect 2848 -2967 3000 -2933
rect 3034 -2967 3072 -2933
rect 3106 -2967 3258 -2933
rect 3292 -2967 3330 -2933
rect 3364 -2967 3590 -2933
rect 2516 -2973 3590 -2967
rect 3667 -2721 4633 -2703
rect 3667 -2773 3721 -2721
rect 3773 -2773 3785 -2721
rect 3837 -2773 3849 -2721
rect 3901 -2773 3917 -2721
rect 3969 -2773 3981 -2721
rect 4033 -2773 4045 -2721
rect 4097 -2773 4207 -2721
rect 4259 -2773 4271 -2721
rect 4323 -2773 4335 -2721
rect 4387 -2773 4403 -2721
rect 4455 -2773 4467 -2721
rect 4519 -2773 4531 -2721
rect 4583 -2773 4633 -2721
rect 3667 -2899 4633 -2773
rect 3667 -2933 3721 -2899
rect 3773 -2933 3785 -2899
rect 3667 -2967 3710 -2933
rect 3773 -2951 3782 -2933
rect 3837 -2951 3849 -2899
rect 3901 -2951 3917 -2899
rect 3969 -2933 3981 -2899
rect 4033 -2933 4045 -2899
rect 4033 -2951 4040 -2933
rect 4097 -2951 4207 -2899
rect 4259 -2933 4271 -2899
rect 4323 -2933 4335 -2899
rect 4260 -2951 4271 -2933
rect 4332 -2951 4335 -2933
rect 4387 -2951 4403 -2899
rect 4455 -2951 4467 -2899
rect 4519 -2951 4531 -2899
rect 4583 -2933 4633 -2899
rect 3744 -2967 3782 -2951
rect 3816 -2967 3968 -2951
rect 4002 -2967 4040 -2951
rect 4074 -2967 4226 -2951
rect 4260 -2967 4298 -2951
rect 4332 -2967 4484 -2951
rect 4518 -2967 4556 -2951
rect 4590 -2967 4633 -2933
rect 3667 -2973 4633 -2967
rect 4836 -2718 5626 -2680
rect 4836 -2752 5214 -2718
rect 5248 -2752 5626 -2718
rect 4836 -2790 5626 -2752
rect 4836 -2824 5214 -2790
rect 5248 -2824 5626 -2790
rect 4836 -2862 5626 -2824
rect 4836 -2896 5214 -2862
rect 5248 -2896 5626 -2862
rect 4836 -2933 5626 -2896
rect 4836 -2967 4935 -2933
rect 4969 -2967 5007 -2933
rect 5041 -2934 5421 -2933
rect 5041 -2967 5214 -2934
rect 4836 -2968 5214 -2967
rect 5248 -2967 5421 -2934
rect 5455 -2967 5493 -2933
rect 5527 -2967 5626 -2933
rect 5248 -2968 5626 -2967
rect 833 -3040 856 -3006
rect 890 -3040 1269 -3006
rect 4836 -3006 5626 -2968
rect 5830 -2721 6796 -2703
rect 5830 -2773 5880 -2721
rect 5932 -2773 5944 -2721
rect 5996 -2773 6008 -2721
rect 6060 -2773 6076 -2721
rect 6128 -2773 6140 -2721
rect 6192 -2773 6204 -2721
rect 6256 -2773 6366 -2721
rect 6418 -2773 6430 -2721
rect 6482 -2773 6494 -2721
rect 6546 -2773 6562 -2721
rect 6614 -2773 6626 -2721
rect 6678 -2773 6690 -2721
rect 6742 -2773 6796 -2721
rect 5830 -2899 6796 -2773
rect 5830 -2933 5880 -2899
rect 5830 -2967 5873 -2933
rect 5932 -2951 5944 -2899
rect 5996 -2951 6008 -2899
rect 6060 -2951 6076 -2899
rect 6128 -2933 6140 -2899
rect 6192 -2933 6204 -2899
rect 6128 -2951 6131 -2933
rect 6192 -2951 6203 -2933
rect 6256 -2951 6366 -2899
rect 6418 -2933 6430 -2899
rect 6482 -2933 6494 -2899
rect 6423 -2951 6430 -2933
rect 6546 -2951 6562 -2899
rect 6614 -2951 6626 -2899
rect 6678 -2933 6690 -2899
rect 6742 -2933 6796 -2899
rect 6681 -2951 6690 -2933
rect 5907 -2967 5945 -2951
rect 5979 -2967 6131 -2951
rect 6165 -2967 6203 -2951
rect 6237 -2967 6389 -2951
rect 6423 -2967 6461 -2951
rect 6495 -2967 6647 -2951
rect 6681 -2967 6719 -2951
rect 6753 -2967 6796 -2933
rect 5830 -2973 6796 -2967
rect 6873 -2885 6934 -2653
rect 7056 -2570 7764 -2564
rect 7056 -2604 7099 -2570
rect 7133 -2604 7171 -2570
rect 7205 -2604 7357 -2570
rect 7391 -2604 7429 -2570
rect 7463 -2604 7615 -2570
rect 7649 -2604 7687 -2570
rect 7721 -2604 7764 -2570
rect 7056 -2721 7764 -2604
rect 7056 -2773 7094 -2721
rect 7146 -2773 7158 -2721
rect 7210 -2773 7222 -2721
rect 7274 -2773 7290 -2721
rect 7342 -2773 7354 -2721
rect 7406 -2773 7418 -2721
rect 7470 -2773 7482 -2721
rect 7534 -2773 7550 -2721
rect 7602 -2773 7614 -2721
rect 7666 -2773 7678 -2721
rect 7730 -2773 7764 -2721
rect 7056 -2791 7764 -2773
rect 7886 -2570 8990 -2564
rect 7886 -2604 8067 -2570
rect 8101 -2583 8139 -2570
rect 8173 -2583 8325 -2570
rect 8359 -2583 8397 -2570
rect 8431 -2583 8583 -2570
rect 8617 -2583 8655 -2570
rect 8689 -2583 8841 -2570
rect 8875 -2583 8913 -2570
rect 8130 -2604 8139 -2583
rect 7886 -2635 8078 -2604
rect 8130 -2635 8142 -2604
rect 8194 -2635 8206 -2583
rect 8258 -2635 8274 -2583
rect 8390 -2604 8397 -2583
rect 8326 -2635 8338 -2604
rect 8390 -2635 8402 -2604
rect 8454 -2635 8564 -2583
rect 8617 -2604 8628 -2583
rect 8689 -2604 8692 -2583
rect 8616 -2635 8628 -2604
rect 8680 -2635 8692 -2604
rect 8744 -2635 8760 -2583
rect 8812 -2635 8824 -2583
rect 8876 -2635 8888 -2583
rect 8947 -2604 8990 -2570
rect 8940 -2635 8990 -2604
rect 7886 -2653 8990 -2635
rect 9194 -2570 9986 -2536
rect 13554 -2536 13932 -2502
rect 13966 -2536 14344 -2502
rect 14491 -2370 14537 -1764
rect 14749 -1995 14795 -1520
rect 15007 -1414 15053 -1367
rect 15007 -1448 15013 -1414
rect 15047 -1448 15053 -1414
rect 15007 -1486 15053 -1448
rect 15007 -1520 15013 -1486
rect 15047 -1520 15053 -1486
rect 15007 -1694 15053 -1520
rect 15265 -1414 15311 -1367
rect 15265 -1448 15271 -1414
rect 15305 -1448 15311 -1414
rect 15265 -1486 15311 -1448
rect 15265 -1520 15271 -1486
rect 15305 -1520 15311 -1486
rect 14931 -1702 15127 -1694
rect 14931 -1754 14940 -1702
rect 14992 -1754 15004 -1702
rect 15056 -1754 15068 -1702
rect 15120 -1754 15127 -1702
rect 14931 -1764 15127 -1754
rect 14671 -2003 14867 -1995
rect 14671 -2055 14680 -2003
rect 14732 -2055 14744 -2003
rect 14796 -2055 14808 -2003
rect 14860 -2055 14867 -2003
rect 14671 -2065 14867 -2055
rect 14491 -2404 14497 -2370
rect 14531 -2404 14537 -2370
rect 14491 -2442 14537 -2404
rect 14491 -2476 14497 -2442
rect 14531 -2476 14537 -2442
rect 14491 -2523 14537 -2476
rect 14749 -2370 14795 -2065
rect 14749 -2404 14755 -2370
rect 14789 -2404 14795 -2370
rect 14749 -2442 14795 -2404
rect 14749 -2476 14755 -2442
rect 14789 -2476 14795 -2442
rect 14749 -2523 14795 -2476
rect 15007 -2370 15053 -1764
rect 15265 -1995 15311 -1520
rect 15523 -1414 15569 -1367
rect 15523 -1448 15529 -1414
rect 15563 -1448 15569 -1414
rect 15523 -1486 15569 -1448
rect 15523 -1520 15529 -1486
rect 15563 -1520 15569 -1486
rect 15523 -1694 15569 -1520
rect 15717 -1414 15763 -1367
rect 15717 -1448 15723 -1414
rect 15757 -1448 15763 -1414
rect 15717 -1486 15763 -1448
rect 15717 -1520 15723 -1486
rect 15757 -1520 15763 -1486
rect 15448 -1702 15644 -1694
rect 15448 -1754 15457 -1702
rect 15509 -1754 15521 -1702
rect 15573 -1754 15585 -1702
rect 15637 -1754 15644 -1702
rect 15448 -1764 15644 -1754
rect 15188 -2003 15384 -1995
rect 15188 -2055 15197 -2003
rect 15249 -2055 15261 -2003
rect 15313 -2055 15325 -2003
rect 15377 -2055 15384 -2003
rect 15188 -2065 15384 -2055
rect 15007 -2404 15013 -2370
rect 15047 -2404 15053 -2370
rect 15007 -2442 15053 -2404
rect 15007 -2476 15013 -2442
rect 15047 -2476 15053 -2442
rect 15007 -2523 15053 -2476
rect 15265 -2370 15311 -2065
rect 15265 -2404 15271 -2370
rect 15305 -2404 15311 -2370
rect 15265 -2442 15311 -2404
rect 15265 -2476 15271 -2442
rect 15305 -2476 15311 -2442
rect 15265 -2523 15311 -2476
rect 15523 -2370 15569 -1764
rect 15717 -1834 15763 -1520
rect 15975 -1414 16021 -1367
rect 15975 -1448 15981 -1414
rect 16015 -1448 16021 -1414
rect 15975 -1486 16021 -1448
rect 15975 -1520 15981 -1486
rect 16015 -1520 16021 -1486
rect 15643 -1842 15839 -1834
rect 15643 -1894 15650 -1842
rect 15702 -1894 15714 -1842
rect 15766 -1894 15778 -1842
rect 15830 -1894 15839 -1842
rect 15643 -1904 15839 -1894
rect 15523 -2404 15529 -2370
rect 15563 -2404 15569 -2370
rect 15523 -2442 15569 -2404
rect 15523 -2476 15529 -2442
rect 15563 -2476 15569 -2442
rect 15523 -2523 15569 -2476
rect 15717 -2370 15763 -1904
rect 15975 -2139 16021 -1520
rect 16233 -1414 16279 -1367
rect 16233 -1448 16239 -1414
rect 16273 -1448 16279 -1414
rect 16233 -1486 16279 -1448
rect 16233 -1520 16239 -1486
rect 16273 -1520 16279 -1486
rect 16233 -1834 16279 -1520
rect 16491 -1414 16537 -1367
rect 16491 -1448 16497 -1414
rect 16531 -1448 16537 -1414
rect 16491 -1486 16537 -1448
rect 16491 -1520 16497 -1486
rect 16531 -1520 16537 -1486
rect 16160 -1842 16356 -1834
rect 16160 -1894 16167 -1842
rect 16219 -1894 16231 -1842
rect 16283 -1894 16295 -1842
rect 16347 -1894 16356 -1842
rect 16160 -1904 16356 -1894
rect 15901 -2147 16097 -2139
rect 15901 -2199 15908 -2147
rect 15960 -2199 15972 -2147
rect 16024 -2199 16036 -2147
rect 16088 -2199 16097 -2147
rect 15901 -2209 16097 -2199
rect 15717 -2404 15723 -2370
rect 15757 -2404 15763 -2370
rect 15717 -2442 15763 -2404
rect 15717 -2476 15723 -2442
rect 15757 -2476 15763 -2442
rect 15717 -2523 15763 -2476
rect 15975 -2370 16021 -2209
rect 15975 -2404 15981 -2370
rect 16015 -2404 16021 -2370
rect 15975 -2442 16021 -2404
rect 15975 -2476 15981 -2442
rect 16015 -2476 16021 -2442
rect 15975 -2523 16021 -2476
rect 16233 -2370 16279 -1904
rect 16491 -2139 16537 -1520
rect 16685 -1414 16731 -1367
rect 16685 -1448 16691 -1414
rect 16725 -1448 16731 -1414
rect 16685 -1486 16731 -1448
rect 16685 -1520 16691 -1486
rect 16725 -1520 16731 -1486
rect 16685 -1694 16731 -1520
rect 16943 -1414 16989 -1367
rect 16943 -1448 16949 -1414
rect 16983 -1448 16989 -1414
rect 16943 -1486 16989 -1448
rect 16943 -1520 16949 -1486
rect 16983 -1520 16989 -1486
rect 16608 -1702 16804 -1694
rect 16608 -1754 16617 -1702
rect 16669 -1754 16681 -1702
rect 16733 -1754 16745 -1702
rect 16797 -1754 16804 -1702
rect 16608 -1764 16804 -1754
rect 16418 -2147 16614 -2139
rect 16418 -2199 16425 -2147
rect 16477 -2199 16489 -2147
rect 16541 -2199 16553 -2147
rect 16605 -2199 16614 -2147
rect 16418 -2209 16614 -2199
rect 16233 -2404 16239 -2370
rect 16273 -2404 16279 -2370
rect 16233 -2442 16279 -2404
rect 16233 -2476 16239 -2442
rect 16273 -2476 16279 -2442
rect 16233 -2523 16279 -2476
rect 16491 -2370 16537 -2209
rect 16491 -2404 16497 -2370
rect 16531 -2404 16537 -2370
rect 16491 -2442 16537 -2404
rect 16491 -2476 16497 -2442
rect 16531 -2476 16537 -2442
rect 16491 -2523 16537 -2476
rect 16685 -2370 16731 -1764
rect 16943 -1995 16989 -1520
rect 17201 -1414 17247 -1367
rect 17201 -1448 17207 -1414
rect 17241 -1448 17247 -1414
rect 17201 -1486 17247 -1448
rect 17201 -1520 17207 -1486
rect 17241 -1520 17247 -1486
rect 17201 -1694 17247 -1520
rect 17459 -1414 17505 -1367
rect 17459 -1448 17465 -1414
rect 17499 -1448 17505 -1414
rect 17459 -1486 17505 -1448
rect 17459 -1520 17465 -1486
rect 17499 -1520 17505 -1486
rect 17126 -1702 17322 -1694
rect 17126 -1754 17135 -1702
rect 17187 -1754 17199 -1702
rect 17251 -1754 17263 -1702
rect 17315 -1754 17322 -1702
rect 17126 -1764 17322 -1754
rect 16865 -2003 17061 -1995
rect 16865 -2055 16874 -2003
rect 16926 -2055 16938 -2003
rect 16990 -2055 17002 -2003
rect 17054 -2055 17061 -2003
rect 16865 -2065 17061 -2055
rect 16685 -2404 16691 -2370
rect 16725 -2404 16731 -2370
rect 16685 -2442 16731 -2404
rect 16685 -2476 16691 -2442
rect 16725 -2476 16731 -2442
rect 16685 -2523 16731 -2476
rect 16943 -2370 16989 -2065
rect 16943 -2404 16949 -2370
rect 16983 -2404 16989 -2370
rect 16943 -2442 16989 -2404
rect 16943 -2476 16949 -2442
rect 16983 -2476 16989 -2442
rect 16943 -2523 16989 -2476
rect 17201 -2370 17247 -1764
rect 17459 -1995 17505 -1520
rect 17717 -1414 17763 -1367
rect 17717 -1448 17723 -1414
rect 17757 -1448 17763 -1414
rect 17717 -1486 17763 -1448
rect 17717 -1520 17723 -1486
rect 17757 -1520 17763 -1486
rect 17717 -1694 17763 -1520
rect 17911 -1384 18290 -1350
rect 18324 -1384 18347 -1350
rect 17911 -1414 18347 -1384
rect 17911 -1448 17917 -1414
rect 17951 -1448 18175 -1414
rect 18209 -1422 18347 -1414
rect 18209 -1448 18290 -1422
rect 17911 -1456 18290 -1448
rect 18324 -1456 18347 -1422
rect 17911 -1486 18347 -1456
rect 17911 -1520 17917 -1486
rect 17951 -1520 18175 -1486
rect 18209 -1494 18347 -1486
rect 18209 -1520 18290 -1494
rect 17911 -1528 18290 -1520
rect 18324 -1528 18347 -1494
rect 17911 -1566 18347 -1528
rect 17911 -1600 18290 -1566
rect 18324 -1600 18347 -1566
rect 17911 -1638 18347 -1600
rect 17911 -1672 18290 -1638
rect 18324 -1672 18347 -1638
rect 17641 -1702 17837 -1694
rect 17641 -1754 17650 -1702
rect 17702 -1754 17714 -1702
rect 17766 -1754 17778 -1702
rect 17830 -1754 17837 -1702
rect 17641 -1764 17837 -1754
rect 17911 -1710 18347 -1672
rect 17911 -1744 18290 -1710
rect 18324 -1744 18347 -1710
rect 17383 -2003 17579 -1995
rect 17383 -2055 17392 -2003
rect 17444 -2055 17456 -2003
rect 17508 -2055 17520 -2003
rect 17572 -2055 17579 -2003
rect 17383 -2065 17579 -2055
rect 17201 -2404 17207 -2370
rect 17241 -2404 17247 -2370
rect 17201 -2442 17247 -2404
rect 17201 -2476 17207 -2442
rect 17241 -2476 17247 -2442
rect 17201 -2523 17247 -2476
rect 17459 -2370 17505 -2065
rect 17459 -2404 17465 -2370
rect 17499 -2404 17505 -2370
rect 17459 -2442 17505 -2404
rect 17459 -2476 17465 -2442
rect 17499 -2476 17505 -2442
rect 17459 -2523 17505 -2476
rect 17717 -2370 17763 -1764
rect 17717 -2404 17723 -2370
rect 17757 -2404 17763 -2370
rect 17717 -2442 17763 -2404
rect 17717 -2476 17723 -2442
rect 17757 -2476 17763 -2442
rect 17717 -2523 17763 -2476
rect 17911 -1782 18347 -1744
rect 17911 -1816 18290 -1782
rect 18324 -1816 18347 -1782
rect 17911 -1854 18347 -1816
rect 17911 -1888 18290 -1854
rect 18324 -1888 18347 -1854
rect 17911 -1926 18347 -1888
rect 17911 -1960 18290 -1926
rect 18324 -1960 18347 -1926
rect 17911 -1998 18347 -1960
rect 17911 -2032 18290 -1998
rect 18324 -2032 18347 -1998
rect 17911 -2070 18347 -2032
rect 17911 -2104 18290 -2070
rect 18324 -2104 18347 -2070
rect 17911 -2142 18347 -2104
rect 17911 -2176 18290 -2142
rect 18324 -2176 18347 -2142
rect 17911 -2214 18347 -2176
rect 17911 -2248 18290 -2214
rect 18324 -2248 18347 -2214
rect 17911 -2286 18347 -2248
rect 17911 -2320 18290 -2286
rect 18324 -2320 18347 -2286
rect 17911 -2358 18347 -2320
rect 17911 -2370 18290 -2358
rect 17911 -2404 17917 -2370
rect 17951 -2404 18175 -2370
rect 18209 -2392 18290 -2370
rect 18324 -2392 18347 -2358
rect 18209 -2404 18347 -2392
rect 17911 -2430 18347 -2404
rect 17911 -2442 18290 -2430
rect 17911 -2476 17917 -2442
rect 17951 -2476 18175 -2442
rect 18209 -2464 18290 -2442
rect 18324 -2464 18347 -2430
rect 18209 -2476 18347 -2464
rect 17911 -2502 18347 -2476
rect 9194 -2604 9293 -2570
rect 9327 -2604 9365 -2570
rect 9399 -2574 9781 -2570
rect 9399 -2604 9573 -2574
rect 9194 -2608 9573 -2604
rect 9607 -2604 9781 -2574
rect 9815 -2604 9853 -2570
rect 9887 -2604 9986 -2570
rect 9607 -2608 9986 -2604
rect 9194 -2646 9986 -2608
rect 7886 -2885 7947 -2653
rect 9194 -2680 9573 -2646
rect 9607 -2680 9986 -2646
rect 10190 -2570 11294 -2564
rect 10190 -2604 10233 -2570
rect 10267 -2583 10305 -2570
rect 10339 -2583 10491 -2570
rect 10525 -2583 10563 -2570
rect 10597 -2583 10749 -2570
rect 10783 -2583 10821 -2570
rect 10855 -2583 11007 -2570
rect 11041 -2583 11079 -2570
rect 10190 -2635 10240 -2604
rect 10292 -2635 10304 -2583
rect 10356 -2635 10368 -2583
rect 10420 -2635 10436 -2583
rect 10488 -2604 10491 -2583
rect 10552 -2604 10563 -2583
rect 10488 -2635 10500 -2604
rect 10552 -2635 10564 -2604
rect 10616 -2635 10726 -2583
rect 10783 -2604 10790 -2583
rect 10778 -2635 10790 -2604
rect 10842 -2635 10854 -2604
rect 10906 -2635 10922 -2583
rect 10974 -2635 10986 -2583
rect 11041 -2604 11050 -2583
rect 11113 -2604 11294 -2570
rect 11038 -2635 11050 -2604
rect 11102 -2635 11294 -2604
rect 10190 -2653 11294 -2635
rect 6873 -2933 7947 -2885
rect 6873 -2967 7099 -2933
rect 7133 -2967 7171 -2933
rect 7205 -2967 7357 -2933
rect 7391 -2967 7429 -2933
rect 7463 -2967 7615 -2933
rect 7649 -2967 7687 -2933
rect 7721 -2967 7947 -2933
rect 6873 -2973 7947 -2967
rect 8024 -2721 8990 -2703
rect 8024 -2773 8078 -2721
rect 8130 -2773 8142 -2721
rect 8194 -2773 8206 -2721
rect 8258 -2773 8274 -2721
rect 8326 -2773 8338 -2721
rect 8390 -2773 8402 -2721
rect 8454 -2773 8564 -2721
rect 8616 -2773 8628 -2721
rect 8680 -2773 8692 -2721
rect 8744 -2773 8760 -2721
rect 8812 -2773 8824 -2721
rect 8876 -2773 8888 -2721
rect 8940 -2773 8990 -2721
rect 8024 -2899 8990 -2773
rect 8024 -2933 8078 -2899
rect 8130 -2933 8142 -2899
rect 8024 -2967 8067 -2933
rect 8130 -2951 8139 -2933
rect 8194 -2951 8206 -2899
rect 8258 -2951 8274 -2899
rect 8326 -2933 8338 -2899
rect 8390 -2933 8402 -2899
rect 8390 -2951 8397 -2933
rect 8454 -2951 8564 -2899
rect 8616 -2933 8628 -2899
rect 8680 -2933 8692 -2899
rect 8617 -2951 8628 -2933
rect 8689 -2951 8692 -2933
rect 8744 -2951 8760 -2899
rect 8812 -2951 8824 -2899
rect 8876 -2951 8888 -2899
rect 8940 -2933 8990 -2899
rect 8101 -2967 8139 -2951
rect 8173 -2967 8325 -2951
rect 8359 -2967 8397 -2951
rect 8431 -2967 8583 -2951
rect 8617 -2967 8655 -2951
rect 8689 -2967 8841 -2951
rect 8875 -2967 8913 -2951
rect 8947 -2967 8990 -2933
rect 8024 -2973 8990 -2967
rect 9194 -2718 9986 -2680
rect 9194 -2752 9573 -2718
rect 9607 -2752 9986 -2718
rect 9194 -2790 9986 -2752
rect 9194 -2824 9573 -2790
rect 9607 -2824 9986 -2790
rect 9194 -2862 9986 -2824
rect 9194 -2896 9573 -2862
rect 9607 -2896 9986 -2862
rect 9194 -2933 9986 -2896
rect 9194 -2967 9293 -2933
rect 9327 -2967 9365 -2933
rect 9399 -2934 9781 -2933
rect 9399 -2967 9573 -2934
rect 9194 -2968 9573 -2967
rect 9607 -2967 9781 -2934
rect 9815 -2967 9853 -2933
rect 9887 -2967 9986 -2933
rect 9607 -2968 9986 -2967
rect 833 -3061 1269 -3040
rect 833 -3078 971 -3061
rect 833 -3112 856 -3078
rect 890 -3095 971 -3078
rect 1005 -3095 1229 -3061
rect 1263 -3095 1269 -3061
rect 890 -3112 1269 -3095
rect 833 -3133 1269 -3112
rect 833 -3150 971 -3133
rect 833 -3184 856 -3150
rect 890 -3167 971 -3150
rect 1005 -3167 1229 -3133
rect 1263 -3167 1269 -3133
rect 890 -3184 1269 -3167
rect 833 -3222 1269 -3184
rect 833 -3256 856 -3222
rect 890 -3256 1269 -3222
rect 833 -3294 1269 -3256
rect 833 -3328 856 -3294
rect 890 -3328 1269 -3294
rect 833 -3366 1269 -3328
rect 833 -3400 856 -3366
rect 890 -3400 1269 -3366
rect 833 -3438 1269 -3400
rect 833 -3472 856 -3438
rect 890 -3472 1269 -3438
rect 833 -3510 1269 -3472
rect 833 -3544 856 -3510
rect 890 -3544 1269 -3510
rect 833 -3582 1269 -3544
rect 833 -3616 856 -3582
rect 890 -3616 1269 -3582
rect 833 -3654 1269 -3616
rect 1417 -3061 1463 -3014
rect 1417 -3095 1423 -3061
rect 1457 -3095 1463 -3061
rect 1417 -3133 1463 -3095
rect 1417 -3167 1423 -3133
rect 1457 -3167 1463 -3133
rect 1417 -3647 1463 -3167
rect 1675 -3061 1721 -3014
rect 1675 -3095 1681 -3061
rect 1715 -3095 1721 -3061
rect 1675 -3133 1721 -3095
rect 1675 -3167 1681 -3133
rect 1715 -3167 1721 -3133
rect 1675 -3316 1721 -3167
rect 1933 -3061 1979 -3014
rect 1933 -3095 1939 -3061
rect 1973 -3095 1979 -3061
rect 1933 -3133 1979 -3095
rect 1933 -3167 1939 -3133
rect 1973 -3167 1979 -3133
rect 1598 -3326 1794 -3316
rect 1598 -3378 1607 -3326
rect 1659 -3378 1671 -3326
rect 1723 -3378 1735 -3326
rect 1787 -3378 1794 -3326
rect 1598 -3386 1794 -3378
rect 1933 -3647 1979 -3167
rect 2191 -3061 2237 -3014
rect 2191 -3095 2197 -3061
rect 2231 -3095 2237 -3061
rect 2191 -3133 2237 -3095
rect 2191 -3167 2197 -3133
rect 2231 -3167 2237 -3133
rect 2191 -3316 2237 -3167
rect 2449 -3061 2495 -3014
rect 2449 -3095 2455 -3061
rect 2489 -3095 2495 -3061
rect 2449 -3133 2495 -3095
rect 2449 -3167 2455 -3133
rect 2489 -3167 2495 -3133
rect 2116 -3326 2312 -3316
rect 2116 -3378 2125 -3326
rect 2177 -3378 2189 -3326
rect 2241 -3378 2253 -3326
rect 2305 -3378 2312 -3326
rect 2116 -3386 2312 -3378
rect 2449 -3647 2495 -3167
rect 2643 -3061 2689 -3014
rect 2643 -3095 2649 -3061
rect 2683 -3095 2689 -3061
rect 2643 -3133 2689 -3095
rect 2643 -3167 2649 -3133
rect 2683 -3167 2689 -3133
rect 2643 -3485 2689 -3167
rect 2901 -3061 2947 -3014
rect 2901 -3095 2907 -3061
rect 2941 -3095 2947 -3061
rect 2901 -3133 2947 -3095
rect 2901 -3167 2907 -3133
rect 2941 -3167 2947 -3133
rect 2570 -3495 2766 -3485
rect 2570 -3547 2577 -3495
rect 2629 -3547 2641 -3495
rect 2693 -3547 2705 -3495
rect 2757 -3547 2766 -3495
rect 2570 -3555 2766 -3547
rect 833 -3688 856 -3654
rect 890 -3688 1269 -3654
rect 833 -3726 1269 -3688
rect 1339 -3657 1535 -3647
rect 1339 -3709 1348 -3657
rect 1400 -3709 1412 -3657
rect 1464 -3709 1476 -3657
rect 1528 -3709 1535 -3657
rect 1339 -3717 1535 -3709
rect 1856 -3657 2052 -3647
rect 1856 -3709 1865 -3657
rect 1917 -3709 1929 -3657
rect 1981 -3709 1993 -3657
rect 2045 -3709 2052 -3657
rect 1856 -3717 2052 -3709
rect 2373 -3657 2569 -3647
rect 2373 -3709 2382 -3657
rect 2434 -3709 2446 -3657
rect 2498 -3709 2510 -3657
rect 2562 -3709 2569 -3657
rect 2373 -3717 2569 -3709
rect 833 -3760 856 -3726
rect 890 -3760 1269 -3726
rect 833 -3798 1269 -3760
rect 833 -3832 856 -3798
rect 890 -3832 1269 -3798
rect 2901 -3816 2947 -3167
rect 3159 -3061 3205 -3014
rect 3159 -3095 3165 -3061
rect 3199 -3095 3205 -3061
rect 3159 -3133 3205 -3095
rect 3159 -3167 3165 -3133
rect 3199 -3167 3205 -3133
rect 3159 -3485 3205 -3167
rect 3417 -3061 3463 -3014
rect 3417 -3095 3423 -3061
rect 3457 -3095 3463 -3061
rect 3417 -3133 3463 -3095
rect 3417 -3167 3423 -3133
rect 3457 -3167 3463 -3133
rect 3087 -3495 3283 -3485
rect 3087 -3547 3094 -3495
rect 3146 -3547 3158 -3495
rect 3210 -3547 3222 -3495
rect 3274 -3547 3283 -3495
rect 3087 -3555 3283 -3547
rect 3417 -3816 3463 -3167
rect 3611 -3061 3657 -3014
rect 3611 -3095 3617 -3061
rect 3651 -3095 3657 -3061
rect 3611 -3133 3657 -3095
rect 3611 -3167 3617 -3133
rect 3651 -3167 3657 -3133
rect 3611 -3647 3657 -3167
rect 3869 -3061 3915 -3014
rect 3869 -3095 3875 -3061
rect 3909 -3095 3915 -3061
rect 3869 -3133 3915 -3095
rect 3869 -3167 3875 -3133
rect 3909 -3167 3915 -3133
rect 3869 -3316 3915 -3167
rect 4127 -3061 4173 -3014
rect 4127 -3095 4133 -3061
rect 4167 -3095 4173 -3061
rect 4127 -3133 4173 -3095
rect 4127 -3167 4133 -3133
rect 4167 -3167 4173 -3133
rect 3793 -3326 3989 -3316
rect 3793 -3378 3802 -3326
rect 3854 -3378 3866 -3326
rect 3918 -3378 3930 -3326
rect 3982 -3378 3989 -3326
rect 3793 -3386 3989 -3378
rect 4127 -3647 4173 -3167
rect 4385 -3061 4431 -3014
rect 4385 -3095 4391 -3061
rect 4425 -3095 4431 -3061
rect 4385 -3133 4431 -3095
rect 4385 -3167 4391 -3133
rect 4425 -3167 4431 -3133
rect 4385 -3316 4431 -3167
rect 4643 -3061 4689 -3014
rect 4643 -3095 4649 -3061
rect 4683 -3095 4689 -3061
rect 4643 -3133 4689 -3095
rect 4643 -3167 4649 -3133
rect 4683 -3167 4689 -3133
rect 4310 -3326 4506 -3316
rect 4310 -3378 4319 -3326
rect 4371 -3378 4383 -3326
rect 4435 -3378 4447 -3326
rect 4499 -3378 4506 -3326
rect 4310 -3386 4506 -3378
rect 4643 -3647 4689 -3167
rect 4836 -3040 5214 -3006
rect 5248 -3040 5626 -3006
rect 9194 -3006 9986 -2968
rect 10190 -2721 11156 -2703
rect 10190 -2773 10240 -2721
rect 10292 -2773 10304 -2721
rect 10356 -2773 10368 -2721
rect 10420 -2773 10436 -2721
rect 10488 -2773 10500 -2721
rect 10552 -2773 10564 -2721
rect 10616 -2773 10726 -2721
rect 10778 -2773 10790 -2721
rect 10842 -2773 10854 -2721
rect 10906 -2773 10922 -2721
rect 10974 -2773 10986 -2721
rect 11038 -2773 11050 -2721
rect 11102 -2773 11156 -2721
rect 10190 -2899 11156 -2773
rect 10190 -2933 10240 -2899
rect 10190 -2967 10233 -2933
rect 10292 -2951 10304 -2899
rect 10356 -2951 10368 -2899
rect 10420 -2951 10436 -2899
rect 10488 -2933 10500 -2899
rect 10552 -2933 10564 -2899
rect 10488 -2951 10491 -2933
rect 10552 -2951 10563 -2933
rect 10616 -2951 10726 -2899
rect 10778 -2933 10790 -2899
rect 10842 -2933 10854 -2899
rect 10783 -2951 10790 -2933
rect 10906 -2951 10922 -2899
rect 10974 -2951 10986 -2899
rect 11038 -2933 11050 -2899
rect 11102 -2933 11156 -2899
rect 11041 -2951 11050 -2933
rect 10267 -2967 10305 -2951
rect 10339 -2967 10491 -2951
rect 10525 -2967 10563 -2951
rect 10597 -2967 10749 -2951
rect 10783 -2967 10821 -2951
rect 10855 -2967 11007 -2951
rect 11041 -2967 11079 -2951
rect 11113 -2967 11156 -2933
rect 10190 -2973 11156 -2967
rect 11233 -2885 11294 -2653
rect 11416 -2570 12124 -2564
rect 11416 -2604 11459 -2570
rect 11493 -2604 11531 -2570
rect 11565 -2604 11717 -2570
rect 11751 -2604 11789 -2570
rect 11823 -2604 11975 -2570
rect 12009 -2604 12047 -2570
rect 12081 -2604 12124 -2570
rect 11416 -2721 12124 -2604
rect 11416 -2773 11450 -2721
rect 11502 -2773 11514 -2721
rect 11566 -2773 11578 -2721
rect 11630 -2773 11646 -2721
rect 11698 -2773 11710 -2721
rect 11762 -2773 11774 -2721
rect 11826 -2773 11838 -2721
rect 11890 -2773 11906 -2721
rect 11958 -2773 11970 -2721
rect 12022 -2773 12034 -2721
rect 12086 -2773 12124 -2721
rect 11416 -2791 12124 -2773
rect 12246 -2570 13350 -2564
rect 12246 -2604 12427 -2570
rect 12461 -2583 12499 -2570
rect 12533 -2583 12685 -2570
rect 12719 -2583 12757 -2570
rect 12791 -2583 12943 -2570
rect 12977 -2583 13015 -2570
rect 13049 -2583 13201 -2570
rect 13235 -2583 13273 -2570
rect 12490 -2604 12499 -2583
rect 12246 -2635 12438 -2604
rect 12490 -2635 12502 -2604
rect 12554 -2635 12566 -2583
rect 12618 -2635 12634 -2583
rect 12750 -2604 12757 -2583
rect 12686 -2635 12698 -2604
rect 12750 -2635 12762 -2604
rect 12814 -2635 12924 -2583
rect 12977 -2604 12988 -2583
rect 13049 -2604 13052 -2583
rect 12976 -2635 12988 -2604
rect 13040 -2635 13052 -2604
rect 13104 -2635 13120 -2583
rect 13172 -2635 13184 -2583
rect 13236 -2635 13248 -2583
rect 13307 -2604 13350 -2570
rect 13300 -2635 13350 -2604
rect 12246 -2653 13350 -2635
rect 13554 -2570 14344 -2536
rect 17911 -2536 18290 -2502
rect 18324 -2536 18347 -2502
rect 13554 -2604 13653 -2570
rect 13687 -2604 13725 -2570
rect 13759 -2574 14139 -2570
rect 13759 -2604 13932 -2574
rect 13554 -2608 13932 -2604
rect 13966 -2604 14139 -2574
rect 14173 -2604 14211 -2570
rect 14245 -2604 14344 -2570
rect 13966 -2608 14344 -2604
rect 13554 -2646 14344 -2608
rect 12246 -2885 12307 -2653
rect 13554 -2680 13932 -2646
rect 13966 -2680 14344 -2646
rect 14547 -2570 15651 -2564
rect 14547 -2604 14590 -2570
rect 14624 -2583 14662 -2570
rect 14696 -2583 14848 -2570
rect 14882 -2583 14920 -2570
rect 14954 -2583 15106 -2570
rect 15140 -2583 15178 -2570
rect 15212 -2583 15364 -2570
rect 15398 -2583 15436 -2570
rect 14547 -2635 14597 -2604
rect 14649 -2635 14661 -2583
rect 14713 -2635 14725 -2583
rect 14777 -2635 14793 -2583
rect 14845 -2604 14848 -2583
rect 14909 -2604 14920 -2583
rect 14845 -2635 14857 -2604
rect 14909 -2635 14921 -2604
rect 14973 -2635 15083 -2583
rect 15140 -2604 15147 -2583
rect 15135 -2635 15147 -2604
rect 15199 -2635 15211 -2604
rect 15263 -2635 15279 -2583
rect 15331 -2635 15343 -2583
rect 15398 -2604 15407 -2583
rect 15470 -2604 15651 -2570
rect 15395 -2635 15407 -2604
rect 15459 -2635 15651 -2604
rect 14547 -2653 15651 -2635
rect 11233 -2933 12307 -2885
rect 11233 -2967 11459 -2933
rect 11493 -2967 11531 -2933
rect 11565 -2967 11717 -2933
rect 11751 -2967 11789 -2933
rect 11823 -2967 11975 -2933
rect 12009 -2967 12047 -2933
rect 12081 -2967 12307 -2933
rect 11233 -2973 12307 -2967
rect 12384 -2721 13350 -2703
rect 12384 -2773 12438 -2721
rect 12490 -2773 12502 -2721
rect 12554 -2773 12566 -2721
rect 12618 -2773 12634 -2721
rect 12686 -2773 12698 -2721
rect 12750 -2773 12762 -2721
rect 12814 -2773 12924 -2721
rect 12976 -2773 12988 -2721
rect 13040 -2773 13052 -2721
rect 13104 -2773 13120 -2721
rect 13172 -2773 13184 -2721
rect 13236 -2773 13248 -2721
rect 13300 -2773 13350 -2721
rect 12384 -2899 13350 -2773
rect 12384 -2933 12438 -2899
rect 12490 -2933 12502 -2899
rect 12384 -2967 12427 -2933
rect 12490 -2951 12499 -2933
rect 12554 -2951 12566 -2899
rect 12618 -2951 12634 -2899
rect 12686 -2933 12698 -2899
rect 12750 -2933 12762 -2899
rect 12750 -2951 12757 -2933
rect 12814 -2951 12924 -2899
rect 12976 -2933 12988 -2899
rect 13040 -2933 13052 -2899
rect 12977 -2951 12988 -2933
rect 13049 -2951 13052 -2933
rect 13104 -2951 13120 -2899
rect 13172 -2951 13184 -2899
rect 13236 -2951 13248 -2899
rect 13300 -2933 13350 -2899
rect 12461 -2967 12499 -2951
rect 12533 -2967 12685 -2951
rect 12719 -2967 12757 -2951
rect 12791 -2967 12943 -2951
rect 12977 -2967 13015 -2951
rect 13049 -2967 13201 -2951
rect 13235 -2967 13273 -2951
rect 13307 -2967 13350 -2933
rect 12384 -2973 13350 -2967
rect 13554 -2718 14344 -2680
rect 13554 -2752 13932 -2718
rect 13966 -2752 14344 -2718
rect 13554 -2790 14344 -2752
rect 13554 -2824 13932 -2790
rect 13966 -2824 14344 -2790
rect 13554 -2862 14344 -2824
rect 13554 -2896 13932 -2862
rect 13966 -2896 14344 -2862
rect 13554 -2933 14344 -2896
rect 13554 -2967 13653 -2933
rect 13687 -2967 13725 -2933
rect 13759 -2934 14139 -2933
rect 13759 -2967 13932 -2934
rect 13554 -2968 13932 -2967
rect 13966 -2967 14139 -2934
rect 14173 -2967 14211 -2933
rect 14245 -2967 14344 -2933
rect 13966 -2968 14344 -2967
rect 4836 -3061 5626 -3040
rect 4836 -3095 4842 -3061
rect 4876 -3095 5100 -3061
rect 5134 -3078 5328 -3061
rect 5134 -3095 5214 -3078
rect 4836 -3112 5214 -3095
rect 5248 -3095 5328 -3078
rect 5362 -3095 5586 -3061
rect 5620 -3095 5626 -3061
rect 5248 -3112 5626 -3095
rect 4836 -3133 5626 -3112
rect 4836 -3167 4842 -3133
rect 4876 -3167 5100 -3133
rect 5134 -3150 5328 -3133
rect 5134 -3167 5214 -3150
rect 4836 -3184 5214 -3167
rect 5248 -3167 5328 -3150
rect 5362 -3167 5586 -3133
rect 5620 -3167 5626 -3133
rect 5248 -3184 5626 -3167
rect 4836 -3222 5626 -3184
rect 4836 -3256 5214 -3222
rect 5248 -3256 5626 -3222
rect 4836 -3294 5626 -3256
rect 4836 -3328 5214 -3294
rect 5248 -3328 5626 -3294
rect 4836 -3366 5626 -3328
rect 4836 -3400 5214 -3366
rect 5248 -3400 5626 -3366
rect 4836 -3438 5626 -3400
rect 4836 -3472 5214 -3438
rect 5248 -3472 5626 -3438
rect 4836 -3510 5626 -3472
rect 4836 -3544 5214 -3510
rect 5248 -3544 5626 -3510
rect 4836 -3582 5626 -3544
rect 4836 -3616 5214 -3582
rect 5248 -3616 5626 -3582
rect 3534 -3657 3730 -3647
rect 3534 -3709 3543 -3657
rect 3595 -3709 3607 -3657
rect 3659 -3709 3671 -3657
rect 3723 -3709 3730 -3657
rect 3534 -3717 3730 -3709
rect 4051 -3657 4247 -3647
rect 4051 -3709 4060 -3657
rect 4112 -3709 4124 -3657
rect 4176 -3709 4188 -3657
rect 4240 -3709 4247 -3657
rect 4051 -3717 4247 -3709
rect 4566 -3657 4762 -3647
rect 4566 -3709 4575 -3657
rect 4627 -3709 4639 -3657
rect 4691 -3709 4703 -3657
rect 4755 -3709 4762 -3657
rect 4566 -3717 4762 -3709
rect 4836 -3654 5626 -3616
rect 5774 -3061 5820 -3014
rect 5774 -3095 5780 -3061
rect 5814 -3095 5820 -3061
rect 5774 -3133 5820 -3095
rect 5774 -3167 5780 -3133
rect 5814 -3167 5820 -3133
rect 5774 -3647 5820 -3167
rect 6032 -3061 6078 -3014
rect 6032 -3095 6038 -3061
rect 6072 -3095 6078 -3061
rect 6032 -3133 6078 -3095
rect 6032 -3167 6038 -3133
rect 6072 -3167 6078 -3133
rect 6032 -3316 6078 -3167
rect 6290 -3061 6336 -3014
rect 6290 -3095 6296 -3061
rect 6330 -3095 6336 -3061
rect 6290 -3133 6336 -3095
rect 6290 -3167 6296 -3133
rect 6330 -3167 6336 -3133
rect 5957 -3326 6153 -3316
rect 5957 -3378 5964 -3326
rect 6016 -3378 6028 -3326
rect 6080 -3378 6092 -3326
rect 6144 -3378 6153 -3326
rect 5957 -3386 6153 -3378
rect 6290 -3647 6336 -3167
rect 6548 -3061 6594 -3014
rect 6548 -3095 6554 -3061
rect 6588 -3095 6594 -3061
rect 6548 -3133 6594 -3095
rect 6548 -3167 6554 -3133
rect 6588 -3167 6594 -3133
rect 6548 -3316 6594 -3167
rect 6806 -3061 6852 -3014
rect 6806 -3095 6812 -3061
rect 6846 -3095 6852 -3061
rect 6806 -3133 6852 -3095
rect 6806 -3167 6812 -3133
rect 6846 -3167 6852 -3133
rect 6474 -3326 6670 -3316
rect 6474 -3378 6481 -3326
rect 6533 -3378 6545 -3326
rect 6597 -3378 6609 -3326
rect 6661 -3378 6670 -3326
rect 6474 -3386 6670 -3378
rect 6806 -3647 6852 -3167
rect 7000 -3061 7046 -3014
rect 7000 -3095 7006 -3061
rect 7040 -3095 7046 -3061
rect 7000 -3133 7046 -3095
rect 7000 -3167 7006 -3133
rect 7040 -3167 7046 -3133
rect 4836 -3688 5214 -3654
rect 5248 -3688 5626 -3654
rect 4836 -3726 5626 -3688
rect 5701 -3657 5897 -3647
rect 5701 -3709 5708 -3657
rect 5760 -3709 5772 -3657
rect 5824 -3709 5836 -3657
rect 5888 -3709 5897 -3657
rect 5701 -3717 5897 -3709
rect 6216 -3657 6412 -3647
rect 6216 -3709 6223 -3657
rect 6275 -3709 6287 -3657
rect 6339 -3709 6351 -3657
rect 6403 -3709 6412 -3657
rect 6216 -3717 6412 -3709
rect 6733 -3657 6929 -3647
rect 6733 -3709 6740 -3657
rect 6792 -3709 6804 -3657
rect 6856 -3709 6868 -3657
rect 6920 -3709 6929 -3657
rect 6733 -3717 6929 -3709
rect 4836 -3760 5214 -3726
rect 5248 -3760 5626 -3726
rect 4836 -3798 5626 -3760
rect 833 -3870 1269 -3832
rect 833 -3904 856 -3870
rect 890 -3904 1269 -3870
rect 2827 -3826 3023 -3816
rect 2827 -3878 2834 -3826
rect 2886 -3878 2898 -3826
rect 2950 -3878 2962 -3826
rect 3014 -3878 3023 -3826
rect 2827 -3886 3023 -3878
rect 3344 -3826 3540 -3816
rect 3344 -3878 3351 -3826
rect 3403 -3878 3415 -3826
rect 3467 -3878 3479 -3826
rect 3531 -3878 3540 -3826
rect 3344 -3886 3540 -3878
rect 4836 -3832 5214 -3798
rect 5248 -3832 5626 -3798
rect 7000 -3816 7046 -3167
rect 7258 -3061 7304 -3014
rect 7258 -3095 7264 -3061
rect 7298 -3095 7304 -3061
rect 7258 -3133 7304 -3095
rect 7258 -3167 7264 -3133
rect 7298 -3167 7304 -3133
rect 7258 -3485 7304 -3167
rect 7516 -3061 7562 -3014
rect 7516 -3095 7522 -3061
rect 7556 -3095 7562 -3061
rect 7516 -3133 7562 -3095
rect 7516 -3167 7522 -3133
rect 7556 -3167 7562 -3133
rect 7180 -3495 7376 -3485
rect 7180 -3547 7189 -3495
rect 7241 -3547 7253 -3495
rect 7305 -3547 7317 -3495
rect 7369 -3547 7376 -3495
rect 7180 -3555 7376 -3547
rect 7516 -3816 7562 -3167
rect 7774 -3061 7820 -3014
rect 7774 -3095 7780 -3061
rect 7814 -3095 7820 -3061
rect 7774 -3133 7820 -3095
rect 7774 -3167 7780 -3133
rect 7814 -3167 7820 -3133
rect 7774 -3485 7820 -3167
rect 7968 -3061 8014 -3014
rect 7968 -3095 7974 -3061
rect 8008 -3095 8014 -3061
rect 7968 -3133 8014 -3095
rect 7968 -3167 7974 -3133
rect 8008 -3167 8014 -3133
rect 7697 -3495 7893 -3485
rect 7697 -3547 7706 -3495
rect 7758 -3547 7770 -3495
rect 7822 -3547 7834 -3495
rect 7886 -3547 7893 -3495
rect 7697 -3555 7893 -3547
rect 7968 -3647 8014 -3167
rect 8226 -3061 8272 -3014
rect 8226 -3095 8232 -3061
rect 8266 -3095 8272 -3061
rect 8226 -3133 8272 -3095
rect 8226 -3167 8232 -3133
rect 8266 -3167 8272 -3133
rect 8226 -3316 8272 -3167
rect 8484 -3061 8530 -3014
rect 8484 -3095 8490 -3061
rect 8524 -3095 8530 -3061
rect 8484 -3133 8530 -3095
rect 8484 -3167 8490 -3133
rect 8524 -3167 8530 -3133
rect 8151 -3326 8347 -3316
rect 8151 -3378 8158 -3326
rect 8210 -3378 8222 -3326
rect 8274 -3378 8286 -3326
rect 8338 -3378 8347 -3326
rect 8151 -3386 8347 -3378
rect 8484 -3647 8530 -3167
rect 8742 -3061 8788 -3014
rect 8742 -3095 8748 -3061
rect 8782 -3095 8788 -3061
rect 8742 -3133 8788 -3095
rect 8742 -3167 8748 -3133
rect 8782 -3167 8788 -3133
rect 8742 -3316 8788 -3167
rect 9000 -3061 9046 -3014
rect 9000 -3095 9006 -3061
rect 9040 -3095 9046 -3061
rect 9000 -3133 9046 -3095
rect 9000 -3167 9006 -3133
rect 9040 -3167 9046 -3133
rect 8668 -3326 8864 -3316
rect 8668 -3378 8675 -3326
rect 8727 -3378 8739 -3326
rect 8791 -3378 8803 -3326
rect 8855 -3378 8864 -3326
rect 8668 -3386 8864 -3378
rect 9000 -3647 9046 -3167
rect 9194 -3040 9573 -3006
rect 9607 -3040 9986 -3006
rect 13554 -3006 14344 -2968
rect 14547 -2721 15513 -2703
rect 14547 -2773 14597 -2721
rect 14649 -2773 14661 -2721
rect 14713 -2773 14725 -2721
rect 14777 -2773 14793 -2721
rect 14845 -2773 14857 -2721
rect 14909 -2773 14921 -2721
rect 14973 -2773 15083 -2721
rect 15135 -2773 15147 -2721
rect 15199 -2773 15211 -2721
rect 15263 -2773 15279 -2721
rect 15331 -2773 15343 -2721
rect 15395 -2773 15407 -2721
rect 15459 -2773 15513 -2721
rect 14547 -2899 15513 -2773
rect 14547 -2933 14597 -2899
rect 14547 -2967 14590 -2933
rect 14649 -2951 14661 -2899
rect 14713 -2951 14725 -2899
rect 14777 -2951 14793 -2899
rect 14845 -2933 14857 -2899
rect 14909 -2933 14921 -2899
rect 14845 -2951 14848 -2933
rect 14909 -2951 14920 -2933
rect 14973 -2951 15083 -2899
rect 15135 -2933 15147 -2899
rect 15199 -2933 15211 -2899
rect 15140 -2951 15147 -2933
rect 15263 -2951 15279 -2899
rect 15331 -2951 15343 -2899
rect 15395 -2933 15407 -2899
rect 15459 -2933 15513 -2899
rect 15398 -2951 15407 -2933
rect 14624 -2967 14662 -2951
rect 14696 -2967 14848 -2951
rect 14882 -2967 14920 -2951
rect 14954 -2967 15106 -2951
rect 15140 -2967 15178 -2951
rect 15212 -2967 15364 -2951
rect 15398 -2967 15436 -2951
rect 15470 -2967 15513 -2933
rect 14547 -2973 15513 -2967
rect 15590 -2885 15651 -2653
rect 15773 -2570 16481 -2564
rect 15773 -2604 15816 -2570
rect 15850 -2604 15888 -2570
rect 15922 -2604 16074 -2570
rect 16108 -2604 16146 -2570
rect 16180 -2604 16332 -2570
rect 16366 -2604 16404 -2570
rect 16438 -2604 16481 -2570
rect 15773 -2721 16481 -2604
rect 15773 -2773 15811 -2721
rect 15863 -2773 15875 -2721
rect 15927 -2773 15939 -2721
rect 15991 -2773 16007 -2721
rect 16059 -2773 16071 -2721
rect 16123 -2773 16135 -2721
rect 16187 -2773 16199 -2721
rect 16251 -2773 16267 -2721
rect 16319 -2773 16331 -2721
rect 16383 -2773 16395 -2721
rect 16447 -2773 16481 -2721
rect 15773 -2791 16481 -2773
rect 16603 -2570 17707 -2564
rect 16603 -2604 16784 -2570
rect 16818 -2583 16856 -2570
rect 16890 -2583 17042 -2570
rect 17076 -2583 17114 -2570
rect 17148 -2583 17300 -2570
rect 17334 -2583 17372 -2570
rect 17406 -2583 17558 -2570
rect 17592 -2583 17630 -2570
rect 16847 -2604 16856 -2583
rect 16603 -2635 16795 -2604
rect 16847 -2635 16859 -2604
rect 16911 -2635 16923 -2583
rect 16975 -2635 16991 -2583
rect 17107 -2604 17114 -2583
rect 17043 -2635 17055 -2604
rect 17107 -2635 17119 -2604
rect 17171 -2635 17281 -2583
rect 17334 -2604 17345 -2583
rect 17406 -2604 17409 -2583
rect 17333 -2635 17345 -2604
rect 17397 -2635 17409 -2604
rect 17461 -2635 17477 -2583
rect 17529 -2635 17541 -2583
rect 17593 -2635 17605 -2583
rect 17664 -2604 17707 -2570
rect 17657 -2635 17707 -2604
rect 16603 -2653 17707 -2635
rect 17911 -2570 18347 -2536
rect 17911 -2604 18010 -2570
rect 18044 -2604 18082 -2570
rect 18116 -2574 18347 -2570
rect 18116 -2604 18290 -2574
rect 17911 -2608 18290 -2604
rect 18324 -2608 18347 -2574
rect 17911 -2646 18347 -2608
rect 16603 -2885 16664 -2653
rect 17911 -2680 18290 -2646
rect 18324 -2680 18347 -2646
rect 15590 -2933 16664 -2885
rect 15590 -2967 15816 -2933
rect 15850 -2967 15888 -2933
rect 15922 -2967 16074 -2933
rect 16108 -2967 16146 -2933
rect 16180 -2967 16332 -2933
rect 16366 -2967 16404 -2933
rect 16438 -2967 16664 -2933
rect 15590 -2973 16664 -2967
rect 16741 -2721 17707 -2703
rect 16741 -2773 16795 -2721
rect 16847 -2773 16859 -2721
rect 16911 -2773 16923 -2721
rect 16975 -2773 16991 -2721
rect 17043 -2773 17055 -2721
rect 17107 -2773 17119 -2721
rect 17171 -2773 17281 -2721
rect 17333 -2773 17345 -2721
rect 17397 -2773 17409 -2721
rect 17461 -2773 17477 -2721
rect 17529 -2773 17541 -2721
rect 17593 -2773 17605 -2721
rect 17657 -2773 17707 -2721
rect 16741 -2899 17707 -2773
rect 16741 -2933 16795 -2899
rect 16847 -2933 16859 -2899
rect 16741 -2967 16784 -2933
rect 16847 -2951 16856 -2933
rect 16911 -2951 16923 -2899
rect 16975 -2951 16991 -2899
rect 17043 -2933 17055 -2899
rect 17107 -2933 17119 -2899
rect 17107 -2951 17114 -2933
rect 17171 -2951 17281 -2899
rect 17333 -2933 17345 -2899
rect 17397 -2933 17409 -2899
rect 17334 -2951 17345 -2933
rect 17406 -2951 17409 -2933
rect 17461 -2951 17477 -2899
rect 17529 -2951 17541 -2899
rect 17593 -2951 17605 -2899
rect 17657 -2933 17707 -2899
rect 16818 -2967 16856 -2951
rect 16890 -2967 17042 -2951
rect 17076 -2967 17114 -2951
rect 17148 -2967 17300 -2951
rect 17334 -2967 17372 -2951
rect 17406 -2967 17558 -2951
rect 17592 -2967 17630 -2951
rect 17664 -2967 17707 -2933
rect 16741 -2973 17707 -2967
rect 17911 -2718 18347 -2680
rect 17911 -2752 18290 -2718
rect 18324 -2752 18347 -2718
rect 17911 -2790 18347 -2752
rect 17911 -2824 18290 -2790
rect 18324 -2824 18347 -2790
rect 17911 -2862 18347 -2824
rect 17911 -2896 18290 -2862
rect 18324 -2896 18347 -2862
rect 17911 -2933 18347 -2896
rect 17911 -2967 18010 -2933
rect 18044 -2967 18082 -2933
rect 18116 -2934 18347 -2933
rect 18116 -2967 18290 -2934
rect 17911 -2968 18290 -2967
rect 18324 -2968 18347 -2934
rect 9194 -3061 9986 -3040
rect 9194 -3095 9200 -3061
rect 9234 -3095 9458 -3061
rect 9492 -3078 9688 -3061
rect 9492 -3095 9573 -3078
rect 9194 -3112 9573 -3095
rect 9607 -3095 9688 -3078
rect 9722 -3095 9946 -3061
rect 9980 -3095 9986 -3061
rect 9607 -3112 9986 -3095
rect 9194 -3133 9986 -3112
rect 9194 -3167 9200 -3133
rect 9234 -3167 9458 -3133
rect 9492 -3150 9688 -3133
rect 9492 -3167 9573 -3150
rect 9194 -3184 9573 -3167
rect 9607 -3167 9688 -3150
rect 9722 -3167 9946 -3133
rect 9980 -3167 9986 -3133
rect 9607 -3184 9986 -3167
rect 9194 -3222 9986 -3184
rect 9194 -3256 9573 -3222
rect 9607 -3256 9986 -3222
rect 9194 -3294 9986 -3256
rect 9194 -3328 9573 -3294
rect 9607 -3328 9986 -3294
rect 9194 -3366 9986 -3328
rect 9194 -3400 9573 -3366
rect 9607 -3400 9986 -3366
rect 9194 -3438 9986 -3400
rect 9194 -3472 9573 -3438
rect 9607 -3472 9986 -3438
rect 9194 -3510 9986 -3472
rect 9194 -3544 9573 -3510
rect 9607 -3544 9986 -3510
rect 9194 -3582 9986 -3544
rect 9194 -3616 9573 -3582
rect 9607 -3616 9986 -3582
rect 7894 -3657 8090 -3647
rect 7894 -3709 7901 -3657
rect 7953 -3709 7965 -3657
rect 8017 -3709 8029 -3657
rect 8081 -3709 8090 -3657
rect 7894 -3717 8090 -3709
rect 8410 -3657 8606 -3647
rect 8410 -3709 8417 -3657
rect 8469 -3709 8481 -3657
rect 8533 -3709 8545 -3657
rect 8597 -3709 8606 -3657
rect 8410 -3717 8606 -3709
rect 8928 -3657 9124 -3647
rect 8928 -3709 8935 -3657
rect 8987 -3709 8999 -3657
rect 9051 -3709 9063 -3657
rect 9115 -3709 9124 -3657
rect 8928 -3717 9124 -3709
rect 9194 -3654 9986 -3616
rect 10134 -3061 10180 -3014
rect 10134 -3095 10140 -3061
rect 10174 -3095 10180 -3061
rect 10134 -3133 10180 -3095
rect 10134 -3167 10140 -3133
rect 10174 -3167 10180 -3133
rect 10134 -3647 10180 -3167
rect 10392 -3061 10438 -3014
rect 10392 -3095 10398 -3061
rect 10432 -3095 10438 -3061
rect 10392 -3133 10438 -3095
rect 10392 -3167 10398 -3133
rect 10432 -3167 10438 -3133
rect 10392 -3316 10438 -3167
rect 10650 -3061 10696 -3014
rect 10650 -3095 10656 -3061
rect 10690 -3095 10696 -3061
rect 10650 -3133 10696 -3095
rect 10650 -3167 10656 -3133
rect 10690 -3167 10696 -3133
rect 10316 -3326 10512 -3316
rect 10316 -3378 10325 -3326
rect 10377 -3378 10389 -3326
rect 10441 -3378 10453 -3326
rect 10505 -3378 10512 -3326
rect 10316 -3386 10512 -3378
rect 10650 -3647 10696 -3167
rect 10908 -3061 10954 -3014
rect 10908 -3095 10914 -3061
rect 10948 -3095 10954 -3061
rect 10908 -3133 10954 -3095
rect 10908 -3167 10914 -3133
rect 10948 -3167 10954 -3133
rect 10908 -3316 10954 -3167
rect 11166 -3061 11212 -3014
rect 11166 -3095 11172 -3061
rect 11206 -3095 11212 -3061
rect 11166 -3133 11212 -3095
rect 11166 -3167 11172 -3133
rect 11206 -3167 11212 -3133
rect 10833 -3326 11029 -3316
rect 10833 -3378 10842 -3326
rect 10894 -3378 10906 -3326
rect 10958 -3378 10970 -3326
rect 11022 -3378 11029 -3326
rect 10833 -3386 11029 -3378
rect 11166 -3647 11212 -3167
rect 11360 -3061 11406 -3014
rect 11360 -3095 11366 -3061
rect 11400 -3095 11406 -3061
rect 11360 -3133 11406 -3095
rect 11360 -3167 11366 -3133
rect 11400 -3167 11406 -3133
rect 11360 -3485 11406 -3167
rect 11618 -3061 11664 -3014
rect 11618 -3095 11624 -3061
rect 11658 -3095 11664 -3061
rect 11618 -3133 11664 -3095
rect 11618 -3167 11624 -3133
rect 11658 -3167 11664 -3133
rect 11287 -3495 11483 -3485
rect 11287 -3547 11294 -3495
rect 11346 -3547 11358 -3495
rect 11410 -3547 11422 -3495
rect 11474 -3547 11483 -3495
rect 11287 -3555 11483 -3547
rect 9194 -3688 9573 -3654
rect 9607 -3688 9986 -3654
rect 9194 -3726 9986 -3688
rect 10056 -3657 10252 -3647
rect 10056 -3709 10065 -3657
rect 10117 -3709 10129 -3657
rect 10181 -3709 10193 -3657
rect 10245 -3709 10252 -3657
rect 10056 -3717 10252 -3709
rect 10574 -3657 10770 -3647
rect 10574 -3709 10583 -3657
rect 10635 -3709 10647 -3657
rect 10699 -3709 10711 -3657
rect 10763 -3709 10770 -3657
rect 10574 -3717 10770 -3709
rect 11090 -3657 11286 -3647
rect 11090 -3709 11099 -3657
rect 11151 -3709 11163 -3657
rect 11215 -3709 11227 -3657
rect 11279 -3709 11286 -3657
rect 11090 -3717 11286 -3709
rect 9194 -3760 9573 -3726
rect 9607 -3760 9986 -3726
rect 9194 -3798 9986 -3760
rect 4836 -3870 5626 -3832
rect 833 -3942 1269 -3904
rect 833 -3976 856 -3942
rect 890 -3976 1269 -3942
rect 833 -4014 1269 -3976
rect 4836 -3904 5214 -3870
rect 5248 -3904 5626 -3870
rect 6922 -3826 7118 -3816
rect 6922 -3878 6931 -3826
rect 6983 -3878 6995 -3826
rect 7047 -3878 7059 -3826
rect 7111 -3878 7118 -3826
rect 6922 -3886 7118 -3878
rect 7440 -3826 7636 -3816
rect 7440 -3878 7449 -3826
rect 7501 -3878 7513 -3826
rect 7565 -3878 7577 -3826
rect 7629 -3878 7636 -3826
rect 7440 -3886 7636 -3878
rect 9194 -3832 9573 -3798
rect 9607 -3832 9986 -3798
rect 11618 -3816 11664 -3167
rect 11876 -3061 11922 -3014
rect 11876 -3095 11882 -3061
rect 11916 -3095 11922 -3061
rect 11876 -3133 11922 -3095
rect 11876 -3167 11882 -3133
rect 11916 -3167 11922 -3133
rect 11876 -3485 11922 -3167
rect 12134 -3061 12180 -3014
rect 12134 -3095 12140 -3061
rect 12174 -3095 12180 -3061
rect 12134 -3133 12180 -3095
rect 12134 -3167 12140 -3133
rect 12174 -3167 12180 -3133
rect 11804 -3495 12000 -3485
rect 11804 -3547 11811 -3495
rect 11863 -3547 11875 -3495
rect 11927 -3547 11939 -3495
rect 11991 -3547 12000 -3495
rect 11804 -3555 12000 -3547
rect 12134 -3816 12180 -3167
rect 12328 -3061 12374 -3014
rect 12328 -3095 12334 -3061
rect 12368 -3095 12374 -3061
rect 12328 -3133 12374 -3095
rect 12328 -3167 12334 -3133
rect 12368 -3167 12374 -3133
rect 12328 -3647 12374 -3167
rect 12586 -3061 12632 -3014
rect 12586 -3095 12592 -3061
rect 12626 -3095 12632 -3061
rect 12586 -3133 12632 -3095
rect 12586 -3167 12592 -3133
rect 12626 -3167 12632 -3133
rect 12586 -3316 12632 -3167
rect 12844 -3061 12890 -3014
rect 12844 -3095 12850 -3061
rect 12884 -3095 12890 -3061
rect 12844 -3133 12890 -3095
rect 12844 -3167 12850 -3133
rect 12884 -3167 12890 -3133
rect 12510 -3326 12706 -3316
rect 12510 -3378 12519 -3326
rect 12571 -3378 12583 -3326
rect 12635 -3378 12647 -3326
rect 12699 -3378 12706 -3326
rect 12510 -3386 12706 -3378
rect 12844 -3647 12890 -3167
rect 13102 -3061 13148 -3014
rect 13102 -3095 13108 -3061
rect 13142 -3095 13148 -3061
rect 13102 -3133 13148 -3095
rect 13102 -3167 13108 -3133
rect 13142 -3167 13148 -3133
rect 13102 -3316 13148 -3167
rect 13360 -3061 13406 -3014
rect 13360 -3095 13366 -3061
rect 13400 -3095 13406 -3061
rect 13360 -3133 13406 -3095
rect 13360 -3167 13366 -3133
rect 13400 -3167 13406 -3133
rect 13027 -3326 13223 -3316
rect 13027 -3378 13036 -3326
rect 13088 -3378 13100 -3326
rect 13152 -3378 13164 -3326
rect 13216 -3378 13223 -3326
rect 13027 -3386 13223 -3378
rect 13360 -3647 13406 -3167
rect 13554 -3040 13932 -3006
rect 13966 -3040 14344 -3006
rect 17911 -3006 18347 -2968
rect 13554 -3061 14344 -3040
rect 13554 -3095 13560 -3061
rect 13594 -3095 13818 -3061
rect 13852 -3078 14046 -3061
rect 13852 -3095 13932 -3078
rect 13554 -3112 13932 -3095
rect 13966 -3095 14046 -3078
rect 14080 -3095 14304 -3061
rect 14338 -3095 14344 -3061
rect 13966 -3112 14344 -3095
rect 13554 -3133 14344 -3112
rect 13554 -3167 13560 -3133
rect 13594 -3167 13818 -3133
rect 13852 -3150 14046 -3133
rect 13852 -3167 13932 -3150
rect 13554 -3184 13932 -3167
rect 13966 -3167 14046 -3150
rect 14080 -3167 14304 -3133
rect 14338 -3167 14344 -3133
rect 13966 -3184 14344 -3167
rect 13554 -3222 14344 -3184
rect 13554 -3256 13932 -3222
rect 13966 -3256 14344 -3222
rect 13554 -3294 14344 -3256
rect 13554 -3328 13932 -3294
rect 13966 -3328 14344 -3294
rect 13554 -3366 14344 -3328
rect 13554 -3400 13932 -3366
rect 13966 -3400 14344 -3366
rect 13554 -3438 14344 -3400
rect 13554 -3472 13932 -3438
rect 13966 -3472 14344 -3438
rect 13554 -3510 14344 -3472
rect 13554 -3544 13932 -3510
rect 13966 -3544 14344 -3510
rect 13554 -3582 14344 -3544
rect 13554 -3616 13932 -3582
rect 13966 -3616 14344 -3582
rect 12251 -3657 12447 -3647
rect 12251 -3709 12260 -3657
rect 12312 -3709 12324 -3657
rect 12376 -3709 12388 -3657
rect 12440 -3709 12447 -3657
rect 12251 -3717 12447 -3709
rect 12768 -3657 12964 -3647
rect 12768 -3709 12777 -3657
rect 12829 -3709 12841 -3657
rect 12893 -3709 12905 -3657
rect 12957 -3709 12964 -3657
rect 12768 -3717 12964 -3709
rect 13283 -3657 13479 -3647
rect 13283 -3709 13292 -3657
rect 13344 -3709 13356 -3657
rect 13408 -3709 13420 -3657
rect 13472 -3709 13479 -3657
rect 13283 -3717 13479 -3709
rect 13554 -3654 14344 -3616
rect 14491 -3061 14537 -3014
rect 14491 -3095 14497 -3061
rect 14531 -3095 14537 -3061
rect 14491 -3133 14537 -3095
rect 14491 -3167 14497 -3133
rect 14531 -3167 14537 -3133
rect 14491 -3647 14537 -3167
rect 14749 -3061 14795 -3014
rect 14749 -3095 14755 -3061
rect 14789 -3095 14795 -3061
rect 14749 -3133 14795 -3095
rect 14749 -3167 14755 -3133
rect 14789 -3167 14795 -3133
rect 14749 -3316 14795 -3167
rect 15007 -3061 15053 -3014
rect 15007 -3095 15013 -3061
rect 15047 -3095 15053 -3061
rect 15007 -3133 15053 -3095
rect 15007 -3167 15013 -3133
rect 15047 -3167 15053 -3133
rect 14674 -3326 14870 -3316
rect 14674 -3378 14681 -3326
rect 14733 -3378 14745 -3326
rect 14797 -3378 14809 -3326
rect 14861 -3378 14870 -3326
rect 14674 -3386 14870 -3378
rect 15007 -3647 15053 -3167
rect 15265 -3061 15311 -3014
rect 15265 -3095 15271 -3061
rect 15305 -3095 15311 -3061
rect 15265 -3133 15311 -3095
rect 15265 -3167 15271 -3133
rect 15305 -3167 15311 -3133
rect 15265 -3316 15311 -3167
rect 15523 -3061 15569 -3014
rect 15523 -3095 15529 -3061
rect 15563 -3095 15569 -3061
rect 15523 -3133 15569 -3095
rect 15523 -3167 15529 -3133
rect 15563 -3167 15569 -3133
rect 15191 -3326 15387 -3316
rect 15191 -3378 15198 -3326
rect 15250 -3378 15262 -3326
rect 15314 -3378 15326 -3326
rect 15378 -3378 15387 -3326
rect 15191 -3386 15387 -3378
rect 15523 -3647 15569 -3167
rect 15717 -3061 15763 -3014
rect 15717 -3095 15723 -3061
rect 15757 -3095 15763 -3061
rect 15717 -3133 15763 -3095
rect 15717 -3167 15723 -3133
rect 15757 -3167 15763 -3133
rect 13554 -3688 13932 -3654
rect 13966 -3688 14344 -3654
rect 13554 -3726 14344 -3688
rect 14418 -3657 14614 -3647
rect 14418 -3709 14425 -3657
rect 14477 -3709 14489 -3657
rect 14541 -3709 14553 -3657
rect 14605 -3709 14614 -3657
rect 14418 -3717 14614 -3709
rect 14933 -3657 15129 -3647
rect 14933 -3709 14940 -3657
rect 14992 -3709 15004 -3657
rect 15056 -3709 15068 -3657
rect 15120 -3709 15129 -3657
rect 14933 -3717 15129 -3709
rect 15450 -3657 15646 -3647
rect 15450 -3709 15457 -3657
rect 15509 -3709 15521 -3657
rect 15573 -3709 15585 -3657
rect 15637 -3709 15646 -3657
rect 15450 -3717 15646 -3709
rect 13554 -3760 13932 -3726
rect 13966 -3760 14344 -3726
rect 13554 -3798 14344 -3760
rect 9194 -3870 9986 -3832
rect 4836 -3942 5626 -3904
rect 4836 -3976 5214 -3942
rect 5248 -3976 5626 -3942
rect 833 -4048 856 -4014
rect 890 -4048 1269 -4014
rect 833 -4051 1269 -4048
rect 833 -4085 971 -4051
rect 1005 -4085 1229 -4051
rect 1263 -4085 1269 -4051
rect 833 -4086 1269 -4085
rect 833 -4120 856 -4086
rect 890 -4120 1269 -4086
rect 833 -4123 1269 -4120
rect 833 -4157 971 -4123
rect 1005 -4157 1229 -4123
rect 1263 -4157 1269 -4123
rect 833 -4158 1269 -4157
rect 833 -4192 856 -4158
rect 890 -4192 1269 -4158
rect 833 -4230 1269 -4192
rect 833 -4245 856 -4230
rect 831 -4264 856 -4245
rect 890 -4245 1269 -4230
rect 1417 -4051 1463 -4004
rect 1417 -4085 1423 -4051
rect 1457 -4085 1463 -4051
rect 1417 -4123 1463 -4085
rect 1417 -4157 1423 -4123
rect 1457 -4157 1463 -4123
rect 1417 -4245 1463 -4157
rect 1675 -4051 1721 -4004
rect 1675 -4085 1681 -4051
rect 1715 -4085 1721 -4051
rect 1675 -4123 1721 -4085
rect 1675 -4157 1681 -4123
rect 1715 -4157 1721 -4123
rect 1675 -4245 1721 -4157
rect 1933 -4051 1979 -4004
rect 1933 -4085 1939 -4051
rect 1973 -4085 1979 -4051
rect 1933 -4123 1979 -4085
rect 1933 -4157 1939 -4123
rect 1973 -4157 1979 -4123
rect 1933 -4245 1979 -4157
rect 2191 -4051 2237 -4004
rect 2191 -4085 2197 -4051
rect 2231 -4085 2237 -4051
rect 2191 -4123 2237 -4085
rect 2191 -4157 2197 -4123
rect 2231 -4157 2237 -4123
rect 2191 -4245 2237 -4157
rect 2449 -4051 2495 -4004
rect 2449 -4085 2455 -4051
rect 2489 -4085 2495 -4051
rect 2449 -4123 2495 -4085
rect 2449 -4157 2455 -4123
rect 2489 -4157 2495 -4123
rect 2449 -4245 2495 -4157
rect 2643 -4051 2689 -4004
rect 2643 -4085 2649 -4051
rect 2683 -4085 2689 -4051
rect 2643 -4123 2689 -4085
rect 2643 -4157 2649 -4123
rect 2683 -4157 2689 -4123
rect 2643 -4245 2689 -4157
rect 2901 -4051 2947 -4004
rect 2901 -4085 2907 -4051
rect 2941 -4085 2947 -4051
rect 2901 -4123 2947 -4085
rect 2901 -4157 2907 -4123
rect 2941 -4157 2947 -4123
rect 2901 -4245 2947 -4157
rect 3159 -4051 3205 -4004
rect 3159 -4085 3165 -4051
rect 3199 -4085 3205 -4051
rect 3159 -4123 3205 -4085
rect 3159 -4157 3165 -4123
rect 3199 -4157 3205 -4123
rect 3159 -4245 3205 -4157
rect 3417 -4051 3463 -4004
rect 3417 -4085 3423 -4051
rect 3457 -4085 3463 -4051
rect 3417 -4123 3463 -4085
rect 3417 -4157 3423 -4123
rect 3457 -4157 3463 -4123
rect 3417 -4245 3463 -4157
rect 3611 -4051 3657 -4004
rect 3611 -4085 3617 -4051
rect 3651 -4085 3657 -4051
rect 3611 -4123 3657 -4085
rect 3611 -4157 3617 -4123
rect 3651 -4157 3657 -4123
rect 3611 -4245 3657 -4157
rect 3869 -4051 3915 -4004
rect 3869 -4085 3875 -4051
rect 3909 -4085 3915 -4051
rect 3869 -4123 3915 -4085
rect 3869 -4157 3875 -4123
rect 3909 -4157 3915 -4123
rect 3869 -4245 3915 -4157
rect 4127 -4051 4173 -4004
rect 4127 -4085 4133 -4051
rect 4167 -4085 4173 -4051
rect 4127 -4123 4173 -4085
rect 4127 -4157 4133 -4123
rect 4167 -4157 4173 -4123
rect 4127 -4245 4173 -4157
rect 4385 -4051 4431 -4004
rect 4385 -4085 4391 -4051
rect 4425 -4085 4431 -4051
rect 4385 -4123 4431 -4085
rect 4385 -4157 4391 -4123
rect 4425 -4157 4431 -4123
rect 4385 -4245 4431 -4157
rect 4643 -4051 4689 -4004
rect 4643 -4085 4649 -4051
rect 4683 -4085 4689 -4051
rect 4643 -4123 4689 -4085
rect 4643 -4157 4649 -4123
rect 4683 -4157 4689 -4123
rect 4643 -4245 4689 -4157
rect 4836 -4014 5626 -3976
rect 9194 -3904 9573 -3870
rect 9607 -3904 9986 -3870
rect 11544 -3826 11740 -3816
rect 11544 -3878 11551 -3826
rect 11603 -3878 11615 -3826
rect 11667 -3878 11679 -3826
rect 11731 -3878 11740 -3826
rect 11544 -3886 11740 -3878
rect 12062 -3826 12258 -3816
rect 12062 -3878 12069 -3826
rect 12121 -3878 12133 -3826
rect 12185 -3878 12197 -3826
rect 12249 -3878 12258 -3826
rect 12062 -3886 12258 -3878
rect 13554 -3832 13932 -3798
rect 13966 -3832 14344 -3798
rect 15717 -3816 15763 -3167
rect 15975 -3061 16021 -3014
rect 15975 -3095 15981 -3061
rect 16015 -3095 16021 -3061
rect 15975 -3133 16021 -3095
rect 15975 -3167 15981 -3133
rect 16015 -3167 16021 -3133
rect 15975 -3485 16021 -3167
rect 16233 -3061 16279 -3014
rect 16233 -3095 16239 -3061
rect 16273 -3095 16279 -3061
rect 16233 -3133 16279 -3095
rect 16233 -3167 16239 -3133
rect 16273 -3167 16279 -3133
rect 15897 -3495 16093 -3485
rect 15897 -3547 15906 -3495
rect 15958 -3547 15970 -3495
rect 16022 -3547 16034 -3495
rect 16086 -3547 16093 -3495
rect 15897 -3555 16093 -3547
rect 16233 -3816 16279 -3167
rect 16491 -3061 16537 -3014
rect 16491 -3095 16497 -3061
rect 16531 -3095 16537 -3061
rect 16491 -3133 16537 -3095
rect 16491 -3167 16497 -3133
rect 16531 -3167 16537 -3133
rect 16491 -3485 16537 -3167
rect 16685 -3061 16731 -3014
rect 16685 -3095 16691 -3061
rect 16725 -3095 16731 -3061
rect 16685 -3133 16731 -3095
rect 16685 -3167 16691 -3133
rect 16725 -3167 16731 -3133
rect 16414 -3495 16610 -3485
rect 16414 -3547 16423 -3495
rect 16475 -3547 16487 -3495
rect 16539 -3547 16551 -3495
rect 16603 -3547 16610 -3495
rect 16414 -3555 16610 -3547
rect 16685 -3647 16731 -3167
rect 16943 -3061 16989 -3014
rect 16943 -3095 16949 -3061
rect 16983 -3095 16989 -3061
rect 16943 -3133 16989 -3095
rect 16943 -3167 16949 -3133
rect 16983 -3167 16989 -3133
rect 16943 -3316 16989 -3167
rect 17201 -3061 17247 -3014
rect 17201 -3095 17207 -3061
rect 17241 -3095 17247 -3061
rect 17201 -3133 17247 -3095
rect 17201 -3167 17207 -3133
rect 17241 -3167 17247 -3133
rect 16868 -3326 17064 -3316
rect 16868 -3378 16875 -3326
rect 16927 -3378 16939 -3326
rect 16991 -3378 17003 -3326
rect 17055 -3378 17064 -3326
rect 16868 -3386 17064 -3378
rect 17201 -3647 17247 -3167
rect 17459 -3061 17505 -3014
rect 17459 -3095 17465 -3061
rect 17499 -3095 17505 -3061
rect 17459 -3133 17505 -3095
rect 17459 -3167 17465 -3133
rect 17499 -3167 17505 -3133
rect 17459 -3316 17505 -3167
rect 17717 -3061 17763 -3014
rect 17717 -3095 17723 -3061
rect 17757 -3095 17763 -3061
rect 17717 -3133 17763 -3095
rect 17717 -3167 17723 -3133
rect 17757 -3167 17763 -3133
rect 17386 -3326 17582 -3316
rect 17386 -3378 17393 -3326
rect 17445 -3378 17457 -3326
rect 17509 -3378 17521 -3326
rect 17573 -3378 17582 -3326
rect 17386 -3386 17582 -3378
rect 17717 -3647 17763 -3167
rect 17911 -3040 18290 -3006
rect 18324 -3040 18347 -3006
rect 17911 -3061 18347 -3040
rect 17911 -3095 17917 -3061
rect 17951 -3095 18175 -3061
rect 18209 -3078 18347 -3061
rect 18209 -3095 18290 -3078
rect 17911 -3112 18290 -3095
rect 18324 -3112 18347 -3078
rect 17911 -3133 18347 -3112
rect 17911 -3167 17917 -3133
rect 17951 -3167 18175 -3133
rect 18209 -3150 18347 -3133
rect 18209 -3167 18290 -3150
rect 17911 -3184 18290 -3167
rect 18324 -3184 18347 -3150
rect 17911 -3222 18347 -3184
rect 17911 -3256 18290 -3222
rect 18324 -3256 18347 -3222
rect 17911 -3294 18347 -3256
rect 17911 -3328 18290 -3294
rect 18324 -3328 18347 -3294
rect 17911 -3366 18347 -3328
rect 17911 -3400 18290 -3366
rect 18324 -3400 18347 -3366
rect 17911 -3438 18347 -3400
rect 17911 -3472 18290 -3438
rect 18324 -3472 18347 -3438
rect 17911 -3510 18347 -3472
rect 17911 -3544 18290 -3510
rect 18324 -3544 18347 -3510
rect 17911 -3582 18347 -3544
rect 17911 -3616 18290 -3582
rect 18324 -3616 18347 -3582
rect 16611 -3657 16807 -3647
rect 16611 -3709 16618 -3657
rect 16670 -3709 16682 -3657
rect 16734 -3709 16746 -3657
rect 16798 -3709 16807 -3657
rect 16611 -3717 16807 -3709
rect 17128 -3657 17324 -3647
rect 17128 -3709 17135 -3657
rect 17187 -3709 17199 -3657
rect 17251 -3709 17263 -3657
rect 17315 -3709 17324 -3657
rect 17128 -3717 17324 -3709
rect 17645 -3657 17841 -3647
rect 17645 -3709 17652 -3657
rect 17704 -3709 17716 -3657
rect 17768 -3709 17780 -3657
rect 17832 -3709 17841 -3657
rect 17645 -3717 17841 -3709
rect 17911 -3654 18347 -3616
rect 17911 -3688 18290 -3654
rect 18324 -3688 18347 -3654
rect 17911 -3726 18347 -3688
rect 17911 -3760 18290 -3726
rect 18324 -3760 18347 -3726
rect 17911 -3798 18347 -3760
rect 13554 -3870 14344 -3832
rect 9194 -3942 9986 -3904
rect 9194 -3976 9573 -3942
rect 9607 -3976 9986 -3942
rect 4836 -4048 5214 -4014
rect 5248 -4048 5626 -4014
rect 4836 -4051 5626 -4048
rect 4836 -4085 4842 -4051
rect 4876 -4085 5100 -4051
rect 5134 -4085 5328 -4051
rect 5362 -4085 5586 -4051
rect 5620 -4085 5626 -4051
rect 4836 -4086 5626 -4085
rect 4836 -4120 5214 -4086
rect 5248 -4120 5626 -4086
rect 4836 -4123 5626 -4120
rect 4836 -4157 4842 -4123
rect 4876 -4157 5100 -4123
rect 5134 -4157 5328 -4123
rect 5362 -4157 5586 -4123
rect 5620 -4157 5626 -4123
rect 4836 -4158 5626 -4157
rect 4836 -4192 5214 -4158
rect 5248 -4192 5626 -4158
rect 4836 -4230 5626 -4192
rect 4836 -4245 5214 -4230
rect 890 -4251 5214 -4245
rect 890 -4264 1064 -4251
rect 831 -4285 1064 -4264
rect 1098 -4285 1136 -4251
rect 1170 -4285 1516 -4251
rect 1550 -4285 1588 -4251
rect 1622 -4285 1774 -4251
rect 1808 -4285 1846 -4251
rect 1880 -4285 2032 -4251
rect 2066 -4285 2104 -4251
rect 2138 -4285 2290 -4251
rect 2324 -4285 2362 -4251
rect 2396 -4285 2742 -4251
rect 2776 -4285 2814 -4251
rect 2848 -4285 3000 -4251
rect 3034 -4285 3072 -4251
rect 3106 -4285 3258 -4251
rect 3292 -4285 3330 -4251
rect 3364 -4285 3710 -4251
rect 3744 -4285 3782 -4251
rect 3816 -4285 3968 -4251
rect 4002 -4285 4040 -4251
rect 4074 -4285 4226 -4251
rect 4260 -4285 4298 -4251
rect 4332 -4285 4484 -4251
rect 4518 -4285 4556 -4251
rect 4590 -4285 4935 -4251
rect 4969 -4285 5007 -4251
rect 5041 -4264 5214 -4251
rect 5248 -4245 5626 -4230
rect 5774 -4051 5820 -4004
rect 5774 -4085 5780 -4051
rect 5814 -4085 5820 -4051
rect 5774 -4123 5820 -4085
rect 5774 -4157 5780 -4123
rect 5814 -4157 5820 -4123
rect 5774 -4245 5820 -4157
rect 6032 -4051 6078 -4004
rect 6032 -4085 6038 -4051
rect 6072 -4085 6078 -4051
rect 6032 -4123 6078 -4085
rect 6032 -4157 6038 -4123
rect 6072 -4157 6078 -4123
rect 6032 -4245 6078 -4157
rect 6290 -4051 6336 -4004
rect 6290 -4085 6296 -4051
rect 6330 -4085 6336 -4051
rect 6290 -4123 6336 -4085
rect 6290 -4157 6296 -4123
rect 6330 -4157 6336 -4123
rect 6290 -4245 6336 -4157
rect 6548 -4051 6594 -4004
rect 6548 -4085 6554 -4051
rect 6588 -4085 6594 -4051
rect 6548 -4123 6594 -4085
rect 6548 -4157 6554 -4123
rect 6588 -4157 6594 -4123
rect 6548 -4245 6594 -4157
rect 6806 -4051 6852 -4004
rect 6806 -4085 6812 -4051
rect 6846 -4085 6852 -4051
rect 6806 -4123 6852 -4085
rect 6806 -4157 6812 -4123
rect 6846 -4157 6852 -4123
rect 6806 -4245 6852 -4157
rect 7000 -4051 7046 -4004
rect 7000 -4085 7006 -4051
rect 7040 -4085 7046 -4051
rect 7000 -4123 7046 -4085
rect 7000 -4157 7006 -4123
rect 7040 -4157 7046 -4123
rect 7000 -4245 7046 -4157
rect 7258 -4051 7304 -4004
rect 7258 -4085 7264 -4051
rect 7298 -4085 7304 -4051
rect 7258 -4123 7304 -4085
rect 7258 -4157 7264 -4123
rect 7298 -4157 7304 -4123
rect 7258 -4245 7304 -4157
rect 7516 -4051 7562 -4004
rect 7516 -4085 7522 -4051
rect 7556 -4085 7562 -4051
rect 7516 -4123 7562 -4085
rect 7516 -4157 7522 -4123
rect 7556 -4157 7562 -4123
rect 7516 -4245 7562 -4157
rect 7774 -4051 7820 -4004
rect 7774 -4085 7780 -4051
rect 7814 -4085 7820 -4051
rect 7774 -4123 7820 -4085
rect 7774 -4157 7780 -4123
rect 7814 -4157 7820 -4123
rect 7774 -4245 7820 -4157
rect 7968 -4051 8014 -4004
rect 7968 -4085 7974 -4051
rect 8008 -4085 8014 -4051
rect 7968 -4123 8014 -4085
rect 7968 -4157 7974 -4123
rect 8008 -4157 8014 -4123
rect 7968 -4245 8014 -4157
rect 8226 -4051 8272 -4004
rect 8226 -4085 8232 -4051
rect 8266 -4085 8272 -4051
rect 8226 -4123 8272 -4085
rect 8226 -4157 8232 -4123
rect 8266 -4157 8272 -4123
rect 8226 -4245 8272 -4157
rect 8484 -4051 8530 -4004
rect 8484 -4085 8490 -4051
rect 8524 -4085 8530 -4051
rect 8484 -4123 8530 -4085
rect 8484 -4157 8490 -4123
rect 8524 -4157 8530 -4123
rect 8484 -4245 8530 -4157
rect 8742 -4051 8788 -4004
rect 8742 -4085 8748 -4051
rect 8782 -4085 8788 -4051
rect 8742 -4123 8788 -4085
rect 8742 -4157 8748 -4123
rect 8782 -4157 8788 -4123
rect 8742 -4245 8788 -4157
rect 9000 -4051 9046 -4004
rect 9000 -4085 9006 -4051
rect 9040 -4085 9046 -4051
rect 9000 -4123 9046 -4085
rect 9000 -4157 9006 -4123
rect 9040 -4157 9046 -4123
rect 9000 -4245 9046 -4157
rect 9194 -4014 9986 -3976
rect 13554 -3904 13932 -3870
rect 13966 -3904 14344 -3870
rect 15640 -3826 15836 -3816
rect 15640 -3878 15649 -3826
rect 15701 -3878 15713 -3826
rect 15765 -3878 15777 -3826
rect 15829 -3878 15836 -3826
rect 15640 -3886 15836 -3878
rect 16157 -3826 16353 -3816
rect 16157 -3878 16166 -3826
rect 16218 -3878 16230 -3826
rect 16282 -3878 16294 -3826
rect 16346 -3878 16353 -3826
rect 16157 -3886 16353 -3878
rect 17911 -3832 18290 -3798
rect 18324 -3832 18347 -3798
rect 17911 -3870 18347 -3832
rect 13554 -3942 14344 -3904
rect 13554 -3976 13932 -3942
rect 13966 -3976 14344 -3942
rect 9194 -4048 9573 -4014
rect 9607 -4048 9986 -4014
rect 9194 -4051 9986 -4048
rect 9194 -4085 9200 -4051
rect 9234 -4085 9458 -4051
rect 9492 -4085 9688 -4051
rect 9722 -4085 9946 -4051
rect 9980 -4085 9986 -4051
rect 9194 -4086 9986 -4085
rect 9194 -4120 9573 -4086
rect 9607 -4120 9986 -4086
rect 9194 -4123 9986 -4120
rect 9194 -4157 9200 -4123
rect 9234 -4157 9458 -4123
rect 9492 -4157 9688 -4123
rect 9722 -4157 9946 -4123
rect 9980 -4157 9986 -4123
rect 9194 -4158 9986 -4157
rect 9194 -4192 9573 -4158
rect 9607 -4192 9986 -4158
rect 9194 -4230 9986 -4192
rect 9194 -4245 9573 -4230
rect 5248 -4251 9573 -4245
rect 5248 -4264 5421 -4251
rect 5041 -4285 5421 -4264
rect 5455 -4285 5493 -4251
rect 5527 -4285 5873 -4251
rect 5907 -4285 5945 -4251
rect 5979 -4285 6131 -4251
rect 6165 -4285 6203 -4251
rect 6237 -4285 6389 -4251
rect 6423 -4285 6461 -4251
rect 6495 -4285 6647 -4251
rect 6681 -4285 6719 -4251
rect 6753 -4285 7099 -4251
rect 7133 -4285 7171 -4251
rect 7205 -4285 7357 -4251
rect 7391 -4285 7429 -4251
rect 7463 -4285 7615 -4251
rect 7649 -4285 7687 -4251
rect 7721 -4285 8067 -4251
rect 8101 -4285 8139 -4251
rect 8173 -4285 8325 -4251
rect 8359 -4285 8397 -4251
rect 8431 -4285 8583 -4251
rect 8617 -4285 8655 -4251
rect 8689 -4285 8841 -4251
rect 8875 -4285 8913 -4251
rect 8947 -4285 9293 -4251
rect 9327 -4285 9365 -4251
rect 9399 -4264 9573 -4251
rect 9607 -4245 9986 -4230
rect 10134 -4051 10180 -4004
rect 10134 -4085 10140 -4051
rect 10174 -4085 10180 -4051
rect 10134 -4123 10180 -4085
rect 10134 -4157 10140 -4123
rect 10174 -4157 10180 -4123
rect 10134 -4245 10180 -4157
rect 10392 -4051 10438 -4004
rect 10392 -4085 10398 -4051
rect 10432 -4085 10438 -4051
rect 10392 -4123 10438 -4085
rect 10392 -4157 10398 -4123
rect 10432 -4157 10438 -4123
rect 10392 -4245 10438 -4157
rect 10650 -4051 10696 -4004
rect 10650 -4085 10656 -4051
rect 10690 -4085 10696 -4051
rect 10650 -4123 10696 -4085
rect 10650 -4157 10656 -4123
rect 10690 -4157 10696 -4123
rect 10650 -4245 10696 -4157
rect 10908 -4051 10954 -4004
rect 10908 -4085 10914 -4051
rect 10948 -4085 10954 -4051
rect 10908 -4123 10954 -4085
rect 10908 -4157 10914 -4123
rect 10948 -4157 10954 -4123
rect 10908 -4245 10954 -4157
rect 11166 -4051 11212 -4004
rect 11166 -4085 11172 -4051
rect 11206 -4085 11212 -4051
rect 11166 -4123 11212 -4085
rect 11166 -4157 11172 -4123
rect 11206 -4157 11212 -4123
rect 11166 -4245 11212 -4157
rect 11360 -4051 11406 -4004
rect 11360 -4085 11366 -4051
rect 11400 -4085 11406 -4051
rect 11360 -4123 11406 -4085
rect 11360 -4157 11366 -4123
rect 11400 -4157 11406 -4123
rect 11360 -4245 11406 -4157
rect 11618 -4051 11664 -4004
rect 11618 -4085 11624 -4051
rect 11658 -4085 11664 -4051
rect 11618 -4123 11664 -4085
rect 11618 -4157 11624 -4123
rect 11658 -4157 11664 -4123
rect 11618 -4245 11664 -4157
rect 11876 -4051 11922 -4004
rect 11876 -4085 11882 -4051
rect 11916 -4085 11922 -4051
rect 11876 -4123 11922 -4085
rect 11876 -4157 11882 -4123
rect 11916 -4157 11922 -4123
rect 11876 -4245 11922 -4157
rect 12134 -4051 12180 -4004
rect 12134 -4085 12140 -4051
rect 12174 -4085 12180 -4051
rect 12134 -4123 12180 -4085
rect 12134 -4157 12140 -4123
rect 12174 -4157 12180 -4123
rect 12134 -4245 12180 -4157
rect 12328 -4051 12374 -4004
rect 12328 -4085 12334 -4051
rect 12368 -4085 12374 -4051
rect 12328 -4123 12374 -4085
rect 12328 -4157 12334 -4123
rect 12368 -4157 12374 -4123
rect 12328 -4245 12374 -4157
rect 12586 -4051 12632 -4004
rect 12586 -4085 12592 -4051
rect 12626 -4085 12632 -4051
rect 12586 -4123 12632 -4085
rect 12586 -4157 12592 -4123
rect 12626 -4157 12632 -4123
rect 12586 -4245 12632 -4157
rect 12844 -4051 12890 -4004
rect 12844 -4085 12850 -4051
rect 12884 -4085 12890 -4051
rect 12844 -4123 12890 -4085
rect 12844 -4157 12850 -4123
rect 12884 -4157 12890 -4123
rect 12844 -4245 12890 -4157
rect 13102 -4051 13148 -4004
rect 13102 -4085 13108 -4051
rect 13142 -4085 13148 -4051
rect 13102 -4123 13148 -4085
rect 13102 -4157 13108 -4123
rect 13142 -4157 13148 -4123
rect 13102 -4245 13148 -4157
rect 13360 -4051 13406 -4004
rect 13360 -4085 13366 -4051
rect 13400 -4085 13406 -4051
rect 13360 -4123 13406 -4085
rect 13360 -4157 13366 -4123
rect 13400 -4157 13406 -4123
rect 13360 -4245 13406 -4157
rect 13554 -4014 14344 -3976
rect 17911 -3904 18290 -3870
rect 18324 -3904 18347 -3870
rect 17911 -3942 18347 -3904
rect 17911 -3976 18290 -3942
rect 18324 -3976 18347 -3942
rect 13554 -4048 13932 -4014
rect 13966 -4048 14344 -4014
rect 13554 -4051 14344 -4048
rect 13554 -4085 13560 -4051
rect 13594 -4085 13818 -4051
rect 13852 -4085 14046 -4051
rect 14080 -4085 14304 -4051
rect 14338 -4085 14344 -4051
rect 13554 -4086 14344 -4085
rect 13554 -4120 13932 -4086
rect 13966 -4120 14344 -4086
rect 13554 -4123 14344 -4120
rect 13554 -4157 13560 -4123
rect 13594 -4157 13818 -4123
rect 13852 -4157 14046 -4123
rect 14080 -4157 14304 -4123
rect 14338 -4157 14344 -4123
rect 13554 -4158 14344 -4157
rect 13554 -4192 13932 -4158
rect 13966 -4192 14344 -4158
rect 13554 -4230 14344 -4192
rect 13554 -4245 13932 -4230
rect 9607 -4251 13932 -4245
rect 9607 -4264 9781 -4251
rect 9399 -4285 9781 -4264
rect 9815 -4285 9853 -4251
rect 9887 -4285 10233 -4251
rect 10267 -4285 10305 -4251
rect 10339 -4285 10491 -4251
rect 10525 -4285 10563 -4251
rect 10597 -4285 10749 -4251
rect 10783 -4285 10821 -4251
rect 10855 -4285 11007 -4251
rect 11041 -4285 11079 -4251
rect 11113 -4285 11459 -4251
rect 11493 -4285 11531 -4251
rect 11565 -4285 11717 -4251
rect 11751 -4285 11789 -4251
rect 11823 -4285 11975 -4251
rect 12009 -4285 12047 -4251
rect 12081 -4285 12427 -4251
rect 12461 -4285 12499 -4251
rect 12533 -4285 12685 -4251
rect 12719 -4285 12757 -4251
rect 12791 -4285 12943 -4251
rect 12977 -4285 13015 -4251
rect 13049 -4285 13201 -4251
rect 13235 -4285 13273 -4251
rect 13307 -4285 13653 -4251
rect 13687 -4285 13725 -4251
rect 13759 -4264 13932 -4251
rect 13966 -4245 14344 -4230
rect 14491 -4051 14537 -4004
rect 14491 -4085 14497 -4051
rect 14531 -4085 14537 -4051
rect 14491 -4123 14537 -4085
rect 14491 -4157 14497 -4123
rect 14531 -4157 14537 -4123
rect 14491 -4245 14537 -4157
rect 14749 -4051 14795 -4004
rect 14749 -4085 14755 -4051
rect 14789 -4085 14795 -4051
rect 14749 -4123 14795 -4085
rect 14749 -4157 14755 -4123
rect 14789 -4157 14795 -4123
rect 14749 -4245 14795 -4157
rect 15007 -4051 15053 -4004
rect 15007 -4085 15013 -4051
rect 15047 -4085 15053 -4051
rect 15007 -4123 15053 -4085
rect 15007 -4157 15013 -4123
rect 15047 -4157 15053 -4123
rect 15007 -4245 15053 -4157
rect 15265 -4051 15311 -4004
rect 15265 -4085 15271 -4051
rect 15305 -4085 15311 -4051
rect 15265 -4123 15311 -4085
rect 15265 -4157 15271 -4123
rect 15305 -4157 15311 -4123
rect 15265 -4245 15311 -4157
rect 15523 -4051 15569 -4004
rect 15523 -4085 15529 -4051
rect 15563 -4085 15569 -4051
rect 15523 -4123 15569 -4085
rect 15523 -4157 15529 -4123
rect 15563 -4157 15569 -4123
rect 15523 -4245 15569 -4157
rect 15717 -4051 15763 -4004
rect 15717 -4085 15723 -4051
rect 15757 -4085 15763 -4051
rect 15717 -4123 15763 -4085
rect 15717 -4157 15723 -4123
rect 15757 -4157 15763 -4123
rect 15717 -4245 15763 -4157
rect 15975 -4051 16021 -4004
rect 15975 -4085 15981 -4051
rect 16015 -4085 16021 -4051
rect 15975 -4123 16021 -4085
rect 15975 -4157 15981 -4123
rect 16015 -4157 16021 -4123
rect 15975 -4245 16021 -4157
rect 16233 -4051 16279 -4004
rect 16233 -4085 16239 -4051
rect 16273 -4085 16279 -4051
rect 16233 -4123 16279 -4085
rect 16233 -4157 16239 -4123
rect 16273 -4157 16279 -4123
rect 16233 -4245 16279 -4157
rect 16491 -4051 16537 -4004
rect 16491 -4085 16497 -4051
rect 16531 -4085 16537 -4051
rect 16491 -4123 16537 -4085
rect 16491 -4157 16497 -4123
rect 16531 -4157 16537 -4123
rect 16491 -4245 16537 -4157
rect 16685 -4051 16731 -4004
rect 16685 -4085 16691 -4051
rect 16725 -4085 16731 -4051
rect 16685 -4123 16731 -4085
rect 16685 -4157 16691 -4123
rect 16725 -4157 16731 -4123
rect 16685 -4245 16731 -4157
rect 16943 -4051 16989 -4004
rect 16943 -4085 16949 -4051
rect 16983 -4085 16989 -4051
rect 16943 -4123 16989 -4085
rect 16943 -4157 16949 -4123
rect 16983 -4157 16989 -4123
rect 16943 -4245 16989 -4157
rect 17201 -4051 17247 -4004
rect 17201 -4085 17207 -4051
rect 17241 -4085 17247 -4051
rect 17201 -4123 17247 -4085
rect 17201 -4157 17207 -4123
rect 17241 -4157 17247 -4123
rect 17201 -4245 17247 -4157
rect 17459 -4051 17505 -4004
rect 17459 -4085 17465 -4051
rect 17499 -4085 17505 -4051
rect 17459 -4123 17505 -4085
rect 17459 -4157 17465 -4123
rect 17499 -4157 17505 -4123
rect 17459 -4245 17505 -4157
rect 17717 -4051 17763 -4004
rect 17717 -4085 17723 -4051
rect 17757 -4085 17763 -4051
rect 17717 -4123 17763 -4085
rect 17717 -4157 17723 -4123
rect 17757 -4157 17763 -4123
rect 17717 -4245 17763 -4157
rect 17911 -4014 18347 -3976
rect 17911 -4048 18290 -4014
rect 18324 -4048 18347 -4014
rect 17911 -4051 18347 -4048
rect 17911 -4085 17917 -4051
rect 17951 -4085 18175 -4051
rect 18209 -4085 18347 -4051
rect 17911 -4086 18347 -4085
rect 17911 -4120 18290 -4086
rect 18324 -4120 18347 -4086
rect 17911 -4123 18347 -4120
rect 17911 -4157 17917 -4123
rect 17951 -4157 18175 -4123
rect 18209 -4157 18347 -4123
rect 17911 -4158 18347 -4157
rect 17911 -4192 18290 -4158
rect 18324 -4192 18347 -4158
rect 17911 -4230 18347 -4192
rect 17911 -4245 18290 -4230
rect 13966 -4251 18290 -4245
rect 13966 -4264 14139 -4251
rect 13759 -4285 14139 -4264
rect 14173 -4285 14211 -4251
rect 14245 -4285 14590 -4251
rect 14624 -4285 14662 -4251
rect 14696 -4285 14848 -4251
rect 14882 -4285 14920 -4251
rect 14954 -4285 15106 -4251
rect 15140 -4285 15178 -4251
rect 15212 -4285 15364 -4251
rect 15398 -4285 15436 -4251
rect 15470 -4285 15816 -4251
rect 15850 -4285 15888 -4251
rect 15922 -4285 16074 -4251
rect 16108 -4285 16146 -4251
rect 16180 -4285 16332 -4251
rect 16366 -4285 16404 -4251
rect 16438 -4285 16784 -4251
rect 16818 -4285 16856 -4251
rect 16890 -4285 17042 -4251
rect 17076 -4285 17114 -4251
rect 17148 -4285 17300 -4251
rect 17334 -4285 17372 -4251
rect 17406 -4285 17558 -4251
rect 17592 -4285 17630 -4251
rect 17664 -4285 18010 -4251
rect 18044 -4285 18082 -4251
rect 18116 -4264 18290 -4251
rect 18324 -4245 18347 -4230
rect 18324 -4264 18349 -4245
rect 18116 -4285 18349 -4264
rect 831 -4302 18349 -4285
rect 831 -4336 856 -4302
rect 890 -4336 5214 -4302
rect 5248 -4336 9573 -4302
rect 9607 -4336 13932 -4302
rect 13966 -4336 18290 -4302
rect 18324 -4336 18349 -4302
rect 831 -4365 18349 -4336
rect 831 -4399 930 -4365
rect 964 -4399 1002 -4365
rect 1036 -4399 1074 -4365
rect 1108 -4399 1146 -4365
rect 1180 -4399 1218 -4365
rect 1252 -4399 1290 -4365
rect 1324 -4399 1362 -4365
rect 1396 -4399 1434 -4365
rect 1468 -4399 1506 -4365
rect 1540 -4399 1578 -4365
rect 1612 -4399 1650 -4365
rect 1684 -4399 1722 -4365
rect 1756 -4399 1794 -4365
rect 1828 -4399 1866 -4365
rect 1900 -4399 1938 -4365
rect 1972 -4399 2010 -4365
rect 2044 -4399 2082 -4365
rect 2116 -4399 2154 -4365
rect 2188 -4399 2226 -4365
rect 2260 -4399 2298 -4365
rect 2332 -4399 2370 -4365
rect 2404 -4399 2442 -4365
rect 2476 -4399 2514 -4365
rect 2548 -4399 2586 -4365
rect 2620 -4399 2658 -4365
rect 2692 -4399 2730 -4365
rect 2764 -4399 2802 -4365
rect 2836 -4399 2874 -4365
rect 2908 -4399 2946 -4365
rect 2980 -4399 3018 -4365
rect 3052 -4399 3090 -4365
rect 3124 -4399 3162 -4365
rect 3196 -4399 3234 -4365
rect 3268 -4399 3306 -4365
rect 3340 -4399 3378 -4365
rect 3412 -4399 3450 -4365
rect 3484 -4399 3522 -4365
rect 3556 -4399 3594 -4365
rect 3628 -4399 3666 -4365
rect 3700 -4399 3738 -4365
rect 3772 -4399 3810 -4365
rect 3844 -4399 3882 -4365
rect 3916 -4399 3954 -4365
rect 3988 -4399 4026 -4365
rect 4060 -4399 4098 -4365
rect 4132 -4399 4170 -4365
rect 4204 -4399 4242 -4365
rect 4276 -4399 4314 -4365
rect 4348 -4399 4386 -4365
rect 4420 -4399 4458 -4365
rect 4492 -4399 4530 -4365
rect 4564 -4399 4602 -4365
rect 4636 -4399 4674 -4365
rect 4708 -4399 4746 -4365
rect 4780 -4399 4818 -4365
rect 4852 -4399 4890 -4365
rect 4924 -4399 4962 -4365
rect 4996 -4399 5034 -4365
rect 5068 -4399 5106 -4365
rect 5140 -4399 5323 -4365
rect 5357 -4399 5395 -4365
rect 5429 -4399 5467 -4365
rect 5501 -4399 5539 -4365
rect 5573 -4399 5611 -4365
rect 5645 -4399 5683 -4365
rect 5717 -4399 5755 -4365
rect 5789 -4399 5827 -4365
rect 5861 -4399 5899 -4365
rect 5933 -4399 5971 -4365
rect 6005 -4399 6043 -4365
rect 6077 -4399 6115 -4365
rect 6149 -4399 6187 -4365
rect 6221 -4399 6259 -4365
rect 6293 -4399 6331 -4365
rect 6365 -4399 6403 -4365
rect 6437 -4399 6475 -4365
rect 6509 -4399 6547 -4365
rect 6581 -4399 6619 -4365
rect 6653 -4399 6691 -4365
rect 6725 -4399 6763 -4365
rect 6797 -4399 6835 -4365
rect 6869 -4399 6907 -4365
rect 6941 -4399 6979 -4365
rect 7013 -4399 7051 -4365
rect 7085 -4399 7123 -4365
rect 7157 -4399 7195 -4365
rect 7229 -4399 7267 -4365
rect 7301 -4399 7339 -4365
rect 7373 -4399 7411 -4365
rect 7445 -4399 7483 -4365
rect 7517 -4399 7555 -4365
rect 7589 -4399 7627 -4365
rect 7661 -4399 7699 -4365
rect 7733 -4399 7771 -4365
rect 7805 -4399 7843 -4365
rect 7877 -4399 7915 -4365
rect 7949 -4399 7987 -4365
rect 8021 -4399 8059 -4365
rect 8093 -4399 8131 -4365
rect 8165 -4399 8203 -4365
rect 8237 -4399 8275 -4365
rect 8309 -4399 8347 -4365
rect 8381 -4399 8419 -4365
rect 8453 -4399 8491 -4365
rect 8525 -4399 8563 -4365
rect 8597 -4399 8635 -4365
rect 8669 -4399 8707 -4365
rect 8741 -4399 8779 -4365
rect 8813 -4399 8851 -4365
rect 8885 -4399 8923 -4365
rect 8957 -4399 8995 -4365
rect 9029 -4399 9067 -4365
rect 9101 -4399 9139 -4365
rect 9173 -4399 9211 -4365
rect 9245 -4399 9283 -4365
rect 9317 -4399 9355 -4365
rect 9389 -4399 9427 -4365
rect 9461 -4399 9499 -4365
rect 9533 -4399 9647 -4365
rect 9681 -4399 9719 -4365
rect 9753 -4399 9791 -4365
rect 9825 -4399 9863 -4365
rect 9897 -4399 9935 -4365
rect 9969 -4399 10007 -4365
rect 10041 -4399 10079 -4365
rect 10113 -4399 10151 -4365
rect 10185 -4399 10223 -4365
rect 10257 -4399 10295 -4365
rect 10329 -4399 10367 -4365
rect 10401 -4399 10439 -4365
rect 10473 -4399 10511 -4365
rect 10545 -4399 10583 -4365
rect 10617 -4399 10655 -4365
rect 10689 -4399 10727 -4365
rect 10761 -4399 10799 -4365
rect 10833 -4399 10871 -4365
rect 10905 -4399 10943 -4365
rect 10977 -4399 11015 -4365
rect 11049 -4399 11087 -4365
rect 11121 -4399 11159 -4365
rect 11193 -4399 11231 -4365
rect 11265 -4399 11303 -4365
rect 11337 -4399 11375 -4365
rect 11409 -4399 11447 -4365
rect 11481 -4399 11519 -4365
rect 11553 -4399 11591 -4365
rect 11625 -4399 11663 -4365
rect 11697 -4399 11735 -4365
rect 11769 -4399 11807 -4365
rect 11841 -4399 11879 -4365
rect 11913 -4399 11951 -4365
rect 11985 -4399 12023 -4365
rect 12057 -4399 12095 -4365
rect 12129 -4399 12167 -4365
rect 12201 -4399 12239 -4365
rect 12273 -4399 12311 -4365
rect 12345 -4399 12383 -4365
rect 12417 -4399 12455 -4365
rect 12489 -4399 12527 -4365
rect 12561 -4399 12599 -4365
rect 12633 -4399 12671 -4365
rect 12705 -4399 12743 -4365
rect 12777 -4399 12815 -4365
rect 12849 -4399 12887 -4365
rect 12921 -4399 12959 -4365
rect 12993 -4399 13031 -4365
rect 13065 -4399 13103 -4365
rect 13137 -4399 13175 -4365
rect 13209 -4399 13247 -4365
rect 13281 -4399 13319 -4365
rect 13353 -4399 13391 -4365
rect 13425 -4399 13463 -4365
rect 13497 -4399 13535 -4365
rect 13569 -4399 13607 -4365
rect 13641 -4399 13679 -4365
rect 13713 -4399 13751 -4365
rect 13785 -4399 13823 -4365
rect 13857 -4399 14040 -4365
rect 14074 -4399 14112 -4365
rect 14146 -4399 14184 -4365
rect 14218 -4399 14256 -4365
rect 14290 -4399 14328 -4365
rect 14362 -4399 14400 -4365
rect 14434 -4399 14472 -4365
rect 14506 -4399 14544 -4365
rect 14578 -4399 14616 -4365
rect 14650 -4399 14688 -4365
rect 14722 -4399 14760 -4365
rect 14794 -4399 14832 -4365
rect 14866 -4399 14904 -4365
rect 14938 -4399 14976 -4365
rect 15010 -4399 15048 -4365
rect 15082 -4399 15120 -4365
rect 15154 -4399 15192 -4365
rect 15226 -4399 15264 -4365
rect 15298 -4399 15336 -4365
rect 15370 -4399 15408 -4365
rect 15442 -4399 15480 -4365
rect 15514 -4399 15552 -4365
rect 15586 -4399 15624 -4365
rect 15658 -4399 15696 -4365
rect 15730 -4399 15768 -4365
rect 15802 -4399 15840 -4365
rect 15874 -4399 15912 -4365
rect 15946 -4399 15984 -4365
rect 16018 -4399 16056 -4365
rect 16090 -4399 16128 -4365
rect 16162 -4399 16200 -4365
rect 16234 -4399 16272 -4365
rect 16306 -4399 16344 -4365
rect 16378 -4399 16416 -4365
rect 16450 -4399 16488 -4365
rect 16522 -4399 16560 -4365
rect 16594 -4399 16632 -4365
rect 16666 -4399 16704 -4365
rect 16738 -4399 16776 -4365
rect 16810 -4399 16848 -4365
rect 16882 -4399 16920 -4365
rect 16954 -4399 16992 -4365
rect 17026 -4399 17064 -4365
rect 17098 -4399 17136 -4365
rect 17170 -4399 17208 -4365
rect 17242 -4399 17280 -4365
rect 17314 -4399 17352 -4365
rect 17386 -4399 17424 -4365
rect 17458 -4399 17496 -4365
rect 17530 -4399 17568 -4365
rect 17602 -4399 17640 -4365
rect 17674 -4399 17712 -4365
rect 17746 -4399 17784 -4365
rect 17818 -4399 17856 -4365
rect 17890 -4399 17928 -4365
rect 17962 -4399 18000 -4365
rect 18034 -4399 18072 -4365
rect 18106 -4399 18144 -4365
rect 18178 -4399 18216 -4365
rect 18250 -4399 18349 -4365
rect 831 -4428 18349 -4399
rect 831 -4462 856 -4428
rect 890 -4462 5214 -4428
rect 5248 -4462 9573 -4428
rect 9607 -4462 13932 -4428
rect 13966 -4462 18290 -4428
rect 18324 -4462 18349 -4428
rect 831 -4479 18349 -4462
rect 831 -4500 1064 -4479
rect 831 -4519 856 -4500
rect 833 -4534 856 -4519
rect 890 -4513 1064 -4500
rect 1098 -4513 1136 -4479
rect 1170 -4513 1516 -4479
rect 1550 -4513 1588 -4479
rect 1622 -4513 1774 -4479
rect 1808 -4513 1846 -4479
rect 1880 -4513 2032 -4479
rect 2066 -4513 2104 -4479
rect 2138 -4513 2290 -4479
rect 2324 -4513 2362 -4479
rect 2396 -4513 2742 -4479
rect 2776 -4513 2814 -4479
rect 2848 -4513 3000 -4479
rect 3034 -4513 3072 -4479
rect 3106 -4513 3258 -4479
rect 3292 -4513 3330 -4479
rect 3364 -4513 3710 -4479
rect 3744 -4513 3782 -4479
rect 3816 -4513 3968 -4479
rect 4002 -4513 4040 -4479
rect 4074 -4513 4226 -4479
rect 4260 -4513 4298 -4479
rect 4332 -4513 4484 -4479
rect 4518 -4513 4556 -4479
rect 4590 -4513 4935 -4479
rect 4969 -4513 5007 -4479
rect 5041 -4500 5421 -4479
rect 5041 -4513 5214 -4500
rect 890 -4519 5214 -4513
rect 890 -4534 1269 -4519
rect 833 -4572 1269 -4534
rect 833 -4606 856 -4572
rect 890 -4606 1269 -4572
rect 833 -4607 1269 -4606
rect 833 -4641 971 -4607
rect 1005 -4641 1229 -4607
rect 1263 -4641 1269 -4607
rect 833 -4644 1269 -4641
rect 833 -4678 856 -4644
rect 890 -4678 1269 -4644
rect 833 -4679 1269 -4678
rect 833 -4713 971 -4679
rect 1005 -4713 1229 -4679
rect 1263 -4713 1269 -4679
rect 833 -4716 1269 -4713
rect 833 -4750 856 -4716
rect 890 -4750 1269 -4716
rect 833 -4788 1269 -4750
rect 1417 -4607 1463 -4519
rect 1417 -4641 1423 -4607
rect 1457 -4641 1463 -4607
rect 1417 -4679 1463 -4641
rect 1417 -4713 1423 -4679
rect 1457 -4713 1463 -4679
rect 1417 -4760 1463 -4713
rect 1675 -4607 1721 -4519
rect 1675 -4641 1681 -4607
rect 1715 -4641 1721 -4607
rect 1675 -4679 1721 -4641
rect 1675 -4713 1681 -4679
rect 1715 -4713 1721 -4679
rect 1675 -4760 1721 -4713
rect 1933 -4607 1979 -4519
rect 1933 -4641 1939 -4607
rect 1973 -4641 1979 -4607
rect 1933 -4679 1979 -4641
rect 1933 -4713 1939 -4679
rect 1973 -4713 1979 -4679
rect 1933 -4760 1979 -4713
rect 2191 -4607 2237 -4519
rect 2191 -4641 2197 -4607
rect 2231 -4641 2237 -4607
rect 2191 -4679 2237 -4641
rect 2191 -4713 2197 -4679
rect 2231 -4713 2237 -4679
rect 2191 -4760 2237 -4713
rect 2449 -4607 2495 -4519
rect 2449 -4641 2455 -4607
rect 2489 -4641 2495 -4607
rect 2449 -4679 2495 -4641
rect 2449 -4713 2455 -4679
rect 2489 -4713 2495 -4679
rect 2449 -4760 2495 -4713
rect 2643 -4607 2689 -4519
rect 2643 -4641 2649 -4607
rect 2683 -4641 2689 -4607
rect 2643 -4679 2689 -4641
rect 2643 -4713 2649 -4679
rect 2683 -4713 2689 -4679
rect 2643 -4760 2689 -4713
rect 2901 -4607 2947 -4519
rect 2901 -4641 2907 -4607
rect 2941 -4641 2947 -4607
rect 2901 -4679 2947 -4641
rect 2901 -4713 2907 -4679
rect 2941 -4713 2947 -4679
rect 2901 -4760 2947 -4713
rect 3159 -4607 3205 -4519
rect 3159 -4641 3165 -4607
rect 3199 -4641 3205 -4607
rect 3159 -4679 3205 -4641
rect 3159 -4713 3165 -4679
rect 3199 -4713 3205 -4679
rect 3159 -4760 3205 -4713
rect 3417 -4607 3463 -4519
rect 3417 -4641 3423 -4607
rect 3457 -4641 3463 -4607
rect 3417 -4679 3463 -4641
rect 3417 -4713 3423 -4679
rect 3457 -4713 3463 -4679
rect 3417 -4760 3463 -4713
rect 3611 -4607 3657 -4519
rect 3611 -4641 3617 -4607
rect 3651 -4641 3657 -4607
rect 3611 -4679 3657 -4641
rect 3611 -4713 3617 -4679
rect 3651 -4713 3657 -4679
rect 3611 -4760 3657 -4713
rect 3869 -4607 3915 -4519
rect 3869 -4641 3875 -4607
rect 3909 -4641 3915 -4607
rect 3869 -4679 3915 -4641
rect 3869 -4713 3875 -4679
rect 3909 -4713 3915 -4679
rect 3869 -4760 3915 -4713
rect 4127 -4607 4173 -4519
rect 4127 -4641 4133 -4607
rect 4167 -4641 4173 -4607
rect 4127 -4679 4173 -4641
rect 4127 -4713 4133 -4679
rect 4167 -4713 4173 -4679
rect 4127 -4760 4173 -4713
rect 4385 -4607 4431 -4519
rect 4385 -4641 4391 -4607
rect 4425 -4641 4431 -4607
rect 4385 -4679 4431 -4641
rect 4385 -4713 4391 -4679
rect 4425 -4713 4431 -4679
rect 4385 -4760 4431 -4713
rect 4643 -4607 4689 -4519
rect 4643 -4641 4649 -4607
rect 4683 -4641 4689 -4607
rect 4643 -4679 4689 -4641
rect 4643 -4713 4649 -4679
rect 4683 -4713 4689 -4679
rect 4643 -4760 4689 -4713
rect 4836 -4534 5214 -4519
rect 5248 -4513 5421 -4500
rect 5455 -4513 5493 -4479
rect 5527 -4513 5873 -4479
rect 5907 -4513 5945 -4479
rect 5979 -4513 6131 -4479
rect 6165 -4513 6203 -4479
rect 6237 -4513 6389 -4479
rect 6423 -4513 6461 -4479
rect 6495 -4513 6647 -4479
rect 6681 -4513 6719 -4479
rect 6753 -4513 7099 -4479
rect 7133 -4513 7171 -4479
rect 7205 -4513 7357 -4479
rect 7391 -4513 7429 -4479
rect 7463 -4513 7615 -4479
rect 7649 -4513 7687 -4479
rect 7721 -4513 8067 -4479
rect 8101 -4513 8139 -4479
rect 8173 -4513 8325 -4479
rect 8359 -4513 8397 -4479
rect 8431 -4513 8583 -4479
rect 8617 -4513 8655 -4479
rect 8689 -4513 8841 -4479
rect 8875 -4513 8913 -4479
rect 8947 -4513 9293 -4479
rect 9327 -4513 9365 -4479
rect 9399 -4500 9781 -4479
rect 9399 -4513 9573 -4500
rect 5248 -4519 9573 -4513
rect 5248 -4534 5626 -4519
rect 4836 -4572 5626 -4534
rect 4836 -4606 5214 -4572
rect 5248 -4606 5626 -4572
rect 4836 -4607 5626 -4606
rect 4836 -4641 4842 -4607
rect 4876 -4641 5100 -4607
rect 5134 -4641 5328 -4607
rect 5362 -4641 5586 -4607
rect 5620 -4641 5626 -4607
rect 4836 -4644 5626 -4641
rect 4836 -4678 5214 -4644
rect 5248 -4678 5626 -4644
rect 4836 -4679 5626 -4678
rect 4836 -4713 4842 -4679
rect 4876 -4713 5100 -4679
rect 5134 -4713 5328 -4679
rect 5362 -4713 5586 -4679
rect 5620 -4713 5626 -4679
rect 4836 -4716 5626 -4713
rect 4836 -4750 5214 -4716
rect 5248 -4750 5626 -4716
rect 833 -4822 856 -4788
rect 890 -4822 1269 -4788
rect 833 -4860 1269 -4822
rect 833 -4894 856 -4860
rect 890 -4894 1269 -4860
rect 4836 -4788 5626 -4750
rect 5774 -4607 5820 -4519
rect 5774 -4641 5780 -4607
rect 5814 -4641 5820 -4607
rect 5774 -4679 5820 -4641
rect 5774 -4713 5780 -4679
rect 5814 -4713 5820 -4679
rect 5774 -4760 5820 -4713
rect 6032 -4607 6078 -4519
rect 6032 -4641 6038 -4607
rect 6072 -4641 6078 -4607
rect 6032 -4679 6078 -4641
rect 6032 -4713 6038 -4679
rect 6072 -4713 6078 -4679
rect 6032 -4760 6078 -4713
rect 6290 -4607 6336 -4519
rect 6290 -4641 6296 -4607
rect 6330 -4641 6336 -4607
rect 6290 -4679 6336 -4641
rect 6290 -4713 6296 -4679
rect 6330 -4713 6336 -4679
rect 6290 -4760 6336 -4713
rect 6548 -4607 6594 -4519
rect 6548 -4641 6554 -4607
rect 6588 -4641 6594 -4607
rect 6548 -4679 6594 -4641
rect 6548 -4713 6554 -4679
rect 6588 -4713 6594 -4679
rect 6548 -4760 6594 -4713
rect 6806 -4607 6852 -4519
rect 6806 -4641 6812 -4607
rect 6846 -4641 6852 -4607
rect 6806 -4679 6852 -4641
rect 6806 -4713 6812 -4679
rect 6846 -4713 6852 -4679
rect 6806 -4760 6852 -4713
rect 7000 -4607 7046 -4519
rect 7000 -4641 7006 -4607
rect 7040 -4641 7046 -4607
rect 7000 -4679 7046 -4641
rect 7000 -4713 7006 -4679
rect 7040 -4713 7046 -4679
rect 7000 -4760 7046 -4713
rect 7258 -4607 7304 -4519
rect 7258 -4641 7264 -4607
rect 7298 -4641 7304 -4607
rect 7258 -4679 7304 -4641
rect 7258 -4713 7264 -4679
rect 7298 -4713 7304 -4679
rect 7258 -4760 7304 -4713
rect 7516 -4607 7562 -4519
rect 7516 -4641 7522 -4607
rect 7556 -4641 7562 -4607
rect 7516 -4679 7562 -4641
rect 7516 -4713 7522 -4679
rect 7556 -4713 7562 -4679
rect 7516 -4760 7562 -4713
rect 7774 -4607 7820 -4519
rect 7774 -4641 7780 -4607
rect 7814 -4641 7820 -4607
rect 7774 -4679 7820 -4641
rect 7774 -4713 7780 -4679
rect 7814 -4713 7820 -4679
rect 7774 -4760 7820 -4713
rect 7968 -4607 8014 -4519
rect 7968 -4641 7974 -4607
rect 8008 -4641 8014 -4607
rect 7968 -4679 8014 -4641
rect 7968 -4713 7974 -4679
rect 8008 -4713 8014 -4679
rect 7968 -4760 8014 -4713
rect 8226 -4607 8272 -4519
rect 8226 -4641 8232 -4607
rect 8266 -4641 8272 -4607
rect 8226 -4679 8272 -4641
rect 8226 -4713 8232 -4679
rect 8266 -4713 8272 -4679
rect 8226 -4760 8272 -4713
rect 8484 -4607 8530 -4519
rect 8484 -4641 8490 -4607
rect 8524 -4641 8530 -4607
rect 8484 -4679 8530 -4641
rect 8484 -4713 8490 -4679
rect 8524 -4713 8530 -4679
rect 8484 -4760 8530 -4713
rect 8742 -4607 8788 -4519
rect 8742 -4641 8748 -4607
rect 8782 -4641 8788 -4607
rect 8742 -4679 8788 -4641
rect 8742 -4713 8748 -4679
rect 8782 -4713 8788 -4679
rect 8742 -4760 8788 -4713
rect 9000 -4607 9046 -4519
rect 9000 -4641 9006 -4607
rect 9040 -4641 9046 -4607
rect 9000 -4679 9046 -4641
rect 9000 -4713 9006 -4679
rect 9040 -4713 9046 -4679
rect 9000 -4760 9046 -4713
rect 9194 -4534 9573 -4519
rect 9607 -4513 9781 -4500
rect 9815 -4513 9853 -4479
rect 9887 -4513 10233 -4479
rect 10267 -4513 10305 -4479
rect 10339 -4513 10491 -4479
rect 10525 -4513 10563 -4479
rect 10597 -4513 10749 -4479
rect 10783 -4513 10821 -4479
rect 10855 -4513 11007 -4479
rect 11041 -4513 11079 -4479
rect 11113 -4513 11459 -4479
rect 11493 -4513 11531 -4479
rect 11565 -4513 11717 -4479
rect 11751 -4513 11789 -4479
rect 11823 -4513 11975 -4479
rect 12009 -4513 12047 -4479
rect 12081 -4513 12427 -4479
rect 12461 -4513 12499 -4479
rect 12533 -4513 12685 -4479
rect 12719 -4513 12757 -4479
rect 12791 -4513 12943 -4479
rect 12977 -4513 13015 -4479
rect 13049 -4513 13201 -4479
rect 13235 -4513 13273 -4479
rect 13307 -4513 13653 -4479
rect 13687 -4513 13725 -4479
rect 13759 -4500 14139 -4479
rect 13759 -4513 13932 -4500
rect 9607 -4519 13932 -4513
rect 9607 -4534 9986 -4519
rect 9194 -4572 9986 -4534
rect 9194 -4606 9573 -4572
rect 9607 -4606 9986 -4572
rect 9194 -4607 9986 -4606
rect 9194 -4641 9200 -4607
rect 9234 -4641 9458 -4607
rect 9492 -4641 9688 -4607
rect 9722 -4641 9946 -4607
rect 9980 -4641 9986 -4607
rect 9194 -4644 9986 -4641
rect 9194 -4678 9573 -4644
rect 9607 -4678 9986 -4644
rect 9194 -4679 9986 -4678
rect 9194 -4713 9200 -4679
rect 9234 -4713 9458 -4679
rect 9492 -4713 9688 -4679
rect 9722 -4713 9946 -4679
rect 9980 -4713 9986 -4679
rect 9194 -4716 9986 -4713
rect 9194 -4750 9573 -4716
rect 9607 -4750 9986 -4716
rect 4836 -4822 5214 -4788
rect 5248 -4822 5626 -4788
rect 4836 -4860 5626 -4822
rect 833 -4932 1269 -4894
rect 833 -4966 856 -4932
rect 890 -4966 1269 -4932
rect 2827 -4885 3023 -4877
rect 2827 -4937 2834 -4885
rect 2886 -4937 2898 -4885
rect 2950 -4937 2962 -4885
rect 3014 -4937 3023 -4885
rect 2827 -4947 3023 -4937
rect 3344 -4885 3540 -4877
rect 3344 -4937 3351 -4885
rect 3403 -4937 3415 -4885
rect 3467 -4937 3479 -4885
rect 3531 -4937 3540 -4885
rect 3344 -4947 3540 -4937
rect 4836 -4894 5214 -4860
rect 5248 -4894 5626 -4860
rect 9194 -4788 9986 -4750
rect 10134 -4607 10180 -4519
rect 10134 -4641 10140 -4607
rect 10174 -4641 10180 -4607
rect 10134 -4679 10180 -4641
rect 10134 -4713 10140 -4679
rect 10174 -4713 10180 -4679
rect 10134 -4760 10180 -4713
rect 10392 -4607 10438 -4519
rect 10392 -4641 10398 -4607
rect 10432 -4641 10438 -4607
rect 10392 -4679 10438 -4641
rect 10392 -4713 10398 -4679
rect 10432 -4713 10438 -4679
rect 10392 -4760 10438 -4713
rect 10650 -4607 10696 -4519
rect 10650 -4641 10656 -4607
rect 10690 -4641 10696 -4607
rect 10650 -4679 10696 -4641
rect 10650 -4713 10656 -4679
rect 10690 -4713 10696 -4679
rect 10650 -4760 10696 -4713
rect 10908 -4607 10954 -4519
rect 10908 -4641 10914 -4607
rect 10948 -4641 10954 -4607
rect 10908 -4679 10954 -4641
rect 10908 -4713 10914 -4679
rect 10948 -4713 10954 -4679
rect 10908 -4760 10954 -4713
rect 11166 -4607 11212 -4519
rect 11166 -4641 11172 -4607
rect 11206 -4641 11212 -4607
rect 11166 -4679 11212 -4641
rect 11166 -4713 11172 -4679
rect 11206 -4713 11212 -4679
rect 11166 -4760 11212 -4713
rect 11360 -4607 11406 -4519
rect 11360 -4641 11366 -4607
rect 11400 -4641 11406 -4607
rect 11360 -4679 11406 -4641
rect 11360 -4713 11366 -4679
rect 11400 -4713 11406 -4679
rect 11360 -4760 11406 -4713
rect 11618 -4607 11664 -4519
rect 11618 -4641 11624 -4607
rect 11658 -4641 11664 -4607
rect 11618 -4679 11664 -4641
rect 11618 -4713 11624 -4679
rect 11658 -4713 11664 -4679
rect 11618 -4760 11664 -4713
rect 11876 -4607 11922 -4519
rect 11876 -4641 11882 -4607
rect 11916 -4641 11922 -4607
rect 11876 -4679 11922 -4641
rect 11876 -4713 11882 -4679
rect 11916 -4713 11922 -4679
rect 11876 -4760 11922 -4713
rect 12134 -4607 12180 -4519
rect 12134 -4641 12140 -4607
rect 12174 -4641 12180 -4607
rect 12134 -4679 12180 -4641
rect 12134 -4713 12140 -4679
rect 12174 -4713 12180 -4679
rect 12134 -4760 12180 -4713
rect 12328 -4607 12374 -4519
rect 12328 -4641 12334 -4607
rect 12368 -4641 12374 -4607
rect 12328 -4679 12374 -4641
rect 12328 -4713 12334 -4679
rect 12368 -4713 12374 -4679
rect 12328 -4760 12374 -4713
rect 12586 -4607 12632 -4519
rect 12586 -4641 12592 -4607
rect 12626 -4641 12632 -4607
rect 12586 -4679 12632 -4641
rect 12586 -4713 12592 -4679
rect 12626 -4713 12632 -4679
rect 12586 -4760 12632 -4713
rect 12844 -4607 12890 -4519
rect 12844 -4641 12850 -4607
rect 12884 -4641 12890 -4607
rect 12844 -4679 12890 -4641
rect 12844 -4713 12850 -4679
rect 12884 -4713 12890 -4679
rect 12844 -4760 12890 -4713
rect 13102 -4607 13148 -4519
rect 13102 -4641 13108 -4607
rect 13142 -4641 13148 -4607
rect 13102 -4679 13148 -4641
rect 13102 -4713 13108 -4679
rect 13142 -4713 13148 -4679
rect 13102 -4760 13148 -4713
rect 13360 -4607 13406 -4519
rect 13360 -4641 13366 -4607
rect 13400 -4641 13406 -4607
rect 13360 -4679 13406 -4641
rect 13360 -4713 13366 -4679
rect 13400 -4713 13406 -4679
rect 13360 -4760 13406 -4713
rect 13554 -4534 13932 -4519
rect 13966 -4513 14139 -4500
rect 14173 -4513 14211 -4479
rect 14245 -4513 14590 -4479
rect 14624 -4513 14662 -4479
rect 14696 -4513 14848 -4479
rect 14882 -4513 14920 -4479
rect 14954 -4513 15106 -4479
rect 15140 -4513 15178 -4479
rect 15212 -4513 15364 -4479
rect 15398 -4513 15436 -4479
rect 15470 -4513 15816 -4479
rect 15850 -4513 15888 -4479
rect 15922 -4513 16074 -4479
rect 16108 -4513 16146 -4479
rect 16180 -4513 16332 -4479
rect 16366 -4513 16404 -4479
rect 16438 -4513 16784 -4479
rect 16818 -4513 16856 -4479
rect 16890 -4513 17042 -4479
rect 17076 -4513 17114 -4479
rect 17148 -4513 17300 -4479
rect 17334 -4513 17372 -4479
rect 17406 -4513 17558 -4479
rect 17592 -4513 17630 -4479
rect 17664 -4513 18010 -4479
rect 18044 -4513 18082 -4479
rect 18116 -4500 18349 -4479
rect 18116 -4513 18290 -4500
rect 13966 -4519 18290 -4513
rect 13966 -4534 14344 -4519
rect 13554 -4572 14344 -4534
rect 13554 -4606 13932 -4572
rect 13966 -4606 14344 -4572
rect 13554 -4607 14344 -4606
rect 13554 -4641 13560 -4607
rect 13594 -4641 13818 -4607
rect 13852 -4641 14046 -4607
rect 14080 -4641 14304 -4607
rect 14338 -4641 14344 -4607
rect 13554 -4644 14344 -4641
rect 13554 -4678 13932 -4644
rect 13966 -4678 14344 -4644
rect 13554 -4679 14344 -4678
rect 13554 -4713 13560 -4679
rect 13594 -4713 13818 -4679
rect 13852 -4713 14046 -4679
rect 14080 -4713 14304 -4679
rect 14338 -4713 14344 -4679
rect 13554 -4716 14344 -4713
rect 13554 -4750 13932 -4716
rect 13966 -4750 14344 -4716
rect 9194 -4822 9573 -4788
rect 9607 -4822 9986 -4788
rect 9194 -4860 9986 -4822
rect 4836 -4932 5626 -4894
rect 833 -5004 1269 -4966
rect 833 -5038 856 -5004
rect 890 -5038 1269 -5004
rect 833 -5076 1269 -5038
rect 833 -5110 856 -5076
rect 890 -5110 1269 -5076
rect 833 -5148 1269 -5110
rect 1339 -5054 1535 -5046
rect 1339 -5106 1348 -5054
rect 1400 -5106 1412 -5054
rect 1464 -5106 1476 -5054
rect 1528 -5106 1535 -5054
rect 1339 -5116 1535 -5106
rect 1856 -5054 2052 -5046
rect 1856 -5106 1865 -5054
rect 1917 -5106 1929 -5054
rect 1981 -5106 1993 -5054
rect 2045 -5106 2052 -5054
rect 1856 -5116 2052 -5106
rect 2373 -5054 2569 -5046
rect 2373 -5106 2382 -5054
rect 2434 -5106 2446 -5054
rect 2498 -5106 2510 -5054
rect 2562 -5106 2569 -5054
rect 2373 -5116 2569 -5106
rect 833 -5182 856 -5148
rect 890 -5182 1269 -5148
rect 833 -5220 1269 -5182
rect 833 -5254 856 -5220
rect 890 -5254 1269 -5220
rect 833 -5292 1269 -5254
rect 833 -5326 856 -5292
rect 890 -5326 1269 -5292
rect 833 -5364 1269 -5326
rect 833 -5398 856 -5364
rect 890 -5398 1269 -5364
rect 833 -5436 1269 -5398
rect 833 -5470 856 -5436
rect 890 -5470 1269 -5436
rect 833 -5508 1269 -5470
rect 833 -5542 856 -5508
rect 890 -5542 1269 -5508
rect 833 -5580 1269 -5542
rect 833 -5614 856 -5580
rect 890 -5597 1269 -5580
rect 890 -5614 971 -5597
rect 833 -5631 971 -5614
rect 1005 -5631 1229 -5597
rect 1263 -5631 1269 -5597
rect 833 -5652 1269 -5631
rect 833 -5686 856 -5652
rect 890 -5669 1269 -5652
rect 890 -5686 971 -5669
rect 833 -5703 971 -5686
rect 1005 -5703 1229 -5669
rect 1263 -5703 1269 -5669
rect 833 -5724 1269 -5703
rect 833 -5758 856 -5724
rect 890 -5758 1269 -5724
rect 1417 -5597 1463 -5116
rect 1598 -5386 1794 -5378
rect 1598 -5438 1607 -5386
rect 1659 -5438 1671 -5386
rect 1723 -5438 1735 -5386
rect 1787 -5438 1794 -5386
rect 1598 -5448 1794 -5438
rect 1417 -5631 1423 -5597
rect 1457 -5631 1463 -5597
rect 1417 -5669 1463 -5631
rect 1417 -5703 1423 -5669
rect 1457 -5703 1463 -5669
rect 1417 -5750 1463 -5703
rect 1675 -5597 1721 -5448
rect 1675 -5631 1681 -5597
rect 1715 -5631 1721 -5597
rect 1675 -5669 1721 -5631
rect 1675 -5703 1681 -5669
rect 1715 -5703 1721 -5669
rect 1675 -5750 1721 -5703
rect 1933 -5597 1979 -5116
rect 2116 -5386 2312 -5378
rect 2116 -5438 2125 -5386
rect 2177 -5438 2189 -5386
rect 2241 -5438 2253 -5386
rect 2305 -5438 2312 -5386
rect 2116 -5448 2312 -5438
rect 1933 -5631 1939 -5597
rect 1973 -5631 1979 -5597
rect 1933 -5669 1979 -5631
rect 1933 -5703 1939 -5669
rect 1973 -5703 1979 -5669
rect 1933 -5750 1979 -5703
rect 2191 -5597 2237 -5448
rect 2191 -5631 2197 -5597
rect 2231 -5631 2237 -5597
rect 2191 -5669 2237 -5631
rect 2191 -5703 2197 -5669
rect 2231 -5703 2237 -5669
rect 2191 -5750 2237 -5703
rect 2449 -5597 2495 -5116
rect 2570 -5217 2766 -5209
rect 2570 -5269 2577 -5217
rect 2629 -5269 2641 -5217
rect 2693 -5269 2705 -5217
rect 2757 -5269 2766 -5217
rect 2570 -5279 2766 -5269
rect 2449 -5631 2455 -5597
rect 2489 -5631 2495 -5597
rect 2449 -5669 2495 -5631
rect 2449 -5703 2455 -5669
rect 2489 -5703 2495 -5669
rect 2449 -5750 2495 -5703
rect 2643 -5597 2689 -5279
rect 2643 -5631 2649 -5597
rect 2683 -5631 2689 -5597
rect 2643 -5669 2689 -5631
rect 2643 -5703 2649 -5669
rect 2683 -5703 2689 -5669
rect 2643 -5750 2689 -5703
rect 2901 -5597 2947 -4947
rect 3087 -5217 3283 -5209
rect 3087 -5269 3094 -5217
rect 3146 -5269 3158 -5217
rect 3210 -5269 3222 -5217
rect 3274 -5269 3283 -5217
rect 3087 -5279 3283 -5269
rect 2901 -5631 2907 -5597
rect 2941 -5631 2947 -5597
rect 2901 -5669 2947 -5631
rect 2901 -5703 2907 -5669
rect 2941 -5703 2947 -5669
rect 2901 -5750 2947 -5703
rect 3159 -5597 3205 -5279
rect 3159 -5631 3165 -5597
rect 3199 -5631 3205 -5597
rect 3159 -5669 3205 -5631
rect 3159 -5703 3165 -5669
rect 3199 -5703 3205 -5669
rect 3159 -5750 3205 -5703
rect 3417 -5597 3463 -4947
rect 4836 -4966 5214 -4932
rect 5248 -4966 5626 -4932
rect 6922 -4885 7118 -4877
rect 6922 -4937 6931 -4885
rect 6983 -4937 6995 -4885
rect 7047 -4937 7059 -4885
rect 7111 -4937 7118 -4885
rect 6922 -4947 7118 -4937
rect 7440 -4885 7636 -4877
rect 7440 -4937 7449 -4885
rect 7501 -4937 7513 -4885
rect 7565 -4937 7577 -4885
rect 7629 -4937 7636 -4885
rect 7440 -4947 7636 -4937
rect 9194 -4894 9573 -4860
rect 9607 -4894 9986 -4860
rect 13554 -4788 14344 -4750
rect 14491 -4607 14537 -4519
rect 14491 -4641 14497 -4607
rect 14531 -4641 14537 -4607
rect 14491 -4679 14537 -4641
rect 14491 -4713 14497 -4679
rect 14531 -4713 14537 -4679
rect 14491 -4760 14537 -4713
rect 14749 -4607 14795 -4519
rect 14749 -4641 14755 -4607
rect 14789 -4641 14795 -4607
rect 14749 -4679 14795 -4641
rect 14749 -4713 14755 -4679
rect 14789 -4713 14795 -4679
rect 14749 -4760 14795 -4713
rect 15007 -4607 15053 -4519
rect 15007 -4641 15013 -4607
rect 15047 -4641 15053 -4607
rect 15007 -4679 15053 -4641
rect 15007 -4713 15013 -4679
rect 15047 -4713 15053 -4679
rect 15007 -4760 15053 -4713
rect 15265 -4607 15311 -4519
rect 15265 -4641 15271 -4607
rect 15305 -4641 15311 -4607
rect 15265 -4679 15311 -4641
rect 15265 -4713 15271 -4679
rect 15305 -4713 15311 -4679
rect 15265 -4760 15311 -4713
rect 15523 -4607 15569 -4519
rect 15523 -4641 15529 -4607
rect 15563 -4641 15569 -4607
rect 15523 -4679 15569 -4641
rect 15523 -4713 15529 -4679
rect 15563 -4713 15569 -4679
rect 15523 -4760 15569 -4713
rect 15717 -4607 15763 -4519
rect 15717 -4641 15723 -4607
rect 15757 -4641 15763 -4607
rect 15717 -4679 15763 -4641
rect 15717 -4713 15723 -4679
rect 15757 -4713 15763 -4679
rect 15717 -4760 15763 -4713
rect 15975 -4607 16021 -4519
rect 15975 -4641 15981 -4607
rect 16015 -4641 16021 -4607
rect 15975 -4679 16021 -4641
rect 15975 -4713 15981 -4679
rect 16015 -4713 16021 -4679
rect 15975 -4760 16021 -4713
rect 16233 -4607 16279 -4519
rect 16233 -4641 16239 -4607
rect 16273 -4641 16279 -4607
rect 16233 -4679 16279 -4641
rect 16233 -4713 16239 -4679
rect 16273 -4713 16279 -4679
rect 16233 -4760 16279 -4713
rect 16491 -4607 16537 -4519
rect 16491 -4641 16497 -4607
rect 16531 -4641 16537 -4607
rect 16491 -4679 16537 -4641
rect 16491 -4713 16497 -4679
rect 16531 -4713 16537 -4679
rect 16491 -4760 16537 -4713
rect 16685 -4607 16731 -4519
rect 16685 -4641 16691 -4607
rect 16725 -4641 16731 -4607
rect 16685 -4679 16731 -4641
rect 16685 -4713 16691 -4679
rect 16725 -4713 16731 -4679
rect 16685 -4760 16731 -4713
rect 16943 -4607 16989 -4519
rect 16943 -4641 16949 -4607
rect 16983 -4641 16989 -4607
rect 16943 -4679 16989 -4641
rect 16943 -4713 16949 -4679
rect 16983 -4713 16989 -4679
rect 16943 -4760 16989 -4713
rect 17201 -4607 17247 -4519
rect 17201 -4641 17207 -4607
rect 17241 -4641 17247 -4607
rect 17201 -4679 17247 -4641
rect 17201 -4713 17207 -4679
rect 17241 -4713 17247 -4679
rect 17201 -4760 17247 -4713
rect 17459 -4607 17505 -4519
rect 17459 -4641 17465 -4607
rect 17499 -4641 17505 -4607
rect 17459 -4679 17505 -4641
rect 17459 -4713 17465 -4679
rect 17499 -4713 17505 -4679
rect 17459 -4760 17505 -4713
rect 17717 -4607 17763 -4519
rect 17717 -4641 17723 -4607
rect 17757 -4641 17763 -4607
rect 17717 -4679 17763 -4641
rect 17717 -4713 17723 -4679
rect 17757 -4713 17763 -4679
rect 17717 -4760 17763 -4713
rect 17911 -4534 18290 -4519
rect 18324 -4519 18349 -4500
rect 18324 -4534 18347 -4519
rect 17911 -4572 18347 -4534
rect 17911 -4606 18290 -4572
rect 18324 -4606 18347 -4572
rect 17911 -4607 18347 -4606
rect 17911 -4641 17917 -4607
rect 17951 -4641 18175 -4607
rect 18209 -4641 18347 -4607
rect 17911 -4644 18347 -4641
rect 17911 -4678 18290 -4644
rect 18324 -4678 18347 -4644
rect 17911 -4679 18347 -4678
rect 17911 -4713 17917 -4679
rect 17951 -4713 18175 -4679
rect 18209 -4713 18347 -4679
rect 17911 -4716 18347 -4713
rect 17911 -4750 18290 -4716
rect 18324 -4750 18347 -4716
rect 13554 -4822 13932 -4788
rect 13966 -4822 14344 -4788
rect 13554 -4860 14344 -4822
rect 9194 -4932 9986 -4894
rect 4836 -5004 5626 -4966
rect 4836 -5038 5214 -5004
rect 5248 -5038 5626 -5004
rect 3534 -5054 3730 -5046
rect 3534 -5106 3543 -5054
rect 3595 -5106 3607 -5054
rect 3659 -5106 3671 -5054
rect 3723 -5106 3730 -5054
rect 3534 -5116 3730 -5106
rect 4051 -5054 4247 -5046
rect 4051 -5106 4060 -5054
rect 4112 -5106 4124 -5054
rect 4176 -5106 4188 -5054
rect 4240 -5106 4247 -5054
rect 4051 -5116 4247 -5106
rect 4566 -5054 4762 -5046
rect 4566 -5106 4575 -5054
rect 4627 -5106 4639 -5054
rect 4691 -5106 4703 -5054
rect 4755 -5106 4762 -5054
rect 4566 -5116 4762 -5106
rect 4836 -5076 5626 -5038
rect 4836 -5110 5214 -5076
rect 5248 -5110 5626 -5076
rect 3417 -5631 3423 -5597
rect 3457 -5631 3463 -5597
rect 3417 -5669 3463 -5631
rect 3417 -5703 3423 -5669
rect 3457 -5703 3463 -5669
rect 3417 -5750 3463 -5703
rect 3611 -5597 3657 -5116
rect 3793 -5386 3989 -5378
rect 3793 -5438 3802 -5386
rect 3854 -5438 3866 -5386
rect 3918 -5438 3930 -5386
rect 3982 -5438 3989 -5386
rect 3793 -5448 3989 -5438
rect 3611 -5631 3617 -5597
rect 3651 -5631 3657 -5597
rect 3611 -5669 3657 -5631
rect 3611 -5703 3617 -5669
rect 3651 -5703 3657 -5669
rect 3611 -5750 3657 -5703
rect 3869 -5597 3915 -5448
rect 3869 -5631 3875 -5597
rect 3909 -5631 3915 -5597
rect 3869 -5669 3915 -5631
rect 3869 -5703 3875 -5669
rect 3909 -5703 3915 -5669
rect 3869 -5750 3915 -5703
rect 4127 -5597 4173 -5116
rect 4310 -5386 4506 -5378
rect 4310 -5438 4319 -5386
rect 4371 -5438 4383 -5386
rect 4435 -5438 4447 -5386
rect 4499 -5438 4506 -5386
rect 4310 -5448 4506 -5438
rect 4127 -5631 4133 -5597
rect 4167 -5631 4173 -5597
rect 4127 -5669 4173 -5631
rect 4127 -5703 4133 -5669
rect 4167 -5703 4173 -5669
rect 4127 -5750 4173 -5703
rect 4385 -5597 4431 -5448
rect 4385 -5631 4391 -5597
rect 4425 -5631 4431 -5597
rect 4385 -5669 4431 -5631
rect 4385 -5703 4391 -5669
rect 4425 -5703 4431 -5669
rect 4385 -5750 4431 -5703
rect 4643 -5597 4689 -5116
rect 4643 -5631 4649 -5597
rect 4683 -5631 4689 -5597
rect 4643 -5669 4689 -5631
rect 4643 -5703 4649 -5669
rect 4683 -5703 4689 -5669
rect 4643 -5750 4689 -5703
rect 4836 -5148 5626 -5110
rect 5701 -5054 5897 -5046
rect 5701 -5106 5708 -5054
rect 5760 -5106 5772 -5054
rect 5824 -5106 5836 -5054
rect 5888 -5106 5897 -5054
rect 5701 -5116 5897 -5106
rect 6216 -5054 6412 -5046
rect 6216 -5106 6223 -5054
rect 6275 -5106 6287 -5054
rect 6339 -5106 6351 -5054
rect 6403 -5106 6412 -5054
rect 6216 -5116 6412 -5106
rect 6733 -5054 6929 -5046
rect 6733 -5106 6740 -5054
rect 6792 -5106 6804 -5054
rect 6856 -5106 6868 -5054
rect 6920 -5106 6929 -5054
rect 6733 -5116 6929 -5106
rect 4836 -5182 5214 -5148
rect 5248 -5182 5626 -5148
rect 4836 -5220 5626 -5182
rect 4836 -5254 5214 -5220
rect 5248 -5254 5626 -5220
rect 4836 -5292 5626 -5254
rect 4836 -5326 5214 -5292
rect 5248 -5326 5626 -5292
rect 4836 -5364 5626 -5326
rect 4836 -5398 5214 -5364
rect 5248 -5398 5626 -5364
rect 4836 -5436 5626 -5398
rect 4836 -5470 5214 -5436
rect 5248 -5470 5626 -5436
rect 4836 -5508 5626 -5470
rect 4836 -5542 5214 -5508
rect 5248 -5542 5626 -5508
rect 4836 -5580 5626 -5542
rect 4836 -5597 5214 -5580
rect 4836 -5631 4842 -5597
rect 4876 -5631 5100 -5597
rect 5134 -5614 5214 -5597
rect 5248 -5597 5626 -5580
rect 5248 -5614 5328 -5597
rect 5134 -5631 5328 -5614
rect 5362 -5631 5586 -5597
rect 5620 -5631 5626 -5597
rect 4836 -5652 5626 -5631
rect 4836 -5669 5214 -5652
rect 4836 -5703 4842 -5669
rect 4876 -5703 5100 -5669
rect 5134 -5686 5214 -5669
rect 5248 -5669 5626 -5652
rect 5248 -5686 5328 -5669
rect 5134 -5703 5328 -5686
rect 5362 -5703 5586 -5669
rect 5620 -5703 5626 -5669
rect 4836 -5724 5626 -5703
rect 833 -5796 1269 -5758
rect 4836 -5758 5214 -5724
rect 5248 -5758 5626 -5724
rect 5774 -5597 5820 -5116
rect 5957 -5386 6153 -5378
rect 5957 -5438 5964 -5386
rect 6016 -5438 6028 -5386
rect 6080 -5438 6092 -5386
rect 6144 -5438 6153 -5386
rect 5957 -5448 6153 -5438
rect 5774 -5631 5780 -5597
rect 5814 -5631 5820 -5597
rect 5774 -5669 5820 -5631
rect 5774 -5703 5780 -5669
rect 5814 -5703 5820 -5669
rect 5774 -5750 5820 -5703
rect 6032 -5597 6078 -5448
rect 6032 -5631 6038 -5597
rect 6072 -5631 6078 -5597
rect 6032 -5669 6078 -5631
rect 6032 -5703 6038 -5669
rect 6072 -5703 6078 -5669
rect 6032 -5750 6078 -5703
rect 6290 -5597 6336 -5116
rect 6474 -5386 6670 -5378
rect 6474 -5438 6481 -5386
rect 6533 -5438 6545 -5386
rect 6597 -5438 6609 -5386
rect 6661 -5438 6670 -5386
rect 6474 -5448 6670 -5438
rect 6290 -5631 6296 -5597
rect 6330 -5631 6336 -5597
rect 6290 -5669 6336 -5631
rect 6290 -5703 6296 -5669
rect 6330 -5703 6336 -5669
rect 6290 -5750 6336 -5703
rect 6548 -5597 6594 -5448
rect 6548 -5631 6554 -5597
rect 6588 -5631 6594 -5597
rect 6548 -5669 6594 -5631
rect 6548 -5703 6554 -5669
rect 6588 -5703 6594 -5669
rect 6548 -5750 6594 -5703
rect 6806 -5597 6852 -5116
rect 6806 -5631 6812 -5597
rect 6846 -5631 6852 -5597
rect 6806 -5669 6852 -5631
rect 6806 -5703 6812 -5669
rect 6846 -5703 6852 -5669
rect 6806 -5750 6852 -5703
rect 7000 -5597 7046 -4947
rect 7180 -5217 7376 -5209
rect 7180 -5269 7189 -5217
rect 7241 -5269 7253 -5217
rect 7305 -5269 7317 -5217
rect 7369 -5269 7376 -5217
rect 7180 -5279 7376 -5269
rect 7000 -5631 7006 -5597
rect 7040 -5631 7046 -5597
rect 7000 -5669 7046 -5631
rect 7000 -5703 7006 -5669
rect 7040 -5703 7046 -5669
rect 7000 -5750 7046 -5703
rect 7258 -5597 7304 -5279
rect 7258 -5631 7264 -5597
rect 7298 -5631 7304 -5597
rect 7258 -5669 7304 -5631
rect 7258 -5703 7264 -5669
rect 7298 -5703 7304 -5669
rect 7258 -5750 7304 -5703
rect 7516 -5597 7562 -4947
rect 9194 -4966 9573 -4932
rect 9607 -4966 9986 -4932
rect 11544 -4885 11740 -4877
rect 11544 -4937 11551 -4885
rect 11603 -4937 11615 -4885
rect 11667 -4937 11679 -4885
rect 11731 -4937 11740 -4885
rect 11544 -4947 11740 -4937
rect 12062 -4885 12258 -4877
rect 12062 -4937 12069 -4885
rect 12121 -4937 12133 -4885
rect 12185 -4937 12197 -4885
rect 12249 -4937 12258 -4885
rect 12062 -4947 12258 -4937
rect 13554 -4894 13932 -4860
rect 13966 -4894 14344 -4860
rect 17911 -4788 18347 -4750
rect 17911 -4822 18290 -4788
rect 18324 -4822 18347 -4788
rect 17911 -4860 18347 -4822
rect 13554 -4932 14344 -4894
rect 9194 -5004 9986 -4966
rect 9194 -5038 9573 -5004
rect 9607 -5038 9986 -5004
rect 7894 -5054 8090 -5046
rect 7894 -5106 7901 -5054
rect 7953 -5106 7965 -5054
rect 8017 -5106 8029 -5054
rect 8081 -5106 8090 -5054
rect 7894 -5116 8090 -5106
rect 8410 -5054 8606 -5046
rect 8410 -5106 8417 -5054
rect 8469 -5106 8481 -5054
rect 8533 -5106 8545 -5054
rect 8597 -5106 8606 -5054
rect 8410 -5116 8606 -5106
rect 8928 -5054 9124 -5046
rect 8928 -5106 8935 -5054
rect 8987 -5106 8999 -5054
rect 9051 -5106 9063 -5054
rect 9115 -5106 9124 -5054
rect 8928 -5116 9124 -5106
rect 9194 -5076 9986 -5038
rect 9194 -5110 9573 -5076
rect 9607 -5110 9986 -5076
rect 7697 -5217 7893 -5209
rect 7697 -5269 7706 -5217
rect 7758 -5269 7770 -5217
rect 7822 -5269 7834 -5217
rect 7886 -5269 7893 -5217
rect 7697 -5279 7893 -5269
rect 7516 -5631 7522 -5597
rect 7556 -5631 7562 -5597
rect 7516 -5669 7562 -5631
rect 7516 -5703 7522 -5669
rect 7556 -5703 7562 -5669
rect 7516 -5750 7562 -5703
rect 7774 -5597 7820 -5279
rect 7774 -5631 7780 -5597
rect 7814 -5631 7820 -5597
rect 7774 -5669 7820 -5631
rect 7774 -5703 7780 -5669
rect 7814 -5703 7820 -5669
rect 7774 -5750 7820 -5703
rect 7968 -5597 8014 -5116
rect 8151 -5386 8347 -5378
rect 8151 -5438 8158 -5386
rect 8210 -5438 8222 -5386
rect 8274 -5438 8286 -5386
rect 8338 -5438 8347 -5386
rect 8151 -5448 8347 -5438
rect 7968 -5631 7974 -5597
rect 8008 -5631 8014 -5597
rect 7968 -5669 8014 -5631
rect 7968 -5703 7974 -5669
rect 8008 -5703 8014 -5669
rect 7968 -5750 8014 -5703
rect 8226 -5597 8272 -5448
rect 8226 -5631 8232 -5597
rect 8266 -5631 8272 -5597
rect 8226 -5669 8272 -5631
rect 8226 -5703 8232 -5669
rect 8266 -5703 8272 -5669
rect 8226 -5750 8272 -5703
rect 8484 -5597 8530 -5116
rect 8668 -5386 8864 -5378
rect 8668 -5438 8675 -5386
rect 8727 -5438 8739 -5386
rect 8791 -5438 8803 -5386
rect 8855 -5438 8864 -5386
rect 8668 -5448 8864 -5438
rect 8484 -5631 8490 -5597
rect 8524 -5631 8530 -5597
rect 8484 -5669 8530 -5631
rect 8484 -5703 8490 -5669
rect 8524 -5703 8530 -5669
rect 8484 -5750 8530 -5703
rect 8742 -5597 8788 -5448
rect 8742 -5631 8748 -5597
rect 8782 -5631 8788 -5597
rect 8742 -5669 8788 -5631
rect 8742 -5703 8748 -5669
rect 8782 -5703 8788 -5669
rect 8742 -5750 8788 -5703
rect 9000 -5597 9046 -5116
rect 9000 -5631 9006 -5597
rect 9040 -5631 9046 -5597
rect 9000 -5669 9046 -5631
rect 9000 -5703 9006 -5669
rect 9040 -5703 9046 -5669
rect 9000 -5750 9046 -5703
rect 9194 -5148 9986 -5110
rect 10056 -5054 10252 -5046
rect 10056 -5106 10065 -5054
rect 10117 -5106 10129 -5054
rect 10181 -5106 10193 -5054
rect 10245 -5106 10252 -5054
rect 10056 -5116 10252 -5106
rect 10574 -5054 10770 -5046
rect 10574 -5106 10583 -5054
rect 10635 -5106 10647 -5054
rect 10699 -5106 10711 -5054
rect 10763 -5106 10770 -5054
rect 10574 -5116 10770 -5106
rect 11090 -5054 11286 -5046
rect 11090 -5106 11099 -5054
rect 11151 -5106 11163 -5054
rect 11215 -5106 11227 -5054
rect 11279 -5106 11286 -5054
rect 11090 -5116 11286 -5106
rect 9194 -5182 9573 -5148
rect 9607 -5182 9986 -5148
rect 9194 -5220 9986 -5182
rect 9194 -5254 9573 -5220
rect 9607 -5254 9986 -5220
rect 9194 -5292 9986 -5254
rect 9194 -5326 9573 -5292
rect 9607 -5326 9986 -5292
rect 9194 -5364 9986 -5326
rect 9194 -5398 9573 -5364
rect 9607 -5398 9986 -5364
rect 9194 -5436 9986 -5398
rect 9194 -5470 9573 -5436
rect 9607 -5470 9986 -5436
rect 9194 -5508 9986 -5470
rect 9194 -5542 9573 -5508
rect 9607 -5542 9986 -5508
rect 9194 -5580 9986 -5542
rect 9194 -5597 9573 -5580
rect 9194 -5631 9200 -5597
rect 9234 -5631 9458 -5597
rect 9492 -5614 9573 -5597
rect 9607 -5597 9986 -5580
rect 9607 -5614 9688 -5597
rect 9492 -5631 9688 -5614
rect 9722 -5631 9946 -5597
rect 9980 -5631 9986 -5597
rect 9194 -5652 9986 -5631
rect 9194 -5669 9573 -5652
rect 9194 -5703 9200 -5669
rect 9234 -5703 9458 -5669
rect 9492 -5686 9573 -5669
rect 9607 -5669 9986 -5652
rect 9607 -5686 9688 -5669
rect 9492 -5703 9688 -5686
rect 9722 -5703 9946 -5669
rect 9980 -5703 9986 -5669
rect 9194 -5724 9986 -5703
rect 833 -5830 856 -5796
rect 890 -5797 1269 -5796
rect 890 -5830 1064 -5797
rect 833 -5831 1064 -5830
rect 1098 -5831 1136 -5797
rect 1170 -5831 1269 -5797
rect 833 -5868 1269 -5831
rect 833 -5902 856 -5868
rect 890 -5902 1269 -5868
rect 833 -5940 1269 -5902
rect 833 -5974 856 -5940
rect 890 -5974 1269 -5940
rect 833 -6012 1269 -5974
rect 833 -6046 856 -6012
rect 890 -6046 1269 -6012
rect 833 -6084 1269 -6046
rect 1473 -5797 2439 -5791
rect 1473 -5831 1516 -5797
rect 1550 -5812 1588 -5797
rect 1622 -5812 1774 -5797
rect 1808 -5812 1846 -5797
rect 1880 -5812 2032 -5797
rect 2066 -5812 2104 -5797
rect 2138 -5812 2290 -5797
rect 2324 -5812 2362 -5797
rect 1473 -5864 1523 -5831
rect 1575 -5864 1587 -5812
rect 1639 -5864 1651 -5812
rect 1703 -5864 1719 -5812
rect 1771 -5831 1774 -5812
rect 1835 -5831 1846 -5812
rect 1771 -5864 1783 -5831
rect 1835 -5864 1847 -5831
rect 1899 -5864 2009 -5812
rect 2066 -5831 2073 -5812
rect 2061 -5864 2073 -5831
rect 2125 -5864 2137 -5831
rect 2189 -5864 2205 -5812
rect 2257 -5864 2269 -5812
rect 2324 -5831 2333 -5812
rect 2396 -5831 2439 -5797
rect 2321 -5864 2333 -5831
rect 2385 -5864 2439 -5831
rect 1473 -5990 2439 -5864
rect 1473 -6042 1523 -5990
rect 1575 -6042 1587 -5990
rect 1639 -6042 1651 -5990
rect 1703 -6042 1719 -5990
rect 1771 -6042 1783 -5990
rect 1835 -6042 1847 -5990
rect 1899 -6042 2009 -5990
rect 2061 -6042 2073 -5990
rect 2125 -6042 2137 -5990
rect 2189 -6042 2205 -5990
rect 2257 -6042 2269 -5990
rect 2321 -6042 2333 -5990
rect 2385 -6042 2439 -5990
rect 1473 -6061 2439 -6042
rect 2516 -5797 3590 -5791
rect 2516 -5831 2742 -5797
rect 2776 -5831 2814 -5797
rect 2848 -5831 3000 -5797
rect 3034 -5831 3072 -5797
rect 3106 -5831 3258 -5797
rect 3292 -5831 3330 -5797
rect 3364 -5831 3590 -5797
rect 2516 -5879 3590 -5831
rect 833 -6118 856 -6084
rect 890 -6118 1269 -6084
rect 2516 -6111 2577 -5879
rect 833 -6156 1269 -6118
rect 833 -6190 856 -6156
rect 890 -6159 1269 -6156
rect 890 -6190 1064 -6159
rect 833 -6193 1064 -6190
rect 1098 -6193 1136 -6159
rect 1170 -6193 1269 -6159
rect 833 -6228 1269 -6193
rect 1473 -6129 2577 -6111
rect 1473 -6159 1523 -6129
rect 1473 -6193 1516 -6159
rect 1575 -6181 1587 -6129
rect 1639 -6181 1651 -6129
rect 1703 -6181 1719 -6129
rect 1771 -6159 1783 -6129
rect 1835 -6159 1847 -6129
rect 1771 -6181 1774 -6159
rect 1835 -6181 1846 -6159
rect 1899 -6181 2009 -6129
rect 2061 -6159 2073 -6129
rect 2125 -6159 2137 -6129
rect 2066 -6181 2073 -6159
rect 2189 -6181 2205 -6129
rect 2257 -6181 2269 -6129
rect 2321 -6159 2333 -6129
rect 2385 -6159 2577 -6129
rect 2324 -6181 2333 -6159
rect 1550 -6193 1588 -6181
rect 1622 -6193 1774 -6181
rect 1808 -6193 1846 -6181
rect 1880 -6193 2032 -6181
rect 2066 -6193 2104 -6181
rect 2138 -6193 2290 -6181
rect 2324 -6193 2362 -6181
rect 2396 -6193 2577 -6159
rect 1473 -6199 2577 -6193
rect 2699 -5990 3407 -5973
rect 2699 -6042 2733 -5990
rect 2785 -6042 2797 -5990
rect 2849 -6042 2861 -5990
rect 2913 -6042 2929 -5990
rect 2981 -6042 2993 -5990
rect 3045 -6042 3057 -5990
rect 3109 -6042 3121 -5990
rect 3173 -6042 3189 -5990
rect 3241 -6042 3253 -5990
rect 3305 -6042 3317 -5990
rect 3369 -6042 3407 -5990
rect 2699 -6159 3407 -6042
rect 2699 -6193 2742 -6159
rect 2776 -6193 2814 -6159
rect 2848 -6193 3000 -6159
rect 3034 -6193 3072 -6159
rect 3106 -6193 3258 -6159
rect 3292 -6193 3330 -6159
rect 3364 -6193 3407 -6159
rect 2699 -6199 3407 -6193
rect 3529 -6111 3590 -5879
rect 3667 -5797 4633 -5791
rect 3667 -5831 3710 -5797
rect 3744 -5812 3782 -5797
rect 3816 -5812 3968 -5797
rect 4002 -5812 4040 -5797
rect 4074 -5812 4226 -5797
rect 4260 -5812 4298 -5797
rect 4332 -5812 4484 -5797
rect 4518 -5812 4556 -5797
rect 3773 -5831 3782 -5812
rect 3667 -5864 3721 -5831
rect 3773 -5864 3785 -5831
rect 3837 -5864 3849 -5812
rect 3901 -5864 3917 -5812
rect 4033 -5831 4040 -5812
rect 3969 -5864 3981 -5831
rect 4033 -5864 4045 -5831
rect 4097 -5864 4207 -5812
rect 4260 -5831 4271 -5812
rect 4332 -5831 4335 -5812
rect 4259 -5864 4271 -5831
rect 4323 -5864 4335 -5831
rect 4387 -5864 4403 -5812
rect 4455 -5864 4467 -5812
rect 4519 -5864 4531 -5812
rect 4590 -5831 4633 -5797
rect 4583 -5864 4633 -5831
rect 3667 -5990 4633 -5864
rect 3667 -6042 3721 -5990
rect 3773 -6042 3785 -5990
rect 3837 -6042 3849 -5990
rect 3901 -6042 3917 -5990
rect 3969 -6042 3981 -5990
rect 4033 -6042 4045 -5990
rect 4097 -6042 4207 -5990
rect 4259 -6042 4271 -5990
rect 4323 -6042 4335 -5990
rect 4387 -6042 4403 -5990
rect 4455 -6042 4467 -5990
rect 4519 -6042 4531 -5990
rect 4583 -6042 4633 -5990
rect 3667 -6061 4633 -6042
rect 4836 -5796 5626 -5758
rect 9194 -5758 9573 -5724
rect 9607 -5758 9986 -5724
rect 10134 -5597 10180 -5116
rect 10316 -5386 10512 -5378
rect 10316 -5438 10325 -5386
rect 10377 -5438 10389 -5386
rect 10441 -5438 10453 -5386
rect 10505 -5438 10512 -5386
rect 10316 -5448 10512 -5438
rect 10134 -5631 10140 -5597
rect 10174 -5631 10180 -5597
rect 10134 -5669 10180 -5631
rect 10134 -5703 10140 -5669
rect 10174 -5703 10180 -5669
rect 10134 -5750 10180 -5703
rect 10392 -5597 10438 -5448
rect 10392 -5631 10398 -5597
rect 10432 -5631 10438 -5597
rect 10392 -5669 10438 -5631
rect 10392 -5703 10398 -5669
rect 10432 -5703 10438 -5669
rect 10392 -5750 10438 -5703
rect 10650 -5597 10696 -5116
rect 10833 -5386 11029 -5378
rect 10833 -5438 10842 -5386
rect 10894 -5438 10906 -5386
rect 10958 -5438 10970 -5386
rect 11022 -5438 11029 -5386
rect 10833 -5448 11029 -5438
rect 10650 -5631 10656 -5597
rect 10690 -5631 10696 -5597
rect 10650 -5669 10696 -5631
rect 10650 -5703 10656 -5669
rect 10690 -5703 10696 -5669
rect 10650 -5750 10696 -5703
rect 10908 -5597 10954 -5448
rect 10908 -5631 10914 -5597
rect 10948 -5631 10954 -5597
rect 10908 -5669 10954 -5631
rect 10908 -5703 10914 -5669
rect 10948 -5703 10954 -5669
rect 10908 -5750 10954 -5703
rect 11166 -5597 11212 -5116
rect 11287 -5217 11483 -5209
rect 11287 -5269 11294 -5217
rect 11346 -5269 11358 -5217
rect 11410 -5269 11422 -5217
rect 11474 -5269 11483 -5217
rect 11287 -5279 11483 -5269
rect 11166 -5631 11172 -5597
rect 11206 -5631 11212 -5597
rect 11166 -5669 11212 -5631
rect 11166 -5703 11172 -5669
rect 11206 -5703 11212 -5669
rect 11166 -5750 11212 -5703
rect 11360 -5597 11406 -5279
rect 11360 -5631 11366 -5597
rect 11400 -5631 11406 -5597
rect 11360 -5669 11406 -5631
rect 11360 -5703 11366 -5669
rect 11400 -5703 11406 -5669
rect 11360 -5750 11406 -5703
rect 11618 -5597 11664 -4947
rect 11804 -5217 12000 -5209
rect 11804 -5269 11811 -5217
rect 11863 -5269 11875 -5217
rect 11927 -5269 11939 -5217
rect 11991 -5269 12000 -5217
rect 11804 -5279 12000 -5269
rect 11618 -5631 11624 -5597
rect 11658 -5631 11664 -5597
rect 11618 -5669 11664 -5631
rect 11618 -5703 11624 -5669
rect 11658 -5703 11664 -5669
rect 11618 -5750 11664 -5703
rect 11876 -5597 11922 -5279
rect 11876 -5631 11882 -5597
rect 11916 -5631 11922 -5597
rect 11876 -5669 11922 -5631
rect 11876 -5703 11882 -5669
rect 11916 -5703 11922 -5669
rect 11876 -5750 11922 -5703
rect 12134 -5597 12180 -4947
rect 13554 -4966 13932 -4932
rect 13966 -4966 14344 -4932
rect 15640 -4885 15836 -4877
rect 15640 -4937 15649 -4885
rect 15701 -4937 15713 -4885
rect 15765 -4937 15777 -4885
rect 15829 -4937 15836 -4885
rect 15640 -4947 15836 -4937
rect 16157 -4885 16353 -4877
rect 16157 -4937 16166 -4885
rect 16218 -4937 16230 -4885
rect 16282 -4937 16294 -4885
rect 16346 -4937 16353 -4885
rect 16157 -4947 16353 -4937
rect 17911 -4894 18290 -4860
rect 18324 -4894 18347 -4860
rect 17911 -4932 18347 -4894
rect 13554 -5004 14344 -4966
rect 13554 -5038 13932 -5004
rect 13966 -5038 14344 -5004
rect 12251 -5054 12447 -5046
rect 12251 -5106 12260 -5054
rect 12312 -5106 12324 -5054
rect 12376 -5106 12388 -5054
rect 12440 -5106 12447 -5054
rect 12251 -5116 12447 -5106
rect 12768 -5054 12964 -5046
rect 12768 -5106 12777 -5054
rect 12829 -5106 12841 -5054
rect 12893 -5106 12905 -5054
rect 12957 -5106 12964 -5054
rect 12768 -5116 12964 -5106
rect 13283 -5054 13479 -5046
rect 13283 -5106 13292 -5054
rect 13344 -5106 13356 -5054
rect 13408 -5106 13420 -5054
rect 13472 -5106 13479 -5054
rect 13283 -5116 13479 -5106
rect 13554 -5076 14344 -5038
rect 13554 -5110 13932 -5076
rect 13966 -5110 14344 -5076
rect 12134 -5631 12140 -5597
rect 12174 -5631 12180 -5597
rect 12134 -5669 12180 -5631
rect 12134 -5703 12140 -5669
rect 12174 -5703 12180 -5669
rect 12134 -5750 12180 -5703
rect 12328 -5597 12374 -5116
rect 12510 -5386 12706 -5378
rect 12510 -5438 12519 -5386
rect 12571 -5438 12583 -5386
rect 12635 -5438 12647 -5386
rect 12699 -5438 12706 -5386
rect 12510 -5448 12706 -5438
rect 12328 -5631 12334 -5597
rect 12368 -5631 12374 -5597
rect 12328 -5669 12374 -5631
rect 12328 -5703 12334 -5669
rect 12368 -5703 12374 -5669
rect 12328 -5750 12374 -5703
rect 12586 -5597 12632 -5448
rect 12586 -5631 12592 -5597
rect 12626 -5631 12632 -5597
rect 12586 -5669 12632 -5631
rect 12586 -5703 12592 -5669
rect 12626 -5703 12632 -5669
rect 12586 -5750 12632 -5703
rect 12844 -5597 12890 -5116
rect 13027 -5386 13223 -5378
rect 13027 -5438 13036 -5386
rect 13088 -5438 13100 -5386
rect 13152 -5438 13164 -5386
rect 13216 -5438 13223 -5386
rect 13027 -5448 13223 -5438
rect 12844 -5631 12850 -5597
rect 12884 -5631 12890 -5597
rect 12844 -5669 12890 -5631
rect 12844 -5703 12850 -5669
rect 12884 -5703 12890 -5669
rect 12844 -5750 12890 -5703
rect 13102 -5597 13148 -5448
rect 13102 -5631 13108 -5597
rect 13142 -5631 13148 -5597
rect 13102 -5669 13148 -5631
rect 13102 -5703 13108 -5669
rect 13142 -5703 13148 -5669
rect 13102 -5750 13148 -5703
rect 13360 -5597 13406 -5116
rect 13360 -5631 13366 -5597
rect 13400 -5631 13406 -5597
rect 13360 -5669 13406 -5631
rect 13360 -5703 13366 -5669
rect 13400 -5703 13406 -5669
rect 13360 -5750 13406 -5703
rect 13554 -5148 14344 -5110
rect 14418 -5054 14614 -5046
rect 14418 -5106 14425 -5054
rect 14477 -5106 14489 -5054
rect 14541 -5106 14553 -5054
rect 14605 -5106 14614 -5054
rect 14418 -5116 14614 -5106
rect 14933 -5054 15129 -5046
rect 14933 -5106 14940 -5054
rect 14992 -5106 15004 -5054
rect 15056 -5106 15068 -5054
rect 15120 -5106 15129 -5054
rect 14933 -5116 15129 -5106
rect 15450 -5054 15646 -5046
rect 15450 -5106 15457 -5054
rect 15509 -5106 15521 -5054
rect 15573 -5106 15585 -5054
rect 15637 -5106 15646 -5054
rect 15450 -5116 15646 -5106
rect 13554 -5182 13932 -5148
rect 13966 -5182 14344 -5148
rect 13554 -5220 14344 -5182
rect 13554 -5254 13932 -5220
rect 13966 -5254 14344 -5220
rect 13554 -5292 14344 -5254
rect 13554 -5326 13932 -5292
rect 13966 -5326 14344 -5292
rect 13554 -5364 14344 -5326
rect 13554 -5398 13932 -5364
rect 13966 -5398 14344 -5364
rect 13554 -5436 14344 -5398
rect 13554 -5470 13932 -5436
rect 13966 -5470 14344 -5436
rect 13554 -5508 14344 -5470
rect 13554 -5542 13932 -5508
rect 13966 -5542 14344 -5508
rect 13554 -5580 14344 -5542
rect 13554 -5597 13932 -5580
rect 13554 -5631 13560 -5597
rect 13594 -5631 13818 -5597
rect 13852 -5614 13932 -5597
rect 13966 -5597 14344 -5580
rect 13966 -5614 14046 -5597
rect 13852 -5631 14046 -5614
rect 14080 -5631 14304 -5597
rect 14338 -5631 14344 -5597
rect 13554 -5652 14344 -5631
rect 13554 -5669 13932 -5652
rect 13554 -5703 13560 -5669
rect 13594 -5703 13818 -5669
rect 13852 -5686 13932 -5669
rect 13966 -5669 14344 -5652
rect 13966 -5686 14046 -5669
rect 13852 -5703 14046 -5686
rect 14080 -5703 14304 -5669
rect 14338 -5703 14344 -5669
rect 13554 -5724 14344 -5703
rect 4836 -5797 5214 -5796
rect 4836 -5831 4935 -5797
rect 4969 -5831 5007 -5797
rect 5041 -5830 5214 -5797
rect 5248 -5797 5626 -5796
rect 5248 -5830 5421 -5797
rect 5041 -5831 5421 -5830
rect 5455 -5831 5493 -5797
rect 5527 -5831 5626 -5797
rect 4836 -5868 5626 -5831
rect 4836 -5902 5214 -5868
rect 5248 -5902 5626 -5868
rect 4836 -5940 5626 -5902
rect 4836 -5974 5214 -5940
rect 5248 -5974 5626 -5940
rect 4836 -6012 5626 -5974
rect 4836 -6046 5214 -6012
rect 5248 -6046 5626 -6012
rect 4836 -6084 5626 -6046
rect 5830 -5797 6796 -5791
rect 5830 -5831 5873 -5797
rect 5907 -5812 5945 -5797
rect 5979 -5812 6131 -5797
rect 6165 -5812 6203 -5797
rect 6237 -5812 6389 -5797
rect 6423 -5812 6461 -5797
rect 6495 -5812 6647 -5797
rect 6681 -5812 6719 -5797
rect 5830 -5864 5880 -5831
rect 5932 -5864 5944 -5812
rect 5996 -5864 6008 -5812
rect 6060 -5864 6076 -5812
rect 6128 -5831 6131 -5812
rect 6192 -5831 6203 -5812
rect 6128 -5864 6140 -5831
rect 6192 -5864 6204 -5831
rect 6256 -5864 6366 -5812
rect 6423 -5831 6430 -5812
rect 6418 -5864 6430 -5831
rect 6482 -5864 6494 -5831
rect 6546 -5864 6562 -5812
rect 6614 -5864 6626 -5812
rect 6681 -5831 6690 -5812
rect 6753 -5831 6796 -5797
rect 6678 -5864 6690 -5831
rect 6742 -5864 6796 -5831
rect 5830 -5990 6796 -5864
rect 5830 -6042 5880 -5990
rect 5932 -6042 5944 -5990
rect 5996 -6042 6008 -5990
rect 6060 -6042 6076 -5990
rect 6128 -6042 6140 -5990
rect 6192 -6042 6204 -5990
rect 6256 -6042 6366 -5990
rect 6418 -6042 6430 -5990
rect 6482 -6042 6494 -5990
rect 6546 -6042 6562 -5990
rect 6614 -6042 6626 -5990
rect 6678 -6042 6690 -5990
rect 6742 -6042 6796 -5990
rect 5830 -6061 6796 -6042
rect 6873 -5797 7947 -5791
rect 6873 -5831 7099 -5797
rect 7133 -5831 7171 -5797
rect 7205 -5831 7357 -5797
rect 7391 -5831 7429 -5797
rect 7463 -5831 7615 -5797
rect 7649 -5831 7687 -5797
rect 7721 -5831 7947 -5797
rect 6873 -5879 7947 -5831
rect 3529 -6129 4633 -6111
rect 3529 -6159 3721 -6129
rect 3773 -6159 3785 -6129
rect 3529 -6193 3710 -6159
rect 3773 -6181 3782 -6159
rect 3837 -6181 3849 -6129
rect 3901 -6181 3917 -6129
rect 3969 -6159 3981 -6129
rect 4033 -6159 4045 -6129
rect 4033 -6181 4040 -6159
rect 4097 -6181 4207 -6129
rect 4259 -6159 4271 -6129
rect 4323 -6159 4335 -6129
rect 4260 -6181 4271 -6159
rect 4332 -6181 4335 -6159
rect 4387 -6181 4403 -6129
rect 4455 -6181 4467 -6129
rect 4519 -6181 4531 -6129
rect 4583 -6159 4633 -6129
rect 3744 -6193 3782 -6181
rect 3816 -6193 3968 -6181
rect 4002 -6193 4040 -6181
rect 4074 -6193 4226 -6181
rect 4260 -6193 4298 -6181
rect 4332 -6193 4484 -6181
rect 4518 -6193 4556 -6181
rect 4590 -6193 4633 -6159
rect 3529 -6199 4633 -6193
rect 4836 -6118 5214 -6084
rect 5248 -6118 5626 -6084
rect 6873 -6111 6934 -5879
rect 4836 -6156 5626 -6118
rect 4836 -6159 5214 -6156
rect 4836 -6193 4935 -6159
rect 4969 -6193 5007 -6159
rect 5041 -6190 5214 -6159
rect 5248 -6159 5626 -6156
rect 5248 -6190 5421 -6159
rect 5041 -6193 5421 -6190
rect 5455 -6193 5493 -6159
rect 5527 -6193 5626 -6159
rect 833 -6262 856 -6228
rect 890 -6262 1269 -6228
rect 4836 -6228 5626 -6193
rect 5830 -6129 6934 -6111
rect 5830 -6159 5880 -6129
rect 5830 -6193 5873 -6159
rect 5932 -6181 5944 -6129
rect 5996 -6181 6008 -6129
rect 6060 -6181 6076 -6129
rect 6128 -6159 6140 -6129
rect 6192 -6159 6204 -6129
rect 6128 -6181 6131 -6159
rect 6192 -6181 6203 -6159
rect 6256 -6181 6366 -6129
rect 6418 -6159 6430 -6129
rect 6482 -6159 6494 -6129
rect 6423 -6181 6430 -6159
rect 6546 -6181 6562 -6129
rect 6614 -6181 6626 -6129
rect 6678 -6159 6690 -6129
rect 6742 -6159 6934 -6129
rect 6681 -6181 6690 -6159
rect 5907 -6193 5945 -6181
rect 5979 -6193 6131 -6181
rect 6165 -6193 6203 -6181
rect 6237 -6193 6389 -6181
rect 6423 -6193 6461 -6181
rect 6495 -6193 6647 -6181
rect 6681 -6193 6719 -6181
rect 6753 -6193 6934 -6159
rect 5830 -6199 6934 -6193
rect 7056 -5990 7764 -5973
rect 7056 -6042 7094 -5990
rect 7146 -6042 7158 -5990
rect 7210 -6042 7222 -5990
rect 7274 -6042 7290 -5990
rect 7342 -6042 7354 -5990
rect 7406 -6042 7418 -5990
rect 7470 -6042 7482 -5990
rect 7534 -6042 7550 -5990
rect 7602 -6042 7614 -5990
rect 7666 -6042 7678 -5990
rect 7730 -6042 7764 -5990
rect 7056 -6159 7764 -6042
rect 7056 -6193 7099 -6159
rect 7133 -6193 7171 -6159
rect 7205 -6193 7357 -6159
rect 7391 -6193 7429 -6159
rect 7463 -6193 7615 -6159
rect 7649 -6193 7687 -6159
rect 7721 -6193 7764 -6159
rect 7056 -6199 7764 -6193
rect 7886 -6111 7947 -5879
rect 8024 -5797 8990 -5791
rect 8024 -5831 8067 -5797
rect 8101 -5812 8139 -5797
rect 8173 -5812 8325 -5797
rect 8359 -5812 8397 -5797
rect 8431 -5812 8583 -5797
rect 8617 -5812 8655 -5797
rect 8689 -5812 8841 -5797
rect 8875 -5812 8913 -5797
rect 8130 -5831 8139 -5812
rect 8024 -5864 8078 -5831
rect 8130 -5864 8142 -5831
rect 8194 -5864 8206 -5812
rect 8258 -5864 8274 -5812
rect 8390 -5831 8397 -5812
rect 8326 -5864 8338 -5831
rect 8390 -5864 8402 -5831
rect 8454 -5864 8564 -5812
rect 8617 -5831 8628 -5812
rect 8689 -5831 8692 -5812
rect 8616 -5864 8628 -5831
rect 8680 -5864 8692 -5831
rect 8744 -5864 8760 -5812
rect 8812 -5864 8824 -5812
rect 8876 -5864 8888 -5812
rect 8947 -5831 8990 -5797
rect 8940 -5864 8990 -5831
rect 8024 -5990 8990 -5864
rect 8024 -6042 8078 -5990
rect 8130 -6042 8142 -5990
rect 8194 -6042 8206 -5990
rect 8258 -6042 8274 -5990
rect 8326 -6042 8338 -5990
rect 8390 -6042 8402 -5990
rect 8454 -6042 8564 -5990
rect 8616 -6042 8628 -5990
rect 8680 -6042 8692 -5990
rect 8744 -6042 8760 -5990
rect 8812 -6042 8824 -5990
rect 8876 -6042 8888 -5990
rect 8940 -6042 8990 -5990
rect 8024 -6061 8990 -6042
rect 9194 -5796 9986 -5758
rect 13554 -5758 13932 -5724
rect 13966 -5758 14344 -5724
rect 14491 -5597 14537 -5116
rect 14674 -5386 14870 -5378
rect 14674 -5438 14681 -5386
rect 14733 -5438 14745 -5386
rect 14797 -5438 14809 -5386
rect 14861 -5438 14870 -5386
rect 14674 -5448 14870 -5438
rect 14491 -5631 14497 -5597
rect 14531 -5631 14537 -5597
rect 14491 -5669 14537 -5631
rect 14491 -5703 14497 -5669
rect 14531 -5703 14537 -5669
rect 14491 -5750 14537 -5703
rect 14749 -5597 14795 -5448
rect 14749 -5631 14755 -5597
rect 14789 -5631 14795 -5597
rect 14749 -5669 14795 -5631
rect 14749 -5703 14755 -5669
rect 14789 -5703 14795 -5669
rect 14749 -5750 14795 -5703
rect 15007 -5597 15053 -5116
rect 15191 -5386 15387 -5378
rect 15191 -5438 15198 -5386
rect 15250 -5438 15262 -5386
rect 15314 -5438 15326 -5386
rect 15378 -5438 15387 -5386
rect 15191 -5448 15387 -5438
rect 15007 -5631 15013 -5597
rect 15047 -5631 15053 -5597
rect 15007 -5669 15053 -5631
rect 15007 -5703 15013 -5669
rect 15047 -5703 15053 -5669
rect 15007 -5750 15053 -5703
rect 15265 -5597 15311 -5448
rect 15265 -5631 15271 -5597
rect 15305 -5631 15311 -5597
rect 15265 -5669 15311 -5631
rect 15265 -5703 15271 -5669
rect 15305 -5703 15311 -5669
rect 15265 -5750 15311 -5703
rect 15523 -5597 15569 -5116
rect 15523 -5631 15529 -5597
rect 15563 -5631 15569 -5597
rect 15523 -5669 15569 -5631
rect 15523 -5703 15529 -5669
rect 15563 -5703 15569 -5669
rect 15523 -5750 15569 -5703
rect 15717 -5597 15763 -4947
rect 15897 -5217 16093 -5209
rect 15897 -5269 15906 -5217
rect 15958 -5269 15970 -5217
rect 16022 -5269 16034 -5217
rect 16086 -5269 16093 -5217
rect 15897 -5279 16093 -5269
rect 15717 -5631 15723 -5597
rect 15757 -5631 15763 -5597
rect 15717 -5669 15763 -5631
rect 15717 -5703 15723 -5669
rect 15757 -5703 15763 -5669
rect 15717 -5750 15763 -5703
rect 15975 -5597 16021 -5279
rect 15975 -5631 15981 -5597
rect 16015 -5631 16021 -5597
rect 15975 -5669 16021 -5631
rect 15975 -5703 15981 -5669
rect 16015 -5703 16021 -5669
rect 15975 -5750 16021 -5703
rect 16233 -5597 16279 -4947
rect 17911 -4966 18290 -4932
rect 18324 -4966 18347 -4932
rect 17911 -5004 18347 -4966
rect 17911 -5038 18290 -5004
rect 18324 -5038 18347 -5004
rect 16611 -5054 16807 -5046
rect 16611 -5106 16618 -5054
rect 16670 -5106 16682 -5054
rect 16734 -5106 16746 -5054
rect 16798 -5106 16807 -5054
rect 16611 -5116 16807 -5106
rect 17128 -5054 17324 -5046
rect 17128 -5106 17135 -5054
rect 17187 -5106 17199 -5054
rect 17251 -5106 17263 -5054
rect 17315 -5106 17324 -5054
rect 17128 -5116 17324 -5106
rect 17645 -5054 17841 -5046
rect 17645 -5106 17652 -5054
rect 17704 -5106 17716 -5054
rect 17768 -5106 17780 -5054
rect 17832 -5106 17841 -5054
rect 17645 -5116 17841 -5106
rect 17911 -5076 18347 -5038
rect 17911 -5110 18290 -5076
rect 18324 -5110 18347 -5076
rect 16414 -5217 16610 -5209
rect 16414 -5269 16423 -5217
rect 16475 -5269 16487 -5217
rect 16539 -5269 16551 -5217
rect 16603 -5269 16610 -5217
rect 16414 -5279 16610 -5269
rect 16233 -5631 16239 -5597
rect 16273 -5631 16279 -5597
rect 16233 -5669 16279 -5631
rect 16233 -5703 16239 -5669
rect 16273 -5703 16279 -5669
rect 16233 -5750 16279 -5703
rect 16491 -5597 16537 -5279
rect 16491 -5631 16497 -5597
rect 16531 -5631 16537 -5597
rect 16491 -5669 16537 -5631
rect 16491 -5703 16497 -5669
rect 16531 -5703 16537 -5669
rect 16491 -5750 16537 -5703
rect 16685 -5597 16731 -5116
rect 16868 -5386 17064 -5378
rect 16868 -5438 16875 -5386
rect 16927 -5438 16939 -5386
rect 16991 -5438 17003 -5386
rect 17055 -5438 17064 -5386
rect 16868 -5448 17064 -5438
rect 16685 -5631 16691 -5597
rect 16725 -5631 16731 -5597
rect 16685 -5669 16731 -5631
rect 16685 -5703 16691 -5669
rect 16725 -5703 16731 -5669
rect 16685 -5750 16731 -5703
rect 16943 -5597 16989 -5448
rect 16943 -5631 16949 -5597
rect 16983 -5631 16989 -5597
rect 16943 -5669 16989 -5631
rect 16943 -5703 16949 -5669
rect 16983 -5703 16989 -5669
rect 16943 -5750 16989 -5703
rect 17201 -5597 17247 -5116
rect 17386 -5386 17582 -5378
rect 17386 -5438 17393 -5386
rect 17445 -5438 17457 -5386
rect 17509 -5438 17521 -5386
rect 17573 -5438 17582 -5386
rect 17386 -5448 17582 -5438
rect 17201 -5631 17207 -5597
rect 17241 -5631 17247 -5597
rect 17201 -5669 17247 -5631
rect 17201 -5703 17207 -5669
rect 17241 -5703 17247 -5669
rect 17201 -5750 17247 -5703
rect 17459 -5597 17505 -5448
rect 17459 -5631 17465 -5597
rect 17499 -5631 17505 -5597
rect 17459 -5669 17505 -5631
rect 17459 -5703 17465 -5669
rect 17499 -5703 17505 -5669
rect 17459 -5750 17505 -5703
rect 17717 -5597 17763 -5116
rect 17717 -5631 17723 -5597
rect 17757 -5631 17763 -5597
rect 17717 -5669 17763 -5631
rect 17717 -5703 17723 -5669
rect 17757 -5703 17763 -5669
rect 17717 -5750 17763 -5703
rect 17911 -5148 18347 -5110
rect 17911 -5182 18290 -5148
rect 18324 -5182 18347 -5148
rect 17911 -5220 18347 -5182
rect 17911 -5254 18290 -5220
rect 18324 -5254 18347 -5220
rect 17911 -5292 18347 -5254
rect 17911 -5326 18290 -5292
rect 18324 -5326 18347 -5292
rect 17911 -5364 18347 -5326
rect 17911 -5398 18290 -5364
rect 18324 -5398 18347 -5364
rect 17911 -5436 18347 -5398
rect 17911 -5470 18290 -5436
rect 18324 -5470 18347 -5436
rect 17911 -5508 18347 -5470
rect 17911 -5542 18290 -5508
rect 18324 -5542 18347 -5508
rect 17911 -5580 18347 -5542
rect 17911 -5597 18290 -5580
rect 17911 -5631 17917 -5597
rect 17951 -5631 18175 -5597
rect 18209 -5614 18290 -5597
rect 18324 -5614 18347 -5580
rect 18209 -5631 18347 -5614
rect 17911 -5652 18347 -5631
rect 17911 -5669 18290 -5652
rect 17911 -5703 17917 -5669
rect 17951 -5703 18175 -5669
rect 18209 -5686 18290 -5669
rect 18324 -5686 18347 -5652
rect 18209 -5703 18347 -5686
rect 17911 -5724 18347 -5703
rect 9194 -5797 9573 -5796
rect 9194 -5831 9293 -5797
rect 9327 -5831 9365 -5797
rect 9399 -5830 9573 -5797
rect 9607 -5797 9986 -5796
rect 9607 -5830 9781 -5797
rect 9399 -5831 9781 -5830
rect 9815 -5831 9853 -5797
rect 9887 -5831 9986 -5797
rect 9194 -5868 9986 -5831
rect 9194 -5902 9573 -5868
rect 9607 -5902 9986 -5868
rect 9194 -5940 9986 -5902
rect 9194 -5974 9573 -5940
rect 9607 -5974 9986 -5940
rect 9194 -6012 9986 -5974
rect 9194 -6046 9573 -6012
rect 9607 -6046 9986 -6012
rect 9194 -6084 9986 -6046
rect 10190 -5797 11156 -5791
rect 10190 -5831 10233 -5797
rect 10267 -5812 10305 -5797
rect 10339 -5812 10491 -5797
rect 10525 -5812 10563 -5797
rect 10597 -5812 10749 -5797
rect 10783 -5812 10821 -5797
rect 10855 -5812 11007 -5797
rect 11041 -5812 11079 -5797
rect 10190 -5864 10240 -5831
rect 10292 -5864 10304 -5812
rect 10356 -5864 10368 -5812
rect 10420 -5864 10436 -5812
rect 10488 -5831 10491 -5812
rect 10552 -5831 10563 -5812
rect 10488 -5864 10500 -5831
rect 10552 -5864 10564 -5831
rect 10616 -5864 10726 -5812
rect 10783 -5831 10790 -5812
rect 10778 -5864 10790 -5831
rect 10842 -5864 10854 -5831
rect 10906 -5864 10922 -5812
rect 10974 -5864 10986 -5812
rect 11041 -5831 11050 -5812
rect 11113 -5831 11156 -5797
rect 11038 -5864 11050 -5831
rect 11102 -5864 11156 -5831
rect 10190 -5990 11156 -5864
rect 10190 -6042 10240 -5990
rect 10292 -6042 10304 -5990
rect 10356 -6042 10368 -5990
rect 10420 -6042 10436 -5990
rect 10488 -6042 10500 -5990
rect 10552 -6042 10564 -5990
rect 10616 -6042 10726 -5990
rect 10778 -6042 10790 -5990
rect 10842 -6042 10854 -5990
rect 10906 -6042 10922 -5990
rect 10974 -6042 10986 -5990
rect 11038 -6042 11050 -5990
rect 11102 -6042 11156 -5990
rect 10190 -6061 11156 -6042
rect 11233 -5797 12307 -5791
rect 11233 -5831 11459 -5797
rect 11493 -5831 11531 -5797
rect 11565 -5831 11717 -5797
rect 11751 -5831 11789 -5797
rect 11823 -5831 11975 -5797
rect 12009 -5831 12047 -5797
rect 12081 -5831 12307 -5797
rect 11233 -5879 12307 -5831
rect 7886 -6129 8990 -6111
rect 7886 -6159 8078 -6129
rect 8130 -6159 8142 -6129
rect 7886 -6193 8067 -6159
rect 8130 -6181 8139 -6159
rect 8194 -6181 8206 -6129
rect 8258 -6181 8274 -6129
rect 8326 -6159 8338 -6129
rect 8390 -6159 8402 -6129
rect 8390 -6181 8397 -6159
rect 8454 -6181 8564 -6129
rect 8616 -6159 8628 -6129
rect 8680 -6159 8692 -6129
rect 8617 -6181 8628 -6159
rect 8689 -6181 8692 -6159
rect 8744 -6181 8760 -6129
rect 8812 -6181 8824 -6129
rect 8876 -6181 8888 -6129
rect 8940 -6159 8990 -6129
rect 8101 -6193 8139 -6181
rect 8173 -6193 8325 -6181
rect 8359 -6193 8397 -6181
rect 8431 -6193 8583 -6181
rect 8617 -6193 8655 -6181
rect 8689 -6193 8841 -6181
rect 8875 -6193 8913 -6181
rect 8947 -6193 8990 -6159
rect 7886 -6199 8990 -6193
rect 9194 -6118 9573 -6084
rect 9607 -6118 9986 -6084
rect 11233 -6111 11294 -5879
rect 9194 -6156 9986 -6118
rect 9194 -6159 9573 -6156
rect 9194 -6193 9293 -6159
rect 9327 -6193 9365 -6159
rect 9399 -6190 9573 -6159
rect 9607 -6159 9986 -6156
rect 9607 -6190 9781 -6159
rect 9399 -6193 9781 -6190
rect 9815 -6193 9853 -6159
rect 9887 -6193 9986 -6159
rect 833 -6287 1269 -6262
rect 833 -6300 971 -6287
rect 833 -6334 856 -6300
rect 890 -6321 971 -6300
rect 1005 -6321 1229 -6287
rect 1263 -6321 1269 -6287
rect 890 -6334 1269 -6321
rect 833 -6359 1269 -6334
rect 833 -6372 971 -6359
rect 833 -6406 856 -6372
rect 890 -6393 971 -6372
rect 1005 -6393 1229 -6359
rect 1263 -6393 1269 -6359
rect 890 -6406 1269 -6393
rect 833 -6444 1269 -6406
rect 833 -6478 856 -6444
rect 890 -6478 1269 -6444
rect 833 -6516 1269 -6478
rect 833 -6550 856 -6516
rect 890 -6550 1269 -6516
rect 833 -6588 1269 -6550
rect 833 -6622 856 -6588
rect 890 -6622 1269 -6588
rect 833 -6660 1269 -6622
rect 833 -6694 856 -6660
rect 890 -6694 1269 -6660
rect 833 -6732 1269 -6694
rect 833 -6766 856 -6732
rect 890 -6766 1269 -6732
rect 833 -6804 1269 -6766
rect 833 -6838 856 -6804
rect 890 -6838 1269 -6804
rect 833 -6876 1269 -6838
rect 833 -6910 856 -6876
rect 890 -6910 1269 -6876
rect 833 -6948 1269 -6910
rect 833 -6982 856 -6948
rect 890 -6982 1269 -6948
rect 833 -7020 1269 -6982
rect 1417 -6287 1463 -6240
rect 1417 -6321 1423 -6287
rect 1457 -6321 1463 -6287
rect 1417 -6359 1463 -6321
rect 1417 -6393 1423 -6359
rect 1457 -6393 1463 -6359
rect 1417 -7000 1463 -6393
rect 1675 -6287 1721 -6240
rect 1675 -6321 1681 -6287
rect 1715 -6321 1721 -6287
rect 1675 -6359 1721 -6321
rect 1675 -6393 1681 -6359
rect 1715 -6393 1721 -6359
rect 1675 -6699 1721 -6393
rect 1933 -6287 1979 -6240
rect 1933 -6321 1939 -6287
rect 1973 -6321 1979 -6287
rect 1933 -6359 1979 -6321
rect 1933 -6393 1939 -6359
rect 1973 -6393 1979 -6359
rect 1601 -6709 1797 -6699
rect 1601 -6761 1608 -6709
rect 1660 -6761 1672 -6709
rect 1724 -6761 1736 -6709
rect 1788 -6761 1797 -6709
rect 1601 -6769 1797 -6761
rect 833 -7054 856 -7020
rect 890 -7054 1269 -7020
rect 833 -7092 1269 -7054
rect 1343 -7010 1539 -7000
rect 1343 -7062 1350 -7010
rect 1402 -7062 1414 -7010
rect 1466 -7062 1478 -7010
rect 1530 -7062 1539 -7010
rect 1343 -7070 1539 -7062
rect 833 -7126 856 -7092
rect 890 -7126 1269 -7092
rect 833 -7164 1269 -7126
rect 833 -7198 856 -7164
rect 890 -7198 1269 -7164
rect 833 -7236 1269 -7198
rect 833 -7270 856 -7236
rect 890 -7244 1269 -7236
rect 890 -7270 971 -7244
rect 833 -7278 971 -7270
rect 1005 -7278 1229 -7244
rect 1263 -7278 1269 -7244
rect 833 -7308 1269 -7278
rect 833 -7342 856 -7308
rect 890 -7316 1269 -7308
rect 890 -7342 971 -7316
rect 833 -7350 971 -7342
rect 1005 -7350 1229 -7316
rect 1263 -7350 1269 -7316
rect 833 -7380 1269 -7350
rect 833 -7414 856 -7380
rect 890 -7414 1269 -7380
rect 1417 -7244 1463 -7070
rect 1417 -7278 1423 -7244
rect 1457 -7278 1463 -7244
rect 1417 -7316 1463 -7278
rect 1417 -7350 1423 -7316
rect 1457 -7350 1463 -7316
rect 1417 -7397 1463 -7350
rect 1675 -7244 1721 -6769
rect 1933 -7000 1979 -6393
rect 2191 -6287 2237 -6240
rect 2191 -6321 2197 -6287
rect 2231 -6321 2237 -6287
rect 2191 -6359 2237 -6321
rect 2191 -6393 2197 -6359
rect 2231 -6393 2237 -6359
rect 2191 -6699 2237 -6393
rect 2449 -6287 2495 -6240
rect 2449 -6321 2455 -6287
rect 2489 -6321 2495 -6287
rect 2449 -6359 2495 -6321
rect 2449 -6393 2455 -6359
rect 2489 -6393 2495 -6359
rect 2119 -6709 2315 -6699
rect 2119 -6761 2126 -6709
rect 2178 -6761 2190 -6709
rect 2242 -6761 2254 -6709
rect 2306 -6761 2315 -6709
rect 2119 -6769 2315 -6761
rect 1858 -7010 2054 -7000
rect 1858 -7062 1865 -7010
rect 1917 -7062 1929 -7010
rect 1981 -7062 1993 -7010
rect 2045 -7062 2054 -7010
rect 1858 -7070 2054 -7062
rect 1675 -7278 1681 -7244
rect 1715 -7278 1721 -7244
rect 1675 -7316 1721 -7278
rect 1675 -7350 1681 -7316
rect 1715 -7350 1721 -7316
rect 1675 -7397 1721 -7350
rect 1933 -7244 1979 -7070
rect 1933 -7278 1939 -7244
rect 1973 -7278 1979 -7244
rect 1933 -7316 1979 -7278
rect 1933 -7350 1939 -7316
rect 1973 -7350 1979 -7316
rect 1933 -7397 1979 -7350
rect 2191 -7244 2237 -6769
rect 2449 -7000 2495 -6393
rect 2643 -6287 2689 -6240
rect 2643 -6321 2649 -6287
rect 2683 -6321 2689 -6287
rect 2643 -6359 2689 -6321
rect 2643 -6393 2649 -6359
rect 2683 -6393 2689 -6359
rect 2643 -6554 2689 -6393
rect 2901 -6287 2947 -6240
rect 2901 -6321 2907 -6287
rect 2941 -6321 2947 -6287
rect 2901 -6359 2947 -6321
rect 2901 -6393 2907 -6359
rect 2941 -6393 2947 -6359
rect 2566 -6564 2762 -6554
rect 2566 -6616 2575 -6564
rect 2627 -6616 2639 -6564
rect 2691 -6616 2703 -6564
rect 2755 -6616 2762 -6564
rect 2566 -6624 2762 -6616
rect 2376 -7010 2572 -7000
rect 2376 -7062 2383 -7010
rect 2435 -7062 2447 -7010
rect 2499 -7062 2511 -7010
rect 2563 -7062 2572 -7010
rect 2376 -7070 2572 -7062
rect 2191 -7278 2197 -7244
rect 2231 -7278 2237 -7244
rect 2191 -7316 2237 -7278
rect 2191 -7350 2197 -7316
rect 2231 -7350 2237 -7316
rect 2191 -7397 2237 -7350
rect 2449 -7244 2495 -7070
rect 2449 -7278 2455 -7244
rect 2489 -7278 2495 -7244
rect 2449 -7316 2495 -7278
rect 2449 -7350 2455 -7316
rect 2489 -7350 2495 -7316
rect 2449 -7397 2495 -7350
rect 2643 -7244 2689 -6624
rect 2901 -6860 2947 -6393
rect 3159 -6287 3205 -6240
rect 3159 -6321 3165 -6287
rect 3199 -6321 3205 -6287
rect 3159 -6359 3205 -6321
rect 3159 -6393 3165 -6359
rect 3199 -6393 3205 -6359
rect 3159 -6554 3205 -6393
rect 3417 -6287 3463 -6240
rect 3417 -6321 3423 -6287
rect 3457 -6321 3463 -6287
rect 3417 -6359 3463 -6321
rect 3417 -6393 3423 -6359
rect 3457 -6393 3463 -6359
rect 3083 -6564 3279 -6554
rect 3083 -6616 3092 -6564
rect 3144 -6616 3156 -6564
rect 3208 -6616 3220 -6564
rect 3272 -6616 3279 -6564
rect 3083 -6624 3279 -6616
rect 2824 -6870 3020 -6860
rect 2824 -6922 2833 -6870
rect 2885 -6922 2897 -6870
rect 2949 -6922 2961 -6870
rect 3013 -6922 3020 -6870
rect 2824 -6930 3020 -6922
rect 2643 -7278 2649 -7244
rect 2683 -7278 2689 -7244
rect 2643 -7316 2689 -7278
rect 2643 -7350 2649 -7316
rect 2683 -7350 2689 -7316
rect 2643 -7397 2689 -7350
rect 2901 -7244 2947 -6930
rect 2901 -7278 2907 -7244
rect 2941 -7278 2947 -7244
rect 2901 -7316 2947 -7278
rect 2901 -7350 2907 -7316
rect 2941 -7350 2947 -7316
rect 2901 -7397 2947 -7350
rect 3159 -7244 3205 -6624
rect 3417 -6860 3463 -6393
rect 3611 -6287 3657 -6240
rect 3611 -6321 3617 -6287
rect 3651 -6321 3657 -6287
rect 3611 -6359 3657 -6321
rect 3611 -6393 3617 -6359
rect 3651 -6393 3657 -6359
rect 3341 -6870 3537 -6860
rect 3341 -6922 3350 -6870
rect 3402 -6922 3414 -6870
rect 3466 -6922 3478 -6870
rect 3530 -6922 3537 -6870
rect 3341 -6930 3537 -6922
rect 3159 -7278 3165 -7244
rect 3199 -7278 3205 -7244
rect 3159 -7316 3205 -7278
rect 3159 -7350 3165 -7316
rect 3199 -7350 3205 -7316
rect 3159 -7397 3205 -7350
rect 3417 -7244 3463 -6930
rect 3611 -7000 3657 -6393
rect 3869 -6287 3915 -6240
rect 3869 -6321 3875 -6287
rect 3909 -6321 3915 -6287
rect 3869 -6359 3915 -6321
rect 3869 -6393 3875 -6359
rect 3909 -6393 3915 -6359
rect 3869 -6699 3915 -6393
rect 4127 -6287 4173 -6240
rect 4127 -6321 4133 -6287
rect 4167 -6321 4173 -6287
rect 4127 -6359 4173 -6321
rect 4127 -6393 4133 -6359
rect 4167 -6393 4173 -6359
rect 3796 -6709 3992 -6699
rect 3796 -6761 3803 -6709
rect 3855 -6761 3867 -6709
rect 3919 -6761 3931 -6709
rect 3983 -6761 3992 -6709
rect 3796 -6769 3992 -6761
rect 3536 -7010 3732 -7000
rect 3536 -7062 3543 -7010
rect 3595 -7062 3607 -7010
rect 3659 -7062 3671 -7010
rect 3723 -7062 3732 -7010
rect 3536 -7070 3732 -7062
rect 3417 -7278 3423 -7244
rect 3457 -7278 3463 -7244
rect 3417 -7316 3463 -7278
rect 3417 -7350 3423 -7316
rect 3457 -7350 3463 -7316
rect 3417 -7397 3463 -7350
rect 3611 -7244 3657 -7070
rect 3611 -7278 3617 -7244
rect 3651 -7278 3657 -7244
rect 3611 -7316 3657 -7278
rect 3611 -7350 3617 -7316
rect 3651 -7350 3657 -7316
rect 3611 -7397 3657 -7350
rect 3869 -7244 3915 -6769
rect 4127 -7000 4173 -6393
rect 4385 -6287 4431 -6240
rect 4385 -6321 4391 -6287
rect 4425 -6321 4431 -6287
rect 4385 -6359 4431 -6321
rect 4385 -6393 4391 -6359
rect 4425 -6393 4431 -6359
rect 4385 -6699 4431 -6393
rect 4643 -6287 4689 -6240
rect 4643 -6321 4649 -6287
rect 4683 -6321 4689 -6287
rect 4643 -6359 4689 -6321
rect 4643 -6393 4649 -6359
rect 4683 -6393 4689 -6359
rect 4313 -6709 4509 -6699
rect 4313 -6761 4320 -6709
rect 4372 -6761 4384 -6709
rect 4436 -6761 4448 -6709
rect 4500 -6761 4509 -6709
rect 4313 -6769 4509 -6761
rect 4053 -7010 4249 -7000
rect 4053 -7062 4060 -7010
rect 4112 -7062 4124 -7010
rect 4176 -7062 4188 -7010
rect 4240 -7062 4249 -7010
rect 4053 -7070 4249 -7062
rect 3869 -7278 3875 -7244
rect 3909 -7278 3915 -7244
rect 3869 -7316 3915 -7278
rect 3869 -7350 3875 -7316
rect 3909 -7350 3915 -7316
rect 3869 -7397 3915 -7350
rect 4127 -7244 4173 -7070
rect 4127 -7278 4133 -7244
rect 4167 -7278 4173 -7244
rect 4127 -7316 4173 -7278
rect 4127 -7350 4133 -7316
rect 4167 -7350 4173 -7316
rect 4127 -7397 4173 -7350
rect 4385 -7244 4431 -6769
rect 4643 -7000 4689 -6393
rect 4836 -6262 5214 -6228
rect 5248 -6262 5626 -6228
rect 9194 -6228 9986 -6193
rect 10190 -6129 11294 -6111
rect 10190 -6159 10240 -6129
rect 10190 -6193 10233 -6159
rect 10292 -6181 10304 -6129
rect 10356 -6181 10368 -6129
rect 10420 -6181 10436 -6129
rect 10488 -6159 10500 -6129
rect 10552 -6159 10564 -6129
rect 10488 -6181 10491 -6159
rect 10552 -6181 10563 -6159
rect 10616 -6181 10726 -6129
rect 10778 -6159 10790 -6129
rect 10842 -6159 10854 -6129
rect 10783 -6181 10790 -6159
rect 10906 -6181 10922 -6129
rect 10974 -6181 10986 -6129
rect 11038 -6159 11050 -6129
rect 11102 -6159 11294 -6129
rect 11041 -6181 11050 -6159
rect 10267 -6193 10305 -6181
rect 10339 -6193 10491 -6181
rect 10525 -6193 10563 -6181
rect 10597 -6193 10749 -6181
rect 10783 -6193 10821 -6181
rect 10855 -6193 11007 -6181
rect 11041 -6193 11079 -6181
rect 11113 -6193 11294 -6159
rect 10190 -6199 11294 -6193
rect 11416 -5990 12124 -5973
rect 11416 -6042 11450 -5990
rect 11502 -6042 11514 -5990
rect 11566 -6042 11578 -5990
rect 11630 -6042 11646 -5990
rect 11698 -6042 11710 -5990
rect 11762 -6042 11774 -5990
rect 11826 -6042 11838 -5990
rect 11890 -6042 11906 -5990
rect 11958 -6042 11970 -5990
rect 12022 -6042 12034 -5990
rect 12086 -6042 12124 -5990
rect 11416 -6159 12124 -6042
rect 11416 -6193 11459 -6159
rect 11493 -6193 11531 -6159
rect 11565 -6193 11717 -6159
rect 11751 -6193 11789 -6159
rect 11823 -6193 11975 -6159
rect 12009 -6193 12047 -6159
rect 12081 -6193 12124 -6159
rect 11416 -6199 12124 -6193
rect 12246 -6111 12307 -5879
rect 12384 -5797 13350 -5791
rect 12384 -5831 12427 -5797
rect 12461 -5812 12499 -5797
rect 12533 -5812 12685 -5797
rect 12719 -5812 12757 -5797
rect 12791 -5812 12943 -5797
rect 12977 -5812 13015 -5797
rect 13049 -5812 13201 -5797
rect 13235 -5812 13273 -5797
rect 12490 -5831 12499 -5812
rect 12384 -5864 12438 -5831
rect 12490 -5864 12502 -5831
rect 12554 -5864 12566 -5812
rect 12618 -5864 12634 -5812
rect 12750 -5831 12757 -5812
rect 12686 -5864 12698 -5831
rect 12750 -5864 12762 -5831
rect 12814 -5864 12924 -5812
rect 12977 -5831 12988 -5812
rect 13049 -5831 13052 -5812
rect 12976 -5864 12988 -5831
rect 13040 -5864 13052 -5831
rect 13104 -5864 13120 -5812
rect 13172 -5864 13184 -5812
rect 13236 -5864 13248 -5812
rect 13307 -5831 13350 -5797
rect 13300 -5864 13350 -5831
rect 12384 -5990 13350 -5864
rect 12384 -6042 12438 -5990
rect 12490 -6042 12502 -5990
rect 12554 -6042 12566 -5990
rect 12618 -6042 12634 -5990
rect 12686 -6042 12698 -5990
rect 12750 -6042 12762 -5990
rect 12814 -6042 12924 -5990
rect 12976 -6042 12988 -5990
rect 13040 -6042 13052 -5990
rect 13104 -6042 13120 -5990
rect 13172 -6042 13184 -5990
rect 13236 -6042 13248 -5990
rect 13300 -6042 13350 -5990
rect 12384 -6061 13350 -6042
rect 13554 -5796 14344 -5758
rect 17911 -5758 18290 -5724
rect 18324 -5758 18347 -5724
rect 13554 -5797 13932 -5796
rect 13554 -5831 13653 -5797
rect 13687 -5831 13725 -5797
rect 13759 -5830 13932 -5797
rect 13966 -5797 14344 -5796
rect 13966 -5830 14139 -5797
rect 13759 -5831 14139 -5830
rect 14173 -5831 14211 -5797
rect 14245 -5831 14344 -5797
rect 13554 -5868 14344 -5831
rect 13554 -5902 13932 -5868
rect 13966 -5902 14344 -5868
rect 13554 -5940 14344 -5902
rect 13554 -5974 13932 -5940
rect 13966 -5974 14344 -5940
rect 13554 -6012 14344 -5974
rect 13554 -6046 13932 -6012
rect 13966 -6046 14344 -6012
rect 13554 -6084 14344 -6046
rect 14547 -5797 15513 -5791
rect 14547 -5831 14590 -5797
rect 14624 -5812 14662 -5797
rect 14696 -5812 14848 -5797
rect 14882 -5812 14920 -5797
rect 14954 -5812 15106 -5797
rect 15140 -5812 15178 -5797
rect 15212 -5812 15364 -5797
rect 15398 -5812 15436 -5797
rect 14547 -5864 14597 -5831
rect 14649 -5864 14661 -5812
rect 14713 -5864 14725 -5812
rect 14777 -5864 14793 -5812
rect 14845 -5831 14848 -5812
rect 14909 -5831 14920 -5812
rect 14845 -5864 14857 -5831
rect 14909 -5864 14921 -5831
rect 14973 -5864 15083 -5812
rect 15140 -5831 15147 -5812
rect 15135 -5864 15147 -5831
rect 15199 -5864 15211 -5831
rect 15263 -5864 15279 -5812
rect 15331 -5864 15343 -5812
rect 15398 -5831 15407 -5812
rect 15470 -5831 15513 -5797
rect 15395 -5864 15407 -5831
rect 15459 -5864 15513 -5831
rect 14547 -5990 15513 -5864
rect 14547 -6042 14597 -5990
rect 14649 -6042 14661 -5990
rect 14713 -6042 14725 -5990
rect 14777 -6042 14793 -5990
rect 14845 -6042 14857 -5990
rect 14909 -6042 14921 -5990
rect 14973 -6042 15083 -5990
rect 15135 -6042 15147 -5990
rect 15199 -6042 15211 -5990
rect 15263 -6042 15279 -5990
rect 15331 -6042 15343 -5990
rect 15395 -6042 15407 -5990
rect 15459 -6042 15513 -5990
rect 14547 -6061 15513 -6042
rect 15590 -5797 16664 -5791
rect 15590 -5831 15816 -5797
rect 15850 -5831 15888 -5797
rect 15922 -5831 16074 -5797
rect 16108 -5831 16146 -5797
rect 16180 -5831 16332 -5797
rect 16366 -5831 16404 -5797
rect 16438 -5831 16664 -5797
rect 15590 -5879 16664 -5831
rect 12246 -6129 13350 -6111
rect 12246 -6159 12438 -6129
rect 12490 -6159 12502 -6129
rect 12246 -6193 12427 -6159
rect 12490 -6181 12499 -6159
rect 12554 -6181 12566 -6129
rect 12618 -6181 12634 -6129
rect 12686 -6159 12698 -6129
rect 12750 -6159 12762 -6129
rect 12750 -6181 12757 -6159
rect 12814 -6181 12924 -6129
rect 12976 -6159 12988 -6129
rect 13040 -6159 13052 -6129
rect 12977 -6181 12988 -6159
rect 13049 -6181 13052 -6159
rect 13104 -6181 13120 -6129
rect 13172 -6181 13184 -6129
rect 13236 -6181 13248 -6129
rect 13300 -6159 13350 -6129
rect 12461 -6193 12499 -6181
rect 12533 -6193 12685 -6181
rect 12719 -6193 12757 -6181
rect 12791 -6193 12943 -6181
rect 12977 -6193 13015 -6181
rect 13049 -6193 13201 -6181
rect 13235 -6193 13273 -6181
rect 13307 -6193 13350 -6159
rect 12246 -6199 13350 -6193
rect 13554 -6118 13932 -6084
rect 13966 -6118 14344 -6084
rect 15590 -6111 15651 -5879
rect 13554 -6156 14344 -6118
rect 13554 -6159 13932 -6156
rect 13554 -6193 13653 -6159
rect 13687 -6193 13725 -6159
rect 13759 -6190 13932 -6159
rect 13966 -6159 14344 -6156
rect 13966 -6190 14139 -6159
rect 13759 -6193 14139 -6190
rect 14173 -6193 14211 -6159
rect 14245 -6193 14344 -6159
rect 4836 -6287 5626 -6262
rect 4836 -6321 4842 -6287
rect 4876 -6321 5100 -6287
rect 5134 -6300 5328 -6287
rect 5134 -6321 5214 -6300
rect 4836 -6334 5214 -6321
rect 5248 -6321 5328 -6300
rect 5362 -6321 5586 -6287
rect 5620 -6321 5626 -6287
rect 5248 -6334 5626 -6321
rect 4836 -6359 5626 -6334
rect 4836 -6393 4842 -6359
rect 4876 -6393 5100 -6359
rect 5134 -6372 5328 -6359
rect 5134 -6393 5214 -6372
rect 4836 -6406 5214 -6393
rect 5248 -6393 5328 -6372
rect 5362 -6393 5586 -6359
rect 5620 -6393 5626 -6359
rect 5248 -6406 5626 -6393
rect 4836 -6444 5626 -6406
rect 4836 -6478 5214 -6444
rect 5248 -6478 5626 -6444
rect 4836 -6516 5626 -6478
rect 4836 -6550 5214 -6516
rect 5248 -6550 5626 -6516
rect 4836 -6588 5626 -6550
rect 4836 -6622 5214 -6588
rect 5248 -6622 5626 -6588
rect 4836 -6660 5626 -6622
rect 4836 -6694 5214 -6660
rect 5248 -6694 5626 -6660
rect 4836 -6732 5626 -6694
rect 4836 -6766 5214 -6732
rect 5248 -6766 5626 -6732
rect 4836 -6804 5626 -6766
rect 4836 -6838 5214 -6804
rect 5248 -6838 5626 -6804
rect 4836 -6876 5626 -6838
rect 4836 -6910 5214 -6876
rect 5248 -6910 5626 -6876
rect 4836 -6948 5626 -6910
rect 4836 -6982 5214 -6948
rect 5248 -6982 5626 -6948
rect 4570 -7010 4766 -7000
rect 4570 -7062 4577 -7010
rect 4629 -7062 4641 -7010
rect 4693 -7062 4705 -7010
rect 4757 -7062 4766 -7010
rect 4570 -7070 4766 -7062
rect 4836 -7020 5626 -6982
rect 5774 -6287 5820 -6240
rect 5774 -6321 5780 -6287
rect 5814 -6321 5820 -6287
rect 5774 -6359 5820 -6321
rect 5774 -6393 5780 -6359
rect 5814 -6393 5820 -6359
rect 5774 -7000 5820 -6393
rect 6032 -6287 6078 -6240
rect 6032 -6321 6038 -6287
rect 6072 -6321 6078 -6287
rect 6032 -6359 6078 -6321
rect 6032 -6393 6038 -6359
rect 6072 -6393 6078 -6359
rect 6032 -6699 6078 -6393
rect 6290 -6287 6336 -6240
rect 6290 -6321 6296 -6287
rect 6330 -6321 6336 -6287
rect 6290 -6359 6336 -6321
rect 6290 -6393 6296 -6359
rect 6330 -6393 6336 -6359
rect 5954 -6709 6150 -6699
rect 5954 -6761 5963 -6709
rect 6015 -6761 6027 -6709
rect 6079 -6761 6091 -6709
rect 6143 -6761 6150 -6709
rect 5954 -6769 6150 -6761
rect 4836 -7054 5214 -7020
rect 5248 -7054 5626 -7020
rect 4385 -7278 4391 -7244
rect 4425 -7278 4431 -7244
rect 4385 -7316 4431 -7278
rect 4385 -7350 4391 -7316
rect 4425 -7350 4431 -7316
rect 4385 -7397 4431 -7350
rect 4643 -7244 4689 -7070
rect 4643 -7278 4649 -7244
rect 4683 -7278 4689 -7244
rect 4643 -7316 4689 -7278
rect 4643 -7350 4649 -7316
rect 4683 -7350 4689 -7316
rect 4643 -7397 4689 -7350
rect 4836 -7092 5626 -7054
rect 5697 -7010 5893 -7000
rect 5697 -7062 5706 -7010
rect 5758 -7062 5770 -7010
rect 5822 -7062 5834 -7010
rect 5886 -7062 5893 -7010
rect 5697 -7070 5893 -7062
rect 4836 -7126 5214 -7092
rect 5248 -7126 5626 -7092
rect 4836 -7164 5626 -7126
rect 4836 -7198 5214 -7164
rect 5248 -7198 5626 -7164
rect 4836 -7236 5626 -7198
rect 4836 -7244 5214 -7236
rect 4836 -7278 4842 -7244
rect 4876 -7278 5100 -7244
rect 5134 -7270 5214 -7244
rect 5248 -7244 5626 -7236
rect 5248 -7270 5328 -7244
rect 5134 -7278 5328 -7270
rect 5362 -7278 5586 -7244
rect 5620 -7278 5626 -7244
rect 4836 -7308 5626 -7278
rect 4836 -7316 5214 -7308
rect 4836 -7350 4842 -7316
rect 4876 -7350 5100 -7316
rect 5134 -7342 5214 -7316
rect 5248 -7316 5626 -7308
rect 5248 -7342 5328 -7316
rect 5134 -7350 5328 -7342
rect 5362 -7350 5586 -7316
rect 5620 -7350 5626 -7316
rect 4836 -7380 5626 -7350
rect 833 -7444 1269 -7414
rect 4836 -7414 5214 -7380
rect 5248 -7414 5626 -7380
rect 5774 -7244 5820 -7070
rect 5774 -7278 5780 -7244
rect 5814 -7278 5820 -7244
rect 5774 -7316 5820 -7278
rect 5774 -7350 5780 -7316
rect 5814 -7350 5820 -7316
rect 5774 -7397 5820 -7350
rect 6032 -7244 6078 -6769
rect 6290 -7000 6336 -6393
rect 6548 -6287 6594 -6240
rect 6548 -6321 6554 -6287
rect 6588 -6321 6594 -6287
rect 6548 -6359 6594 -6321
rect 6548 -6393 6554 -6359
rect 6588 -6393 6594 -6359
rect 6548 -6699 6594 -6393
rect 6806 -6287 6852 -6240
rect 6806 -6321 6812 -6287
rect 6846 -6321 6852 -6287
rect 6806 -6359 6852 -6321
rect 6806 -6393 6812 -6359
rect 6846 -6393 6852 -6359
rect 6471 -6709 6667 -6699
rect 6471 -6761 6480 -6709
rect 6532 -6761 6544 -6709
rect 6596 -6761 6608 -6709
rect 6660 -6761 6667 -6709
rect 6471 -6769 6667 -6761
rect 6214 -7010 6410 -7000
rect 6214 -7062 6223 -7010
rect 6275 -7062 6287 -7010
rect 6339 -7062 6351 -7010
rect 6403 -7062 6410 -7010
rect 6214 -7070 6410 -7062
rect 6032 -7278 6038 -7244
rect 6072 -7278 6078 -7244
rect 6032 -7316 6078 -7278
rect 6032 -7350 6038 -7316
rect 6072 -7350 6078 -7316
rect 6032 -7397 6078 -7350
rect 6290 -7244 6336 -7070
rect 6290 -7278 6296 -7244
rect 6330 -7278 6336 -7244
rect 6290 -7316 6336 -7278
rect 6290 -7350 6296 -7316
rect 6330 -7350 6336 -7316
rect 6290 -7397 6336 -7350
rect 6548 -7244 6594 -6769
rect 6806 -7000 6852 -6393
rect 7000 -6287 7046 -6240
rect 7000 -6321 7006 -6287
rect 7040 -6321 7046 -6287
rect 7000 -6359 7046 -6321
rect 7000 -6393 7006 -6359
rect 7040 -6393 7046 -6359
rect 7000 -6860 7046 -6393
rect 7258 -6287 7304 -6240
rect 7258 -6321 7264 -6287
rect 7298 -6321 7304 -6287
rect 7258 -6359 7304 -6321
rect 7258 -6393 7264 -6359
rect 7298 -6393 7304 -6359
rect 7258 -6554 7304 -6393
rect 7516 -6287 7562 -6240
rect 7516 -6321 7522 -6287
rect 7556 -6321 7562 -6287
rect 7516 -6359 7562 -6321
rect 7516 -6393 7522 -6359
rect 7556 -6393 7562 -6359
rect 7184 -6564 7380 -6554
rect 7184 -6616 7191 -6564
rect 7243 -6616 7255 -6564
rect 7307 -6616 7319 -6564
rect 7371 -6616 7380 -6564
rect 7184 -6624 7380 -6616
rect 6926 -6870 7122 -6860
rect 6926 -6922 6933 -6870
rect 6985 -6922 6997 -6870
rect 7049 -6922 7061 -6870
rect 7113 -6922 7122 -6870
rect 6926 -6930 7122 -6922
rect 6731 -7010 6927 -7000
rect 6731 -7062 6740 -7010
rect 6792 -7062 6804 -7010
rect 6856 -7062 6868 -7010
rect 6920 -7062 6927 -7010
rect 6731 -7070 6927 -7062
rect 6548 -7278 6554 -7244
rect 6588 -7278 6594 -7244
rect 6548 -7316 6594 -7278
rect 6548 -7350 6554 -7316
rect 6588 -7350 6594 -7316
rect 6548 -7397 6594 -7350
rect 6806 -7244 6852 -7070
rect 6806 -7278 6812 -7244
rect 6846 -7278 6852 -7244
rect 6806 -7316 6852 -7278
rect 6806 -7350 6812 -7316
rect 6846 -7350 6852 -7316
rect 6806 -7397 6852 -7350
rect 7000 -7244 7046 -6930
rect 7000 -7278 7006 -7244
rect 7040 -7278 7046 -7244
rect 7000 -7316 7046 -7278
rect 7000 -7350 7006 -7316
rect 7040 -7350 7046 -7316
rect 7000 -7397 7046 -7350
rect 7258 -7244 7304 -6624
rect 7516 -6860 7562 -6393
rect 7774 -6287 7820 -6240
rect 7774 -6321 7780 -6287
rect 7814 -6321 7820 -6287
rect 7774 -6359 7820 -6321
rect 7774 -6393 7780 -6359
rect 7814 -6393 7820 -6359
rect 7774 -6554 7820 -6393
rect 7968 -6287 8014 -6240
rect 7968 -6321 7974 -6287
rect 8008 -6321 8014 -6287
rect 7968 -6359 8014 -6321
rect 7968 -6393 7974 -6359
rect 8008 -6393 8014 -6359
rect 7701 -6564 7897 -6554
rect 7701 -6616 7708 -6564
rect 7760 -6616 7772 -6564
rect 7824 -6616 7836 -6564
rect 7888 -6616 7897 -6564
rect 7701 -6624 7897 -6616
rect 7443 -6870 7639 -6860
rect 7443 -6922 7450 -6870
rect 7502 -6922 7514 -6870
rect 7566 -6922 7578 -6870
rect 7630 -6922 7639 -6870
rect 7443 -6930 7639 -6922
rect 7258 -7278 7264 -7244
rect 7298 -7278 7304 -7244
rect 7258 -7316 7304 -7278
rect 7258 -7350 7264 -7316
rect 7298 -7350 7304 -7316
rect 7258 -7397 7304 -7350
rect 7516 -7244 7562 -6930
rect 7516 -7278 7522 -7244
rect 7556 -7278 7562 -7244
rect 7516 -7316 7562 -7278
rect 7516 -7350 7522 -7316
rect 7556 -7350 7562 -7316
rect 7516 -7397 7562 -7350
rect 7774 -7244 7820 -6624
rect 7968 -7000 8014 -6393
rect 8226 -6287 8272 -6240
rect 8226 -6321 8232 -6287
rect 8266 -6321 8272 -6287
rect 8226 -6359 8272 -6321
rect 8226 -6393 8232 -6359
rect 8266 -6393 8272 -6359
rect 8226 -6699 8272 -6393
rect 8484 -6287 8530 -6240
rect 8484 -6321 8490 -6287
rect 8524 -6321 8530 -6287
rect 8484 -6359 8530 -6321
rect 8484 -6393 8490 -6359
rect 8524 -6393 8530 -6359
rect 8148 -6709 8344 -6699
rect 8148 -6761 8157 -6709
rect 8209 -6761 8221 -6709
rect 8273 -6761 8285 -6709
rect 8337 -6761 8344 -6709
rect 8148 -6769 8344 -6761
rect 7891 -7010 8087 -7000
rect 7891 -7062 7900 -7010
rect 7952 -7062 7964 -7010
rect 8016 -7062 8028 -7010
rect 8080 -7062 8087 -7010
rect 7891 -7070 8087 -7062
rect 7774 -7278 7780 -7244
rect 7814 -7278 7820 -7244
rect 7774 -7316 7820 -7278
rect 7774 -7350 7780 -7316
rect 7814 -7350 7820 -7316
rect 7774 -7397 7820 -7350
rect 7968 -7244 8014 -7070
rect 7968 -7278 7974 -7244
rect 8008 -7278 8014 -7244
rect 7968 -7316 8014 -7278
rect 7968 -7350 7974 -7316
rect 8008 -7350 8014 -7316
rect 7968 -7397 8014 -7350
rect 8226 -7244 8272 -6769
rect 8484 -7000 8530 -6393
rect 8742 -6287 8788 -6240
rect 8742 -6321 8748 -6287
rect 8782 -6321 8788 -6287
rect 8742 -6359 8788 -6321
rect 8742 -6393 8748 -6359
rect 8782 -6393 8788 -6359
rect 8742 -6699 8788 -6393
rect 9000 -6287 9046 -6240
rect 9000 -6321 9006 -6287
rect 9040 -6321 9046 -6287
rect 9000 -6359 9046 -6321
rect 9000 -6393 9006 -6359
rect 9040 -6393 9046 -6359
rect 8665 -6709 8861 -6699
rect 8665 -6761 8674 -6709
rect 8726 -6761 8738 -6709
rect 8790 -6761 8802 -6709
rect 8854 -6761 8861 -6709
rect 8665 -6769 8861 -6761
rect 8408 -7010 8604 -7000
rect 8408 -7062 8417 -7010
rect 8469 -7062 8481 -7010
rect 8533 -7062 8545 -7010
rect 8597 -7062 8604 -7010
rect 8408 -7070 8604 -7062
rect 8226 -7278 8232 -7244
rect 8266 -7278 8272 -7244
rect 8226 -7316 8272 -7278
rect 8226 -7350 8232 -7316
rect 8266 -7350 8272 -7316
rect 8226 -7397 8272 -7350
rect 8484 -7244 8530 -7070
rect 8484 -7278 8490 -7244
rect 8524 -7278 8530 -7244
rect 8484 -7316 8530 -7278
rect 8484 -7350 8490 -7316
rect 8524 -7350 8530 -7316
rect 8484 -7397 8530 -7350
rect 8742 -7244 8788 -6769
rect 9000 -7000 9046 -6393
rect 9194 -6262 9573 -6228
rect 9607 -6262 9986 -6228
rect 13554 -6228 14344 -6193
rect 14547 -6129 15651 -6111
rect 14547 -6159 14597 -6129
rect 14547 -6193 14590 -6159
rect 14649 -6181 14661 -6129
rect 14713 -6181 14725 -6129
rect 14777 -6181 14793 -6129
rect 14845 -6159 14857 -6129
rect 14909 -6159 14921 -6129
rect 14845 -6181 14848 -6159
rect 14909 -6181 14920 -6159
rect 14973 -6181 15083 -6129
rect 15135 -6159 15147 -6129
rect 15199 -6159 15211 -6129
rect 15140 -6181 15147 -6159
rect 15263 -6181 15279 -6129
rect 15331 -6181 15343 -6129
rect 15395 -6159 15407 -6129
rect 15459 -6159 15651 -6129
rect 15398 -6181 15407 -6159
rect 14624 -6193 14662 -6181
rect 14696 -6193 14848 -6181
rect 14882 -6193 14920 -6181
rect 14954 -6193 15106 -6181
rect 15140 -6193 15178 -6181
rect 15212 -6193 15364 -6181
rect 15398 -6193 15436 -6181
rect 15470 -6193 15651 -6159
rect 14547 -6199 15651 -6193
rect 15773 -5990 16481 -5973
rect 15773 -6042 15811 -5990
rect 15863 -6042 15875 -5990
rect 15927 -6042 15939 -5990
rect 15991 -6042 16007 -5990
rect 16059 -6042 16071 -5990
rect 16123 -6042 16135 -5990
rect 16187 -6042 16199 -5990
rect 16251 -6042 16267 -5990
rect 16319 -6042 16331 -5990
rect 16383 -6042 16395 -5990
rect 16447 -6042 16481 -5990
rect 15773 -6159 16481 -6042
rect 15773 -6193 15816 -6159
rect 15850 -6193 15888 -6159
rect 15922 -6193 16074 -6159
rect 16108 -6193 16146 -6159
rect 16180 -6193 16332 -6159
rect 16366 -6193 16404 -6159
rect 16438 -6193 16481 -6159
rect 15773 -6199 16481 -6193
rect 16603 -6111 16664 -5879
rect 16741 -5797 17707 -5791
rect 16741 -5831 16784 -5797
rect 16818 -5812 16856 -5797
rect 16890 -5812 17042 -5797
rect 17076 -5812 17114 -5797
rect 17148 -5812 17300 -5797
rect 17334 -5812 17372 -5797
rect 17406 -5812 17558 -5797
rect 17592 -5812 17630 -5797
rect 16847 -5831 16856 -5812
rect 16741 -5864 16795 -5831
rect 16847 -5864 16859 -5831
rect 16911 -5864 16923 -5812
rect 16975 -5864 16991 -5812
rect 17107 -5831 17114 -5812
rect 17043 -5864 17055 -5831
rect 17107 -5864 17119 -5831
rect 17171 -5864 17281 -5812
rect 17334 -5831 17345 -5812
rect 17406 -5831 17409 -5812
rect 17333 -5864 17345 -5831
rect 17397 -5864 17409 -5831
rect 17461 -5864 17477 -5812
rect 17529 -5864 17541 -5812
rect 17593 -5864 17605 -5812
rect 17664 -5831 17707 -5797
rect 17657 -5864 17707 -5831
rect 16741 -5990 17707 -5864
rect 16741 -6042 16795 -5990
rect 16847 -6042 16859 -5990
rect 16911 -6042 16923 -5990
rect 16975 -6042 16991 -5990
rect 17043 -6042 17055 -5990
rect 17107 -6042 17119 -5990
rect 17171 -6042 17281 -5990
rect 17333 -6042 17345 -5990
rect 17397 -6042 17409 -5990
rect 17461 -6042 17477 -5990
rect 17529 -6042 17541 -5990
rect 17593 -6042 17605 -5990
rect 17657 -6042 17707 -5990
rect 16741 -6061 17707 -6042
rect 17911 -5796 18347 -5758
rect 17911 -5797 18290 -5796
rect 17911 -5831 18010 -5797
rect 18044 -5831 18082 -5797
rect 18116 -5830 18290 -5797
rect 18324 -5830 18347 -5796
rect 18116 -5831 18347 -5830
rect 17911 -5868 18347 -5831
rect 17911 -5902 18290 -5868
rect 18324 -5902 18347 -5868
rect 17911 -5940 18347 -5902
rect 17911 -5974 18290 -5940
rect 18324 -5974 18347 -5940
rect 17911 -6012 18347 -5974
rect 17911 -6046 18290 -6012
rect 18324 -6046 18347 -6012
rect 17911 -6084 18347 -6046
rect 16603 -6129 17707 -6111
rect 16603 -6159 16795 -6129
rect 16847 -6159 16859 -6129
rect 16603 -6193 16784 -6159
rect 16847 -6181 16856 -6159
rect 16911 -6181 16923 -6129
rect 16975 -6181 16991 -6129
rect 17043 -6159 17055 -6129
rect 17107 -6159 17119 -6129
rect 17107 -6181 17114 -6159
rect 17171 -6181 17281 -6129
rect 17333 -6159 17345 -6129
rect 17397 -6159 17409 -6129
rect 17334 -6181 17345 -6159
rect 17406 -6181 17409 -6159
rect 17461 -6181 17477 -6129
rect 17529 -6181 17541 -6129
rect 17593 -6181 17605 -6129
rect 17657 -6159 17707 -6129
rect 16818 -6193 16856 -6181
rect 16890 -6193 17042 -6181
rect 17076 -6193 17114 -6181
rect 17148 -6193 17300 -6181
rect 17334 -6193 17372 -6181
rect 17406 -6193 17558 -6181
rect 17592 -6193 17630 -6181
rect 17664 -6193 17707 -6159
rect 16603 -6199 17707 -6193
rect 17911 -6118 18290 -6084
rect 18324 -6118 18347 -6084
rect 17911 -6156 18347 -6118
rect 17911 -6159 18290 -6156
rect 17911 -6193 18010 -6159
rect 18044 -6193 18082 -6159
rect 18116 -6190 18290 -6159
rect 18324 -6190 18347 -6156
rect 18116 -6193 18347 -6190
rect 9194 -6287 9986 -6262
rect 9194 -6321 9200 -6287
rect 9234 -6321 9458 -6287
rect 9492 -6300 9688 -6287
rect 9492 -6321 9573 -6300
rect 9194 -6334 9573 -6321
rect 9607 -6321 9688 -6300
rect 9722 -6321 9946 -6287
rect 9980 -6321 9986 -6287
rect 9607 -6334 9986 -6321
rect 9194 -6359 9986 -6334
rect 9194 -6393 9200 -6359
rect 9234 -6393 9458 -6359
rect 9492 -6372 9688 -6359
rect 9492 -6393 9573 -6372
rect 9194 -6406 9573 -6393
rect 9607 -6393 9688 -6372
rect 9722 -6393 9946 -6359
rect 9980 -6393 9986 -6359
rect 9607 -6406 9986 -6393
rect 9194 -6444 9986 -6406
rect 9194 -6478 9573 -6444
rect 9607 -6478 9986 -6444
rect 9194 -6516 9986 -6478
rect 9194 -6550 9573 -6516
rect 9607 -6550 9986 -6516
rect 9194 -6588 9986 -6550
rect 9194 -6622 9573 -6588
rect 9607 -6622 9986 -6588
rect 9194 -6660 9986 -6622
rect 9194 -6694 9573 -6660
rect 9607 -6694 9986 -6660
rect 9194 -6732 9986 -6694
rect 9194 -6766 9573 -6732
rect 9607 -6766 9986 -6732
rect 9194 -6804 9986 -6766
rect 9194 -6838 9573 -6804
rect 9607 -6838 9986 -6804
rect 9194 -6876 9986 -6838
rect 9194 -6910 9573 -6876
rect 9607 -6910 9986 -6876
rect 9194 -6948 9986 -6910
rect 9194 -6982 9573 -6948
rect 9607 -6982 9986 -6948
rect 8923 -7010 9119 -7000
rect 8923 -7062 8932 -7010
rect 8984 -7062 8996 -7010
rect 9048 -7062 9060 -7010
rect 9112 -7062 9119 -7010
rect 8923 -7070 9119 -7062
rect 9194 -7020 9986 -6982
rect 10134 -6287 10180 -6240
rect 10134 -6321 10140 -6287
rect 10174 -6321 10180 -6287
rect 10134 -6359 10180 -6321
rect 10134 -6393 10140 -6359
rect 10174 -6393 10180 -6359
rect 10134 -7000 10180 -6393
rect 10392 -6287 10438 -6240
rect 10392 -6321 10398 -6287
rect 10432 -6321 10438 -6287
rect 10392 -6359 10438 -6321
rect 10392 -6393 10398 -6359
rect 10432 -6393 10438 -6359
rect 10392 -6699 10438 -6393
rect 10650 -6287 10696 -6240
rect 10650 -6321 10656 -6287
rect 10690 -6321 10696 -6287
rect 10650 -6359 10696 -6321
rect 10650 -6393 10656 -6359
rect 10690 -6393 10696 -6359
rect 10319 -6709 10515 -6699
rect 10319 -6761 10326 -6709
rect 10378 -6761 10390 -6709
rect 10442 -6761 10454 -6709
rect 10506 -6761 10515 -6709
rect 10319 -6769 10515 -6761
rect 9194 -7054 9573 -7020
rect 9607 -7054 9986 -7020
rect 8742 -7278 8748 -7244
rect 8782 -7278 8788 -7244
rect 8742 -7316 8788 -7278
rect 8742 -7350 8748 -7316
rect 8782 -7350 8788 -7316
rect 8742 -7397 8788 -7350
rect 9000 -7244 9046 -7070
rect 9000 -7278 9006 -7244
rect 9040 -7278 9046 -7244
rect 9000 -7316 9046 -7278
rect 9000 -7350 9006 -7316
rect 9040 -7350 9046 -7316
rect 9000 -7397 9046 -7350
rect 9194 -7092 9986 -7054
rect 10061 -7010 10257 -7000
rect 10061 -7062 10068 -7010
rect 10120 -7062 10132 -7010
rect 10184 -7062 10196 -7010
rect 10248 -7062 10257 -7010
rect 10061 -7070 10257 -7062
rect 9194 -7126 9573 -7092
rect 9607 -7126 9986 -7092
rect 9194 -7164 9986 -7126
rect 9194 -7198 9573 -7164
rect 9607 -7198 9986 -7164
rect 9194 -7236 9986 -7198
rect 9194 -7244 9573 -7236
rect 9194 -7278 9200 -7244
rect 9234 -7278 9458 -7244
rect 9492 -7270 9573 -7244
rect 9607 -7244 9986 -7236
rect 9607 -7270 9688 -7244
rect 9492 -7278 9688 -7270
rect 9722 -7278 9946 -7244
rect 9980 -7278 9986 -7244
rect 9194 -7308 9986 -7278
rect 9194 -7316 9573 -7308
rect 9194 -7350 9200 -7316
rect 9234 -7350 9458 -7316
rect 9492 -7342 9573 -7316
rect 9607 -7316 9986 -7308
rect 9607 -7342 9688 -7316
rect 9492 -7350 9688 -7342
rect 9722 -7350 9946 -7316
rect 9980 -7350 9986 -7316
rect 9194 -7380 9986 -7350
rect 833 -7452 1064 -7444
rect 833 -7486 856 -7452
rect 890 -7478 1064 -7452
rect 1098 -7478 1136 -7444
rect 1170 -7478 1269 -7444
rect 890 -7486 1269 -7478
rect 833 -7524 1269 -7486
rect 833 -7558 856 -7524
rect 890 -7558 1269 -7524
rect 833 -7596 1269 -7558
rect 833 -7630 856 -7596
rect 890 -7630 1269 -7596
rect 833 -7668 1269 -7630
rect 833 -7702 856 -7668
rect 890 -7702 1269 -7668
rect 833 -7740 1269 -7702
rect 1473 -7444 2439 -7438
rect 1473 -7478 1516 -7444
rect 1550 -7459 1588 -7444
rect 1622 -7459 1774 -7444
rect 1808 -7459 1846 -7444
rect 1880 -7459 2032 -7444
rect 2066 -7459 2104 -7444
rect 2138 -7459 2290 -7444
rect 2324 -7459 2362 -7444
rect 1473 -7511 1523 -7478
rect 1575 -7511 1587 -7459
rect 1639 -7511 1651 -7459
rect 1703 -7511 1719 -7459
rect 1771 -7478 1774 -7459
rect 1835 -7478 1846 -7459
rect 1771 -7511 1783 -7478
rect 1835 -7511 1847 -7478
rect 1899 -7511 2009 -7459
rect 2066 -7478 2073 -7459
rect 2061 -7511 2073 -7478
rect 2125 -7511 2137 -7478
rect 2189 -7511 2205 -7459
rect 2257 -7511 2269 -7459
rect 2324 -7478 2333 -7459
rect 2396 -7478 2439 -7444
rect 2321 -7511 2333 -7478
rect 2385 -7511 2439 -7478
rect 1473 -7637 2439 -7511
rect 1473 -7689 1523 -7637
rect 1575 -7689 1587 -7637
rect 1639 -7689 1651 -7637
rect 1703 -7689 1719 -7637
rect 1771 -7689 1783 -7637
rect 1835 -7689 1847 -7637
rect 1899 -7689 2009 -7637
rect 2061 -7689 2073 -7637
rect 2125 -7689 2137 -7637
rect 2189 -7689 2205 -7637
rect 2257 -7689 2269 -7637
rect 2321 -7689 2333 -7637
rect 2385 -7689 2439 -7637
rect 1473 -7708 2439 -7689
rect 2516 -7444 3590 -7438
rect 2516 -7478 2742 -7444
rect 2776 -7478 2814 -7444
rect 2848 -7478 3000 -7444
rect 3034 -7478 3072 -7444
rect 3106 -7478 3258 -7444
rect 3292 -7478 3330 -7444
rect 3364 -7478 3590 -7444
rect 2516 -7526 3590 -7478
rect 833 -7774 856 -7740
rect 890 -7774 1269 -7740
rect 2516 -7758 2577 -7526
rect 833 -7806 1269 -7774
rect 833 -7812 1064 -7806
rect 833 -7846 856 -7812
rect 890 -7840 1064 -7812
rect 1098 -7840 1136 -7806
rect 1170 -7840 1269 -7806
rect 890 -7846 1269 -7840
rect 1473 -7776 2577 -7758
rect 1473 -7806 1523 -7776
rect 1473 -7840 1516 -7806
rect 1575 -7828 1587 -7776
rect 1639 -7828 1651 -7776
rect 1703 -7828 1719 -7776
rect 1771 -7806 1783 -7776
rect 1835 -7806 1847 -7776
rect 1771 -7828 1774 -7806
rect 1835 -7828 1846 -7806
rect 1899 -7828 2009 -7776
rect 2061 -7806 2073 -7776
rect 2125 -7806 2137 -7776
rect 2066 -7828 2073 -7806
rect 2189 -7828 2205 -7776
rect 2257 -7828 2269 -7776
rect 2321 -7806 2333 -7776
rect 2385 -7806 2577 -7776
rect 2324 -7828 2333 -7806
rect 1550 -7840 1588 -7828
rect 1622 -7840 1774 -7828
rect 1808 -7840 1846 -7828
rect 1880 -7840 2032 -7828
rect 2066 -7840 2104 -7828
rect 2138 -7840 2290 -7828
rect 2324 -7840 2362 -7828
rect 2396 -7840 2577 -7806
rect 1473 -7846 2577 -7840
rect 2699 -7637 3407 -7620
rect 2699 -7689 2733 -7637
rect 2785 -7689 2797 -7637
rect 2849 -7689 2861 -7637
rect 2913 -7689 2929 -7637
rect 2981 -7689 2993 -7637
rect 3045 -7689 3057 -7637
rect 3109 -7689 3121 -7637
rect 3173 -7689 3189 -7637
rect 3241 -7689 3253 -7637
rect 3305 -7689 3317 -7637
rect 3369 -7689 3407 -7637
rect 2699 -7806 3407 -7689
rect 2699 -7840 2742 -7806
rect 2776 -7840 2814 -7806
rect 2848 -7840 3000 -7806
rect 3034 -7840 3072 -7806
rect 3106 -7840 3258 -7806
rect 3292 -7840 3330 -7806
rect 3364 -7840 3407 -7806
rect 2699 -7846 3407 -7840
rect 3529 -7758 3590 -7526
rect 3667 -7444 4633 -7438
rect 3667 -7478 3710 -7444
rect 3744 -7459 3782 -7444
rect 3816 -7459 3968 -7444
rect 4002 -7459 4040 -7444
rect 4074 -7459 4226 -7444
rect 4260 -7459 4298 -7444
rect 4332 -7459 4484 -7444
rect 4518 -7459 4556 -7444
rect 3773 -7478 3782 -7459
rect 3667 -7511 3721 -7478
rect 3773 -7511 3785 -7478
rect 3837 -7511 3849 -7459
rect 3901 -7511 3917 -7459
rect 4033 -7478 4040 -7459
rect 3969 -7511 3981 -7478
rect 4033 -7511 4045 -7478
rect 4097 -7511 4207 -7459
rect 4260 -7478 4271 -7459
rect 4332 -7478 4335 -7459
rect 4259 -7511 4271 -7478
rect 4323 -7511 4335 -7478
rect 4387 -7511 4403 -7459
rect 4455 -7511 4467 -7459
rect 4519 -7511 4531 -7459
rect 4590 -7478 4633 -7444
rect 4583 -7511 4633 -7478
rect 3667 -7637 4633 -7511
rect 3667 -7689 3721 -7637
rect 3773 -7689 3785 -7637
rect 3837 -7689 3849 -7637
rect 3901 -7689 3917 -7637
rect 3969 -7689 3981 -7637
rect 4033 -7689 4045 -7637
rect 4097 -7689 4207 -7637
rect 4259 -7689 4271 -7637
rect 4323 -7689 4335 -7637
rect 4387 -7689 4403 -7637
rect 4455 -7689 4467 -7637
rect 4519 -7689 4531 -7637
rect 4583 -7689 4633 -7637
rect 3667 -7708 4633 -7689
rect 4836 -7444 5626 -7414
rect 9194 -7414 9573 -7380
rect 9607 -7414 9986 -7380
rect 10134 -7244 10180 -7070
rect 10134 -7278 10140 -7244
rect 10174 -7278 10180 -7244
rect 10134 -7316 10180 -7278
rect 10134 -7350 10140 -7316
rect 10174 -7350 10180 -7316
rect 10134 -7397 10180 -7350
rect 10392 -7244 10438 -6769
rect 10650 -7000 10696 -6393
rect 10908 -6287 10954 -6240
rect 10908 -6321 10914 -6287
rect 10948 -6321 10954 -6287
rect 10908 -6359 10954 -6321
rect 10908 -6393 10914 -6359
rect 10948 -6393 10954 -6359
rect 10908 -6699 10954 -6393
rect 11166 -6287 11212 -6240
rect 11166 -6321 11172 -6287
rect 11206 -6321 11212 -6287
rect 11166 -6359 11212 -6321
rect 11166 -6393 11172 -6359
rect 11206 -6393 11212 -6359
rect 10836 -6709 11032 -6699
rect 10836 -6761 10843 -6709
rect 10895 -6761 10907 -6709
rect 10959 -6761 10971 -6709
rect 11023 -6761 11032 -6709
rect 10836 -6769 11032 -6761
rect 10576 -7010 10772 -7000
rect 10576 -7062 10583 -7010
rect 10635 -7062 10647 -7010
rect 10699 -7062 10711 -7010
rect 10763 -7062 10772 -7010
rect 10576 -7070 10772 -7062
rect 10392 -7278 10398 -7244
rect 10432 -7278 10438 -7244
rect 10392 -7316 10438 -7278
rect 10392 -7350 10398 -7316
rect 10432 -7350 10438 -7316
rect 10392 -7397 10438 -7350
rect 10650 -7244 10696 -7070
rect 10650 -7278 10656 -7244
rect 10690 -7278 10696 -7244
rect 10650 -7316 10696 -7278
rect 10650 -7350 10656 -7316
rect 10690 -7350 10696 -7316
rect 10650 -7397 10696 -7350
rect 10908 -7244 10954 -6769
rect 11166 -7000 11212 -6393
rect 11360 -6287 11406 -6240
rect 11360 -6321 11366 -6287
rect 11400 -6321 11406 -6287
rect 11360 -6359 11406 -6321
rect 11360 -6393 11366 -6359
rect 11400 -6393 11406 -6359
rect 11360 -6554 11406 -6393
rect 11618 -6287 11664 -6240
rect 11618 -6321 11624 -6287
rect 11658 -6321 11664 -6287
rect 11618 -6359 11664 -6321
rect 11618 -6393 11624 -6359
rect 11658 -6393 11664 -6359
rect 11283 -6564 11479 -6554
rect 11283 -6616 11292 -6564
rect 11344 -6616 11356 -6564
rect 11408 -6616 11420 -6564
rect 11472 -6616 11479 -6564
rect 11283 -6624 11479 -6616
rect 11093 -7010 11289 -7000
rect 11093 -7062 11100 -7010
rect 11152 -7062 11164 -7010
rect 11216 -7062 11228 -7010
rect 11280 -7062 11289 -7010
rect 11093 -7070 11289 -7062
rect 10908 -7278 10914 -7244
rect 10948 -7278 10954 -7244
rect 10908 -7316 10954 -7278
rect 10908 -7350 10914 -7316
rect 10948 -7350 10954 -7316
rect 10908 -7397 10954 -7350
rect 11166 -7244 11212 -7070
rect 11166 -7278 11172 -7244
rect 11206 -7278 11212 -7244
rect 11166 -7316 11212 -7278
rect 11166 -7350 11172 -7316
rect 11206 -7350 11212 -7316
rect 11166 -7397 11212 -7350
rect 11360 -7244 11406 -6624
rect 11618 -6860 11664 -6393
rect 11876 -6287 11922 -6240
rect 11876 -6321 11882 -6287
rect 11916 -6321 11922 -6287
rect 11876 -6359 11922 -6321
rect 11876 -6393 11882 -6359
rect 11916 -6393 11922 -6359
rect 11876 -6554 11922 -6393
rect 12134 -6287 12180 -6240
rect 12134 -6321 12140 -6287
rect 12174 -6321 12180 -6287
rect 12134 -6359 12180 -6321
rect 12134 -6393 12140 -6359
rect 12174 -6393 12180 -6359
rect 11800 -6564 11996 -6554
rect 11800 -6616 11809 -6564
rect 11861 -6616 11873 -6564
rect 11925 -6616 11937 -6564
rect 11989 -6616 11996 -6564
rect 11800 -6624 11996 -6616
rect 11541 -6870 11737 -6860
rect 11541 -6922 11550 -6870
rect 11602 -6922 11614 -6870
rect 11666 -6922 11678 -6870
rect 11730 -6922 11737 -6870
rect 11541 -6930 11737 -6922
rect 11360 -7278 11366 -7244
rect 11400 -7278 11406 -7244
rect 11360 -7316 11406 -7278
rect 11360 -7350 11366 -7316
rect 11400 -7350 11406 -7316
rect 11360 -7397 11406 -7350
rect 11618 -7244 11664 -6930
rect 11618 -7278 11624 -7244
rect 11658 -7278 11664 -7244
rect 11618 -7316 11664 -7278
rect 11618 -7350 11624 -7316
rect 11658 -7350 11664 -7316
rect 11618 -7397 11664 -7350
rect 11876 -7244 11922 -6624
rect 12134 -6860 12180 -6393
rect 12328 -6287 12374 -6240
rect 12328 -6321 12334 -6287
rect 12368 -6321 12374 -6287
rect 12328 -6359 12374 -6321
rect 12328 -6393 12334 -6359
rect 12368 -6393 12374 -6359
rect 12058 -6870 12254 -6860
rect 12058 -6922 12067 -6870
rect 12119 -6922 12131 -6870
rect 12183 -6922 12195 -6870
rect 12247 -6922 12254 -6870
rect 12058 -6930 12254 -6922
rect 11876 -7278 11882 -7244
rect 11916 -7278 11922 -7244
rect 11876 -7316 11922 -7278
rect 11876 -7350 11882 -7316
rect 11916 -7350 11922 -7316
rect 11876 -7397 11922 -7350
rect 12134 -7244 12180 -6930
rect 12328 -7000 12374 -6393
rect 12586 -6287 12632 -6240
rect 12586 -6321 12592 -6287
rect 12626 -6321 12632 -6287
rect 12586 -6359 12632 -6321
rect 12586 -6393 12592 -6359
rect 12626 -6393 12632 -6359
rect 12586 -6699 12632 -6393
rect 12844 -6287 12890 -6240
rect 12844 -6321 12850 -6287
rect 12884 -6321 12890 -6287
rect 12844 -6359 12890 -6321
rect 12844 -6393 12850 -6359
rect 12884 -6393 12890 -6359
rect 12513 -6709 12709 -6699
rect 12513 -6761 12520 -6709
rect 12572 -6761 12584 -6709
rect 12636 -6761 12648 -6709
rect 12700 -6761 12709 -6709
rect 12513 -6769 12709 -6761
rect 12253 -7010 12449 -7000
rect 12253 -7062 12260 -7010
rect 12312 -7062 12324 -7010
rect 12376 -7062 12388 -7010
rect 12440 -7062 12449 -7010
rect 12253 -7070 12449 -7062
rect 12134 -7278 12140 -7244
rect 12174 -7278 12180 -7244
rect 12134 -7316 12180 -7278
rect 12134 -7350 12140 -7316
rect 12174 -7350 12180 -7316
rect 12134 -7397 12180 -7350
rect 12328 -7244 12374 -7070
rect 12328 -7278 12334 -7244
rect 12368 -7278 12374 -7244
rect 12328 -7316 12374 -7278
rect 12328 -7350 12334 -7316
rect 12368 -7350 12374 -7316
rect 12328 -7397 12374 -7350
rect 12586 -7244 12632 -6769
rect 12844 -7000 12890 -6393
rect 13102 -6287 13148 -6240
rect 13102 -6321 13108 -6287
rect 13142 -6321 13148 -6287
rect 13102 -6359 13148 -6321
rect 13102 -6393 13108 -6359
rect 13142 -6393 13148 -6359
rect 13102 -6699 13148 -6393
rect 13360 -6287 13406 -6240
rect 13360 -6321 13366 -6287
rect 13400 -6321 13406 -6287
rect 13360 -6359 13406 -6321
rect 13360 -6393 13366 -6359
rect 13400 -6393 13406 -6359
rect 13030 -6709 13226 -6699
rect 13030 -6761 13037 -6709
rect 13089 -6761 13101 -6709
rect 13153 -6761 13165 -6709
rect 13217 -6761 13226 -6709
rect 13030 -6769 13226 -6761
rect 12770 -7010 12966 -7000
rect 12770 -7062 12777 -7010
rect 12829 -7062 12841 -7010
rect 12893 -7062 12905 -7010
rect 12957 -7062 12966 -7010
rect 12770 -7070 12966 -7062
rect 12586 -7278 12592 -7244
rect 12626 -7278 12632 -7244
rect 12586 -7316 12632 -7278
rect 12586 -7350 12592 -7316
rect 12626 -7350 12632 -7316
rect 12586 -7397 12632 -7350
rect 12844 -7244 12890 -7070
rect 12844 -7278 12850 -7244
rect 12884 -7278 12890 -7244
rect 12844 -7316 12890 -7278
rect 12844 -7350 12850 -7316
rect 12884 -7350 12890 -7316
rect 12844 -7397 12890 -7350
rect 13102 -7244 13148 -6769
rect 13360 -7000 13406 -6393
rect 13554 -6262 13932 -6228
rect 13966 -6262 14344 -6228
rect 17911 -6228 18347 -6193
rect 13554 -6287 14344 -6262
rect 13554 -6321 13560 -6287
rect 13594 -6321 13818 -6287
rect 13852 -6300 14046 -6287
rect 13852 -6321 13932 -6300
rect 13554 -6334 13932 -6321
rect 13966 -6321 14046 -6300
rect 14080 -6321 14304 -6287
rect 14338 -6321 14344 -6287
rect 13966 -6334 14344 -6321
rect 13554 -6359 14344 -6334
rect 13554 -6393 13560 -6359
rect 13594 -6393 13818 -6359
rect 13852 -6372 14046 -6359
rect 13852 -6393 13932 -6372
rect 13554 -6406 13932 -6393
rect 13966 -6393 14046 -6372
rect 14080 -6393 14304 -6359
rect 14338 -6393 14344 -6359
rect 13966 -6406 14344 -6393
rect 13554 -6444 14344 -6406
rect 13554 -6478 13932 -6444
rect 13966 -6478 14344 -6444
rect 13554 -6516 14344 -6478
rect 13554 -6550 13932 -6516
rect 13966 -6550 14344 -6516
rect 13554 -6588 14344 -6550
rect 13554 -6622 13932 -6588
rect 13966 -6622 14344 -6588
rect 13554 -6660 14344 -6622
rect 13554 -6694 13932 -6660
rect 13966 -6694 14344 -6660
rect 13554 -6732 14344 -6694
rect 13554 -6766 13932 -6732
rect 13966 -6766 14344 -6732
rect 13554 -6804 14344 -6766
rect 13554 -6838 13932 -6804
rect 13966 -6838 14344 -6804
rect 13554 -6876 14344 -6838
rect 13554 -6910 13932 -6876
rect 13966 -6910 14344 -6876
rect 13554 -6948 14344 -6910
rect 13554 -6982 13932 -6948
rect 13966 -6982 14344 -6948
rect 13287 -7010 13483 -7000
rect 13287 -7062 13294 -7010
rect 13346 -7062 13358 -7010
rect 13410 -7062 13422 -7010
rect 13474 -7062 13483 -7010
rect 13287 -7070 13483 -7062
rect 13554 -7020 14344 -6982
rect 14491 -6287 14537 -6240
rect 14491 -6321 14497 -6287
rect 14531 -6321 14537 -6287
rect 14491 -6359 14537 -6321
rect 14491 -6393 14497 -6359
rect 14531 -6393 14537 -6359
rect 14491 -7000 14537 -6393
rect 14749 -6287 14795 -6240
rect 14749 -6321 14755 -6287
rect 14789 -6321 14795 -6287
rect 14749 -6359 14795 -6321
rect 14749 -6393 14755 -6359
rect 14789 -6393 14795 -6359
rect 14749 -6699 14795 -6393
rect 15007 -6287 15053 -6240
rect 15007 -6321 15013 -6287
rect 15047 -6321 15053 -6287
rect 15007 -6359 15053 -6321
rect 15007 -6393 15013 -6359
rect 15047 -6393 15053 -6359
rect 14671 -6709 14867 -6699
rect 14671 -6761 14680 -6709
rect 14732 -6761 14744 -6709
rect 14796 -6761 14808 -6709
rect 14860 -6761 14867 -6709
rect 14671 -6769 14867 -6761
rect 13554 -7054 13932 -7020
rect 13966 -7054 14344 -7020
rect 13102 -7278 13108 -7244
rect 13142 -7278 13148 -7244
rect 13102 -7316 13148 -7278
rect 13102 -7350 13108 -7316
rect 13142 -7350 13148 -7316
rect 13102 -7397 13148 -7350
rect 13360 -7244 13406 -7070
rect 13360 -7278 13366 -7244
rect 13400 -7278 13406 -7244
rect 13360 -7316 13406 -7278
rect 13360 -7350 13366 -7316
rect 13400 -7350 13406 -7316
rect 13360 -7397 13406 -7350
rect 13554 -7092 14344 -7054
rect 14414 -7010 14610 -7000
rect 14414 -7062 14423 -7010
rect 14475 -7062 14487 -7010
rect 14539 -7062 14551 -7010
rect 14603 -7062 14610 -7010
rect 14414 -7070 14610 -7062
rect 13554 -7126 13932 -7092
rect 13966 -7126 14344 -7092
rect 13554 -7164 14344 -7126
rect 13554 -7198 13932 -7164
rect 13966 -7198 14344 -7164
rect 13554 -7236 14344 -7198
rect 13554 -7244 13932 -7236
rect 13554 -7278 13560 -7244
rect 13594 -7278 13818 -7244
rect 13852 -7270 13932 -7244
rect 13966 -7244 14344 -7236
rect 13966 -7270 14046 -7244
rect 13852 -7278 14046 -7270
rect 14080 -7278 14304 -7244
rect 14338 -7278 14344 -7244
rect 13554 -7308 14344 -7278
rect 13554 -7316 13932 -7308
rect 13554 -7350 13560 -7316
rect 13594 -7350 13818 -7316
rect 13852 -7342 13932 -7316
rect 13966 -7316 14344 -7308
rect 13966 -7342 14046 -7316
rect 13852 -7350 14046 -7342
rect 14080 -7350 14304 -7316
rect 14338 -7350 14344 -7316
rect 13554 -7380 14344 -7350
rect 4836 -7478 4935 -7444
rect 4969 -7478 5007 -7444
rect 5041 -7452 5421 -7444
rect 5041 -7478 5214 -7452
rect 4836 -7486 5214 -7478
rect 5248 -7478 5421 -7452
rect 5455 -7478 5493 -7444
rect 5527 -7478 5626 -7444
rect 5248 -7486 5626 -7478
rect 4836 -7524 5626 -7486
rect 4836 -7558 5214 -7524
rect 5248 -7558 5626 -7524
rect 4836 -7596 5626 -7558
rect 4836 -7630 5214 -7596
rect 5248 -7630 5626 -7596
rect 4836 -7668 5626 -7630
rect 4836 -7702 5214 -7668
rect 5248 -7702 5626 -7668
rect 4836 -7740 5626 -7702
rect 5830 -7444 6796 -7438
rect 5830 -7478 5873 -7444
rect 5907 -7459 5945 -7444
rect 5979 -7459 6131 -7444
rect 6165 -7459 6203 -7444
rect 6237 -7459 6389 -7444
rect 6423 -7459 6461 -7444
rect 6495 -7459 6647 -7444
rect 6681 -7459 6719 -7444
rect 5830 -7511 5880 -7478
rect 5932 -7511 5944 -7459
rect 5996 -7511 6008 -7459
rect 6060 -7511 6076 -7459
rect 6128 -7478 6131 -7459
rect 6192 -7478 6203 -7459
rect 6128 -7511 6140 -7478
rect 6192 -7511 6204 -7478
rect 6256 -7511 6366 -7459
rect 6423 -7478 6430 -7459
rect 6418 -7511 6430 -7478
rect 6482 -7511 6494 -7478
rect 6546 -7511 6562 -7459
rect 6614 -7511 6626 -7459
rect 6681 -7478 6690 -7459
rect 6753 -7478 6796 -7444
rect 6678 -7511 6690 -7478
rect 6742 -7511 6796 -7478
rect 5830 -7637 6796 -7511
rect 5830 -7689 5880 -7637
rect 5932 -7689 5944 -7637
rect 5996 -7689 6008 -7637
rect 6060 -7689 6076 -7637
rect 6128 -7689 6140 -7637
rect 6192 -7689 6204 -7637
rect 6256 -7689 6366 -7637
rect 6418 -7689 6430 -7637
rect 6482 -7689 6494 -7637
rect 6546 -7689 6562 -7637
rect 6614 -7689 6626 -7637
rect 6678 -7689 6690 -7637
rect 6742 -7689 6796 -7637
rect 5830 -7708 6796 -7689
rect 6873 -7444 7947 -7438
rect 6873 -7478 7099 -7444
rect 7133 -7478 7171 -7444
rect 7205 -7478 7357 -7444
rect 7391 -7478 7429 -7444
rect 7463 -7478 7615 -7444
rect 7649 -7478 7687 -7444
rect 7721 -7478 7947 -7444
rect 6873 -7526 7947 -7478
rect 3529 -7776 4633 -7758
rect 3529 -7806 3721 -7776
rect 3773 -7806 3785 -7776
rect 3529 -7840 3710 -7806
rect 3773 -7828 3782 -7806
rect 3837 -7828 3849 -7776
rect 3901 -7828 3917 -7776
rect 3969 -7806 3981 -7776
rect 4033 -7806 4045 -7776
rect 4033 -7828 4040 -7806
rect 4097 -7828 4207 -7776
rect 4259 -7806 4271 -7776
rect 4323 -7806 4335 -7776
rect 4260 -7828 4271 -7806
rect 4332 -7828 4335 -7806
rect 4387 -7828 4403 -7776
rect 4455 -7828 4467 -7776
rect 4519 -7828 4531 -7776
rect 4583 -7806 4633 -7776
rect 3744 -7840 3782 -7828
rect 3816 -7840 3968 -7828
rect 4002 -7840 4040 -7828
rect 4074 -7840 4226 -7828
rect 4260 -7840 4298 -7828
rect 4332 -7840 4484 -7828
rect 4518 -7840 4556 -7828
rect 4590 -7840 4633 -7806
rect 3529 -7846 4633 -7840
rect 4836 -7774 5214 -7740
rect 5248 -7774 5626 -7740
rect 6873 -7758 6934 -7526
rect 4836 -7806 5626 -7774
rect 4836 -7840 4935 -7806
rect 4969 -7840 5007 -7806
rect 5041 -7812 5421 -7806
rect 5041 -7840 5214 -7812
rect 4836 -7846 5214 -7840
rect 5248 -7840 5421 -7812
rect 5455 -7840 5493 -7806
rect 5527 -7840 5626 -7806
rect 5248 -7846 5626 -7840
rect 5830 -7776 6934 -7758
rect 5830 -7806 5880 -7776
rect 5830 -7840 5873 -7806
rect 5932 -7828 5944 -7776
rect 5996 -7828 6008 -7776
rect 6060 -7828 6076 -7776
rect 6128 -7806 6140 -7776
rect 6192 -7806 6204 -7776
rect 6128 -7828 6131 -7806
rect 6192 -7828 6203 -7806
rect 6256 -7828 6366 -7776
rect 6418 -7806 6430 -7776
rect 6482 -7806 6494 -7776
rect 6423 -7828 6430 -7806
rect 6546 -7828 6562 -7776
rect 6614 -7828 6626 -7776
rect 6678 -7806 6690 -7776
rect 6742 -7806 6934 -7776
rect 6681 -7828 6690 -7806
rect 5907 -7840 5945 -7828
rect 5979 -7840 6131 -7828
rect 6165 -7840 6203 -7828
rect 6237 -7840 6389 -7828
rect 6423 -7840 6461 -7828
rect 6495 -7840 6647 -7828
rect 6681 -7840 6719 -7828
rect 6753 -7840 6934 -7806
rect 5830 -7846 6934 -7840
rect 7056 -7637 7764 -7620
rect 7056 -7689 7094 -7637
rect 7146 -7689 7158 -7637
rect 7210 -7689 7222 -7637
rect 7274 -7689 7290 -7637
rect 7342 -7689 7354 -7637
rect 7406 -7689 7418 -7637
rect 7470 -7689 7482 -7637
rect 7534 -7689 7550 -7637
rect 7602 -7689 7614 -7637
rect 7666 -7689 7678 -7637
rect 7730 -7689 7764 -7637
rect 7056 -7806 7764 -7689
rect 7056 -7840 7099 -7806
rect 7133 -7840 7171 -7806
rect 7205 -7840 7357 -7806
rect 7391 -7840 7429 -7806
rect 7463 -7840 7615 -7806
rect 7649 -7840 7687 -7806
rect 7721 -7840 7764 -7806
rect 7056 -7846 7764 -7840
rect 7886 -7758 7947 -7526
rect 8024 -7444 8990 -7438
rect 8024 -7478 8067 -7444
rect 8101 -7459 8139 -7444
rect 8173 -7459 8325 -7444
rect 8359 -7459 8397 -7444
rect 8431 -7459 8583 -7444
rect 8617 -7459 8655 -7444
rect 8689 -7459 8841 -7444
rect 8875 -7459 8913 -7444
rect 8130 -7478 8139 -7459
rect 8024 -7511 8078 -7478
rect 8130 -7511 8142 -7478
rect 8194 -7511 8206 -7459
rect 8258 -7511 8274 -7459
rect 8390 -7478 8397 -7459
rect 8326 -7511 8338 -7478
rect 8390 -7511 8402 -7478
rect 8454 -7511 8564 -7459
rect 8617 -7478 8628 -7459
rect 8689 -7478 8692 -7459
rect 8616 -7511 8628 -7478
rect 8680 -7511 8692 -7478
rect 8744 -7511 8760 -7459
rect 8812 -7511 8824 -7459
rect 8876 -7511 8888 -7459
rect 8947 -7478 8990 -7444
rect 8940 -7511 8990 -7478
rect 8024 -7637 8990 -7511
rect 8024 -7689 8078 -7637
rect 8130 -7689 8142 -7637
rect 8194 -7689 8206 -7637
rect 8258 -7689 8274 -7637
rect 8326 -7689 8338 -7637
rect 8390 -7689 8402 -7637
rect 8454 -7689 8564 -7637
rect 8616 -7689 8628 -7637
rect 8680 -7689 8692 -7637
rect 8744 -7689 8760 -7637
rect 8812 -7689 8824 -7637
rect 8876 -7689 8888 -7637
rect 8940 -7689 8990 -7637
rect 8024 -7708 8990 -7689
rect 9194 -7444 9986 -7414
rect 13554 -7414 13932 -7380
rect 13966 -7414 14344 -7380
rect 14491 -7244 14537 -7070
rect 14491 -7278 14497 -7244
rect 14531 -7278 14537 -7244
rect 14491 -7316 14537 -7278
rect 14491 -7350 14497 -7316
rect 14531 -7350 14537 -7316
rect 14491 -7397 14537 -7350
rect 14749 -7244 14795 -6769
rect 15007 -7000 15053 -6393
rect 15265 -6287 15311 -6240
rect 15265 -6321 15271 -6287
rect 15305 -6321 15311 -6287
rect 15265 -6359 15311 -6321
rect 15265 -6393 15271 -6359
rect 15305 -6393 15311 -6359
rect 15265 -6699 15311 -6393
rect 15523 -6287 15569 -6240
rect 15523 -6321 15529 -6287
rect 15563 -6321 15569 -6287
rect 15523 -6359 15569 -6321
rect 15523 -6393 15529 -6359
rect 15563 -6393 15569 -6359
rect 15188 -6709 15384 -6699
rect 15188 -6761 15197 -6709
rect 15249 -6761 15261 -6709
rect 15313 -6761 15325 -6709
rect 15377 -6761 15384 -6709
rect 15188 -6769 15384 -6761
rect 14931 -7010 15127 -7000
rect 14931 -7062 14940 -7010
rect 14992 -7062 15004 -7010
rect 15056 -7062 15068 -7010
rect 15120 -7062 15127 -7010
rect 14931 -7070 15127 -7062
rect 14749 -7278 14755 -7244
rect 14789 -7278 14795 -7244
rect 14749 -7316 14795 -7278
rect 14749 -7350 14755 -7316
rect 14789 -7350 14795 -7316
rect 14749 -7397 14795 -7350
rect 15007 -7244 15053 -7070
rect 15007 -7278 15013 -7244
rect 15047 -7278 15053 -7244
rect 15007 -7316 15053 -7278
rect 15007 -7350 15013 -7316
rect 15047 -7350 15053 -7316
rect 15007 -7397 15053 -7350
rect 15265 -7244 15311 -6769
rect 15523 -7000 15569 -6393
rect 15717 -6287 15763 -6240
rect 15717 -6321 15723 -6287
rect 15757 -6321 15763 -6287
rect 15717 -6359 15763 -6321
rect 15717 -6393 15723 -6359
rect 15757 -6393 15763 -6359
rect 15717 -6860 15763 -6393
rect 15975 -6287 16021 -6240
rect 15975 -6321 15981 -6287
rect 16015 -6321 16021 -6287
rect 15975 -6359 16021 -6321
rect 15975 -6393 15981 -6359
rect 16015 -6393 16021 -6359
rect 15975 -6554 16021 -6393
rect 16233 -6287 16279 -6240
rect 16233 -6321 16239 -6287
rect 16273 -6321 16279 -6287
rect 16233 -6359 16279 -6321
rect 16233 -6393 16239 -6359
rect 16273 -6393 16279 -6359
rect 15901 -6564 16097 -6554
rect 15901 -6616 15908 -6564
rect 15960 -6616 15972 -6564
rect 16024 -6616 16036 -6564
rect 16088 -6616 16097 -6564
rect 15901 -6624 16097 -6616
rect 15643 -6870 15839 -6860
rect 15643 -6922 15650 -6870
rect 15702 -6922 15714 -6870
rect 15766 -6922 15778 -6870
rect 15830 -6922 15839 -6870
rect 15643 -6930 15839 -6922
rect 15448 -7010 15644 -7000
rect 15448 -7062 15457 -7010
rect 15509 -7062 15521 -7010
rect 15573 -7062 15585 -7010
rect 15637 -7062 15644 -7010
rect 15448 -7070 15644 -7062
rect 15265 -7278 15271 -7244
rect 15305 -7278 15311 -7244
rect 15265 -7316 15311 -7278
rect 15265 -7350 15271 -7316
rect 15305 -7350 15311 -7316
rect 15265 -7397 15311 -7350
rect 15523 -7244 15569 -7070
rect 15523 -7278 15529 -7244
rect 15563 -7278 15569 -7244
rect 15523 -7316 15569 -7278
rect 15523 -7350 15529 -7316
rect 15563 -7350 15569 -7316
rect 15523 -7397 15569 -7350
rect 15717 -7244 15763 -6930
rect 15717 -7278 15723 -7244
rect 15757 -7278 15763 -7244
rect 15717 -7316 15763 -7278
rect 15717 -7350 15723 -7316
rect 15757 -7350 15763 -7316
rect 15717 -7397 15763 -7350
rect 15975 -7244 16021 -6624
rect 16233 -6860 16279 -6393
rect 16491 -6287 16537 -6240
rect 16491 -6321 16497 -6287
rect 16531 -6321 16537 -6287
rect 16491 -6359 16537 -6321
rect 16491 -6393 16497 -6359
rect 16531 -6393 16537 -6359
rect 16491 -6554 16537 -6393
rect 16685 -6287 16731 -6240
rect 16685 -6321 16691 -6287
rect 16725 -6321 16731 -6287
rect 16685 -6359 16731 -6321
rect 16685 -6393 16691 -6359
rect 16725 -6393 16731 -6359
rect 16418 -6564 16614 -6554
rect 16418 -6616 16425 -6564
rect 16477 -6616 16489 -6564
rect 16541 -6616 16553 -6564
rect 16605 -6616 16614 -6564
rect 16418 -6624 16614 -6616
rect 16160 -6870 16356 -6860
rect 16160 -6922 16167 -6870
rect 16219 -6922 16231 -6870
rect 16283 -6922 16295 -6870
rect 16347 -6922 16356 -6870
rect 16160 -6930 16356 -6922
rect 15975 -7278 15981 -7244
rect 16015 -7278 16021 -7244
rect 15975 -7316 16021 -7278
rect 15975 -7350 15981 -7316
rect 16015 -7350 16021 -7316
rect 15975 -7397 16021 -7350
rect 16233 -7244 16279 -6930
rect 16233 -7278 16239 -7244
rect 16273 -7278 16279 -7244
rect 16233 -7316 16279 -7278
rect 16233 -7350 16239 -7316
rect 16273 -7350 16279 -7316
rect 16233 -7397 16279 -7350
rect 16491 -7244 16537 -6624
rect 16685 -7000 16731 -6393
rect 16943 -6287 16989 -6240
rect 16943 -6321 16949 -6287
rect 16983 -6321 16989 -6287
rect 16943 -6359 16989 -6321
rect 16943 -6393 16949 -6359
rect 16983 -6393 16989 -6359
rect 16943 -6699 16989 -6393
rect 17201 -6287 17247 -6240
rect 17201 -6321 17207 -6287
rect 17241 -6321 17247 -6287
rect 17201 -6359 17247 -6321
rect 17201 -6393 17207 -6359
rect 17241 -6393 17247 -6359
rect 16865 -6709 17061 -6699
rect 16865 -6761 16874 -6709
rect 16926 -6761 16938 -6709
rect 16990 -6761 17002 -6709
rect 17054 -6761 17061 -6709
rect 16865 -6769 17061 -6761
rect 16608 -7010 16804 -7000
rect 16608 -7062 16617 -7010
rect 16669 -7062 16681 -7010
rect 16733 -7062 16745 -7010
rect 16797 -7062 16804 -7010
rect 16608 -7070 16804 -7062
rect 16491 -7278 16497 -7244
rect 16531 -7278 16537 -7244
rect 16491 -7316 16537 -7278
rect 16491 -7350 16497 -7316
rect 16531 -7350 16537 -7316
rect 16491 -7397 16537 -7350
rect 16685 -7244 16731 -7070
rect 16685 -7278 16691 -7244
rect 16725 -7278 16731 -7244
rect 16685 -7316 16731 -7278
rect 16685 -7350 16691 -7316
rect 16725 -7350 16731 -7316
rect 16685 -7397 16731 -7350
rect 16943 -7244 16989 -6769
rect 17201 -7000 17247 -6393
rect 17459 -6287 17505 -6240
rect 17459 -6321 17465 -6287
rect 17499 -6321 17505 -6287
rect 17459 -6359 17505 -6321
rect 17459 -6393 17465 -6359
rect 17499 -6393 17505 -6359
rect 17459 -6699 17505 -6393
rect 17717 -6287 17763 -6240
rect 17717 -6321 17723 -6287
rect 17757 -6321 17763 -6287
rect 17717 -6359 17763 -6321
rect 17717 -6393 17723 -6359
rect 17757 -6393 17763 -6359
rect 17383 -6709 17579 -6699
rect 17383 -6761 17392 -6709
rect 17444 -6761 17456 -6709
rect 17508 -6761 17520 -6709
rect 17572 -6761 17579 -6709
rect 17383 -6769 17579 -6761
rect 17126 -7010 17322 -7000
rect 17126 -7062 17135 -7010
rect 17187 -7062 17199 -7010
rect 17251 -7062 17263 -7010
rect 17315 -7062 17322 -7010
rect 17126 -7070 17322 -7062
rect 16943 -7278 16949 -7244
rect 16983 -7278 16989 -7244
rect 16943 -7316 16989 -7278
rect 16943 -7350 16949 -7316
rect 16983 -7350 16989 -7316
rect 16943 -7397 16989 -7350
rect 17201 -7244 17247 -7070
rect 17201 -7278 17207 -7244
rect 17241 -7278 17247 -7244
rect 17201 -7316 17247 -7278
rect 17201 -7350 17207 -7316
rect 17241 -7350 17247 -7316
rect 17201 -7397 17247 -7350
rect 17459 -7244 17505 -6769
rect 17717 -7000 17763 -6393
rect 17911 -6262 18290 -6228
rect 18324 -6262 18347 -6228
rect 17911 -6287 18347 -6262
rect 17911 -6321 17917 -6287
rect 17951 -6321 18175 -6287
rect 18209 -6300 18347 -6287
rect 18209 -6321 18290 -6300
rect 17911 -6334 18290 -6321
rect 18324 -6334 18347 -6300
rect 17911 -6359 18347 -6334
rect 17911 -6393 17917 -6359
rect 17951 -6393 18175 -6359
rect 18209 -6372 18347 -6359
rect 18209 -6393 18290 -6372
rect 17911 -6406 18290 -6393
rect 18324 -6406 18347 -6372
rect 17911 -6444 18347 -6406
rect 17911 -6478 18290 -6444
rect 18324 -6478 18347 -6444
rect 17911 -6516 18347 -6478
rect 17911 -6550 18290 -6516
rect 18324 -6550 18347 -6516
rect 17911 -6588 18347 -6550
rect 17911 -6622 18290 -6588
rect 18324 -6622 18347 -6588
rect 17911 -6660 18347 -6622
rect 17911 -6694 18290 -6660
rect 18324 -6694 18347 -6660
rect 17911 -6732 18347 -6694
rect 17911 -6766 18290 -6732
rect 18324 -6766 18347 -6732
rect 17911 -6804 18347 -6766
rect 17911 -6838 18290 -6804
rect 18324 -6838 18347 -6804
rect 17911 -6876 18347 -6838
rect 17911 -6910 18290 -6876
rect 18324 -6910 18347 -6876
rect 17911 -6948 18347 -6910
rect 17911 -6982 18290 -6948
rect 18324 -6982 18347 -6948
rect 17641 -7010 17837 -7000
rect 17641 -7062 17650 -7010
rect 17702 -7062 17714 -7010
rect 17766 -7062 17778 -7010
rect 17830 -7062 17837 -7010
rect 17641 -7070 17837 -7062
rect 17911 -7020 18347 -6982
rect 17911 -7054 18290 -7020
rect 18324 -7054 18347 -7020
rect 17459 -7278 17465 -7244
rect 17499 -7278 17505 -7244
rect 17459 -7316 17505 -7278
rect 17459 -7350 17465 -7316
rect 17499 -7350 17505 -7316
rect 17459 -7397 17505 -7350
rect 17717 -7244 17763 -7070
rect 17717 -7278 17723 -7244
rect 17757 -7278 17763 -7244
rect 17717 -7316 17763 -7278
rect 17717 -7350 17723 -7316
rect 17757 -7350 17763 -7316
rect 17717 -7397 17763 -7350
rect 17911 -7092 18347 -7054
rect 17911 -7126 18290 -7092
rect 18324 -7126 18347 -7092
rect 17911 -7164 18347 -7126
rect 17911 -7198 18290 -7164
rect 18324 -7198 18347 -7164
rect 17911 -7236 18347 -7198
rect 17911 -7244 18290 -7236
rect 17911 -7278 17917 -7244
rect 17951 -7278 18175 -7244
rect 18209 -7270 18290 -7244
rect 18324 -7270 18347 -7236
rect 18209 -7278 18347 -7270
rect 17911 -7308 18347 -7278
rect 17911 -7316 18290 -7308
rect 17911 -7350 17917 -7316
rect 17951 -7350 18175 -7316
rect 18209 -7342 18290 -7316
rect 18324 -7342 18347 -7308
rect 18209 -7350 18347 -7342
rect 17911 -7380 18347 -7350
rect 9194 -7478 9293 -7444
rect 9327 -7478 9365 -7444
rect 9399 -7452 9781 -7444
rect 9399 -7478 9573 -7452
rect 9194 -7486 9573 -7478
rect 9607 -7478 9781 -7452
rect 9815 -7478 9853 -7444
rect 9887 -7478 9986 -7444
rect 9607 -7486 9986 -7478
rect 9194 -7524 9986 -7486
rect 9194 -7558 9573 -7524
rect 9607 -7558 9986 -7524
rect 9194 -7596 9986 -7558
rect 9194 -7630 9573 -7596
rect 9607 -7630 9986 -7596
rect 9194 -7668 9986 -7630
rect 9194 -7702 9573 -7668
rect 9607 -7702 9986 -7668
rect 9194 -7740 9986 -7702
rect 10190 -7444 11156 -7438
rect 10190 -7478 10233 -7444
rect 10267 -7459 10305 -7444
rect 10339 -7459 10491 -7444
rect 10525 -7459 10563 -7444
rect 10597 -7459 10749 -7444
rect 10783 -7459 10821 -7444
rect 10855 -7459 11007 -7444
rect 11041 -7459 11079 -7444
rect 10190 -7511 10240 -7478
rect 10292 -7511 10304 -7459
rect 10356 -7511 10368 -7459
rect 10420 -7511 10436 -7459
rect 10488 -7478 10491 -7459
rect 10552 -7478 10563 -7459
rect 10488 -7511 10500 -7478
rect 10552 -7511 10564 -7478
rect 10616 -7511 10726 -7459
rect 10783 -7478 10790 -7459
rect 10778 -7511 10790 -7478
rect 10842 -7511 10854 -7478
rect 10906 -7511 10922 -7459
rect 10974 -7511 10986 -7459
rect 11041 -7478 11050 -7459
rect 11113 -7478 11156 -7444
rect 11038 -7511 11050 -7478
rect 11102 -7511 11156 -7478
rect 10190 -7637 11156 -7511
rect 10190 -7689 10240 -7637
rect 10292 -7689 10304 -7637
rect 10356 -7689 10368 -7637
rect 10420 -7689 10436 -7637
rect 10488 -7689 10500 -7637
rect 10552 -7689 10564 -7637
rect 10616 -7689 10726 -7637
rect 10778 -7689 10790 -7637
rect 10842 -7689 10854 -7637
rect 10906 -7689 10922 -7637
rect 10974 -7689 10986 -7637
rect 11038 -7689 11050 -7637
rect 11102 -7689 11156 -7637
rect 10190 -7708 11156 -7689
rect 11233 -7444 12307 -7438
rect 11233 -7478 11459 -7444
rect 11493 -7478 11531 -7444
rect 11565 -7478 11717 -7444
rect 11751 -7478 11789 -7444
rect 11823 -7478 11975 -7444
rect 12009 -7478 12047 -7444
rect 12081 -7478 12307 -7444
rect 11233 -7526 12307 -7478
rect 7886 -7776 8990 -7758
rect 7886 -7806 8078 -7776
rect 8130 -7806 8142 -7776
rect 7886 -7840 8067 -7806
rect 8130 -7828 8139 -7806
rect 8194 -7828 8206 -7776
rect 8258 -7828 8274 -7776
rect 8326 -7806 8338 -7776
rect 8390 -7806 8402 -7776
rect 8390 -7828 8397 -7806
rect 8454 -7828 8564 -7776
rect 8616 -7806 8628 -7776
rect 8680 -7806 8692 -7776
rect 8617 -7828 8628 -7806
rect 8689 -7828 8692 -7806
rect 8744 -7828 8760 -7776
rect 8812 -7828 8824 -7776
rect 8876 -7828 8888 -7776
rect 8940 -7806 8990 -7776
rect 8101 -7840 8139 -7828
rect 8173 -7840 8325 -7828
rect 8359 -7840 8397 -7828
rect 8431 -7840 8583 -7828
rect 8617 -7840 8655 -7828
rect 8689 -7840 8841 -7828
rect 8875 -7840 8913 -7828
rect 8947 -7840 8990 -7806
rect 7886 -7846 8990 -7840
rect 9194 -7774 9573 -7740
rect 9607 -7774 9986 -7740
rect 11233 -7758 11294 -7526
rect 9194 -7806 9986 -7774
rect 9194 -7840 9293 -7806
rect 9327 -7840 9365 -7806
rect 9399 -7812 9781 -7806
rect 9399 -7840 9573 -7812
rect 9194 -7846 9573 -7840
rect 9607 -7840 9781 -7812
rect 9815 -7840 9853 -7806
rect 9887 -7840 9986 -7806
rect 9607 -7846 9986 -7840
rect 10190 -7776 11294 -7758
rect 10190 -7806 10240 -7776
rect 10190 -7840 10233 -7806
rect 10292 -7828 10304 -7776
rect 10356 -7828 10368 -7776
rect 10420 -7828 10436 -7776
rect 10488 -7806 10500 -7776
rect 10552 -7806 10564 -7776
rect 10488 -7828 10491 -7806
rect 10552 -7828 10563 -7806
rect 10616 -7828 10726 -7776
rect 10778 -7806 10790 -7776
rect 10842 -7806 10854 -7776
rect 10783 -7828 10790 -7806
rect 10906 -7828 10922 -7776
rect 10974 -7828 10986 -7776
rect 11038 -7806 11050 -7776
rect 11102 -7806 11294 -7776
rect 11041 -7828 11050 -7806
rect 10267 -7840 10305 -7828
rect 10339 -7840 10491 -7828
rect 10525 -7840 10563 -7828
rect 10597 -7840 10749 -7828
rect 10783 -7840 10821 -7828
rect 10855 -7840 11007 -7828
rect 11041 -7840 11079 -7828
rect 11113 -7840 11294 -7806
rect 10190 -7846 11294 -7840
rect 11416 -7637 12124 -7620
rect 11416 -7689 11450 -7637
rect 11502 -7689 11514 -7637
rect 11566 -7689 11578 -7637
rect 11630 -7689 11646 -7637
rect 11698 -7689 11710 -7637
rect 11762 -7689 11774 -7637
rect 11826 -7689 11838 -7637
rect 11890 -7689 11906 -7637
rect 11958 -7689 11970 -7637
rect 12022 -7689 12034 -7637
rect 12086 -7689 12124 -7637
rect 11416 -7806 12124 -7689
rect 11416 -7840 11459 -7806
rect 11493 -7840 11531 -7806
rect 11565 -7840 11717 -7806
rect 11751 -7840 11789 -7806
rect 11823 -7840 11975 -7806
rect 12009 -7840 12047 -7806
rect 12081 -7840 12124 -7806
rect 11416 -7846 12124 -7840
rect 12246 -7758 12307 -7526
rect 12384 -7444 13350 -7438
rect 12384 -7478 12427 -7444
rect 12461 -7459 12499 -7444
rect 12533 -7459 12685 -7444
rect 12719 -7459 12757 -7444
rect 12791 -7459 12943 -7444
rect 12977 -7459 13015 -7444
rect 13049 -7459 13201 -7444
rect 13235 -7459 13273 -7444
rect 12490 -7478 12499 -7459
rect 12384 -7511 12438 -7478
rect 12490 -7511 12502 -7478
rect 12554 -7511 12566 -7459
rect 12618 -7511 12634 -7459
rect 12750 -7478 12757 -7459
rect 12686 -7511 12698 -7478
rect 12750 -7511 12762 -7478
rect 12814 -7511 12924 -7459
rect 12977 -7478 12988 -7459
rect 13049 -7478 13052 -7459
rect 12976 -7511 12988 -7478
rect 13040 -7511 13052 -7478
rect 13104 -7511 13120 -7459
rect 13172 -7511 13184 -7459
rect 13236 -7511 13248 -7459
rect 13307 -7478 13350 -7444
rect 13300 -7511 13350 -7478
rect 12384 -7637 13350 -7511
rect 12384 -7689 12438 -7637
rect 12490 -7689 12502 -7637
rect 12554 -7689 12566 -7637
rect 12618 -7689 12634 -7637
rect 12686 -7689 12698 -7637
rect 12750 -7689 12762 -7637
rect 12814 -7689 12924 -7637
rect 12976 -7689 12988 -7637
rect 13040 -7689 13052 -7637
rect 13104 -7689 13120 -7637
rect 13172 -7689 13184 -7637
rect 13236 -7689 13248 -7637
rect 13300 -7689 13350 -7637
rect 12384 -7708 13350 -7689
rect 13554 -7444 14344 -7414
rect 17911 -7414 18290 -7380
rect 18324 -7414 18347 -7380
rect 13554 -7478 13653 -7444
rect 13687 -7478 13725 -7444
rect 13759 -7452 14139 -7444
rect 13759 -7478 13932 -7452
rect 13554 -7486 13932 -7478
rect 13966 -7478 14139 -7452
rect 14173 -7478 14211 -7444
rect 14245 -7478 14344 -7444
rect 13966 -7486 14344 -7478
rect 13554 -7524 14344 -7486
rect 13554 -7558 13932 -7524
rect 13966 -7558 14344 -7524
rect 13554 -7596 14344 -7558
rect 13554 -7630 13932 -7596
rect 13966 -7630 14344 -7596
rect 13554 -7668 14344 -7630
rect 13554 -7702 13932 -7668
rect 13966 -7702 14344 -7668
rect 13554 -7740 14344 -7702
rect 14547 -7444 15513 -7438
rect 14547 -7478 14590 -7444
rect 14624 -7459 14662 -7444
rect 14696 -7459 14848 -7444
rect 14882 -7459 14920 -7444
rect 14954 -7459 15106 -7444
rect 15140 -7459 15178 -7444
rect 15212 -7459 15364 -7444
rect 15398 -7459 15436 -7444
rect 14547 -7511 14597 -7478
rect 14649 -7511 14661 -7459
rect 14713 -7511 14725 -7459
rect 14777 -7511 14793 -7459
rect 14845 -7478 14848 -7459
rect 14909 -7478 14920 -7459
rect 14845 -7511 14857 -7478
rect 14909 -7511 14921 -7478
rect 14973 -7511 15083 -7459
rect 15140 -7478 15147 -7459
rect 15135 -7511 15147 -7478
rect 15199 -7511 15211 -7478
rect 15263 -7511 15279 -7459
rect 15331 -7511 15343 -7459
rect 15398 -7478 15407 -7459
rect 15470 -7478 15513 -7444
rect 15395 -7511 15407 -7478
rect 15459 -7511 15513 -7478
rect 14547 -7637 15513 -7511
rect 14547 -7689 14597 -7637
rect 14649 -7689 14661 -7637
rect 14713 -7689 14725 -7637
rect 14777 -7689 14793 -7637
rect 14845 -7689 14857 -7637
rect 14909 -7689 14921 -7637
rect 14973 -7689 15083 -7637
rect 15135 -7689 15147 -7637
rect 15199 -7689 15211 -7637
rect 15263 -7689 15279 -7637
rect 15331 -7689 15343 -7637
rect 15395 -7689 15407 -7637
rect 15459 -7689 15513 -7637
rect 14547 -7708 15513 -7689
rect 15590 -7444 16664 -7438
rect 15590 -7478 15816 -7444
rect 15850 -7478 15888 -7444
rect 15922 -7478 16074 -7444
rect 16108 -7478 16146 -7444
rect 16180 -7478 16332 -7444
rect 16366 -7478 16404 -7444
rect 16438 -7478 16664 -7444
rect 15590 -7526 16664 -7478
rect 12246 -7776 13350 -7758
rect 12246 -7806 12438 -7776
rect 12490 -7806 12502 -7776
rect 12246 -7840 12427 -7806
rect 12490 -7828 12499 -7806
rect 12554 -7828 12566 -7776
rect 12618 -7828 12634 -7776
rect 12686 -7806 12698 -7776
rect 12750 -7806 12762 -7776
rect 12750 -7828 12757 -7806
rect 12814 -7828 12924 -7776
rect 12976 -7806 12988 -7776
rect 13040 -7806 13052 -7776
rect 12977 -7828 12988 -7806
rect 13049 -7828 13052 -7806
rect 13104 -7828 13120 -7776
rect 13172 -7828 13184 -7776
rect 13236 -7828 13248 -7776
rect 13300 -7806 13350 -7776
rect 12461 -7840 12499 -7828
rect 12533 -7840 12685 -7828
rect 12719 -7840 12757 -7828
rect 12791 -7840 12943 -7828
rect 12977 -7840 13015 -7828
rect 13049 -7840 13201 -7828
rect 13235 -7840 13273 -7828
rect 13307 -7840 13350 -7806
rect 12246 -7846 13350 -7840
rect 13554 -7774 13932 -7740
rect 13966 -7774 14344 -7740
rect 15590 -7758 15651 -7526
rect 13554 -7806 14344 -7774
rect 13554 -7840 13653 -7806
rect 13687 -7840 13725 -7806
rect 13759 -7812 14139 -7806
rect 13759 -7840 13932 -7812
rect 13554 -7846 13932 -7840
rect 13966 -7840 14139 -7812
rect 14173 -7840 14211 -7806
rect 14245 -7840 14344 -7806
rect 13966 -7846 14344 -7840
rect 14547 -7776 15651 -7758
rect 14547 -7806 14597 -7776
rect 14547 -7840 14590 -7806
rect 14649 -7828 14661 -7776
rect 14713 -7828 14725 -7776
rect 14777 -7828 14793 -7776
rect 14845 -7806 14857 -7776
rect 14909 -7806 14921 -7776
rect 14845 -7828 14848 -7806
rect 14909 -7828 14920 -7806
rect 14973 -7828 15083 -7776
rect 15135 -7806 15147 -7776
rect 15199 -7806 15211 -7776
rect 15140 -7828 15147 -7806
rect 15263 -7828 15279 -7776
rect 15331 -7828 15343 -7776
rect 15395 -7806 15407 -7776
rect 15459 -7806 15651 -7776
rect 15398 -7828 15407 -7806
rect 14624 -7840 14662 -7828
rect 14696 -7840 14848 -7828
rect 14882 -7840 14920 -7828
rect 14954 -7840 15106 -7828
rect 15140 -7840 15178 -7828
rect 15212 -7840 15364 -7828
rect 15398 -7840 15436 -7828
rect 15470 -7840 15651 -7806
rect 14547 -7846 15651 -7840
rect 15773 -7637 16481 -7620
rect 15773 -7689 15811 -7637
rect 15863 -7689 15875 -7637
rect 15927 -7689 15939 -7637
rect 15991 -7689 16007 -7637
rect 16059 -7689 16071 -7637
rect 16123 -7689 16135 -7637
rect 16187 -7689 16199 -7637
rect 16251 -7689 16267 -7637
rect 16319 -7689 16331 -7637
rect 16383 -7689 16395 -7637
rect 16447 -7689 16481 -7637
rect 15773 -7806 16481 -7689
rect 15773 -7840 15816 -7806
rect 15850 -7840 15888 -7806
rect 15922 -7840 16074 -7806
rect 16108 -7840 16146 -7806
rect 16180 -7840 16332 -7806
rect 16366 -7840 16404 -7806
rect 16438 -7840 16481 -7806
rect 15773 -7846 16481 -7840
rect 16603 -7758 16664 -7526
rect 16741 -7444 17707 -7438
rect 16741 -7478 16784 -7444
rect 16818 -7459 16856 -7444
rect 16890 -7459 17042 -7444
rect 17076 -7459 17114 -7444
rect 17148 -7459 17300 -7444
rect 17334 -7459 17372 -7444
rect 17406 -7459 17558 -7444
rect 17592 -7459 17630 -7444
rect 16847 -7478 16856 -7459
rect 16741 -7511 16795 -7478
rect 16847 -7511 16859 -7478
rect 16911 -7511 16923 -7459
rect 16975 -7511 16991 -7459
rect 17107 -7478 17114 -7459
rect 17043 -7511 17055 -7478
rect 17107 -7511 17119 -7478
rect 17171 -7511 17281 -7459
rect 17334 -7478 17345 -7459
rect 17406 -7478 17409 -7459
rect 17333 -7511 17345 -7478
rect 17397 -7511 17409 -7478
rect 17461 -7511 17477 -7459
rect 17529 -7511 17541 -7459
rect 17593 -7511 17605 -7459
rect 17664 -7478 17707 -7444
rect 17657 -7511 17707 -7478
rect 16741 -7637 17707 -7511
rect 16741 -7689 16795 -7637
rect 16847 -7689 16859 -7637
rect 16911 -7689 16923 -7637
rect 16975 -7689 16991 -7637
rect 17043 -7689 17055 -7637
rect 17107 -7689 17119 -7637
rect 17171 -7689 17281 -7637
rect 17333 -7689 17345 -7637
rect 17397 -7689 17409 -7637
rect 17461 -7689 17477 -7637
rect 17529 -7689 17541 -7637
rect 17593 -7689 17605 -7637
rect 17657 -7689 17707 -7637
rect 16741 -7708 17707 -7689
rect 17911 -7444 18347 -7414
rect 17911 -7478 18010 -7444
rect 18044 -7478 18082 -7444
rect 18116 -7452 18347 -7444
rect 18116 -7478 18290 -7452
rect 17911 -7486 18290 -7478
rect 18324 -7486 18347 -7452
rect 17911 -7524 18347 -7486
rect 17911 -7558 18290 -7524
rect 18324 -7558 18347 -7524
rect 17911 -7596 18347 -7558
rect 17911 -7630 18290 -7596
rect 18324 -7630 18347 -7596
rect 17911 -7668 18347 -7630
rect 17911 -7702 18290 -7668
rect 18324 -7702 18347 -7668
rect 17911 -7740 18347 -7702
rect 16603 -7776 17707 -7758
rect 16603 -7806 16795 -7776
rect 16847 -7806 16859 -7776
rect 16603 -7840 16784 -7806
rect 16847 -7828 16856 -7806
rect 16911 -7828 16923 -7776
rect 16975 -7828 16991 -7776
rect 17043 -7806 17055 -7776
rect 17107 -7806 17119 -7776
rect 17107 -7828 17114 -7806
rect 17171 -7828 17281 -7776
rect 17333 -7806 17345 -7776
rect 17397 -7806 17409 -7776
rect 17334 -7828 17345 -7806
rect 17406 -7828 17409 -7806
rect 17461 -7828 17477 -7776
rect 17529 -7828 17541 -7776
rect 17593 -7828 17605 -7776
rect 17657 -7806 17707 -7776
rect 16818 -7840 16856 -7828
rect 16890 -7840 17042 -7828
rect 17076 -7840 17114 -7828
rect 17148 -7840 17300 -7828
rect 17334 -7840 17372 -7828
rect 17406 -7840 17558 -7828
rect 17592 -7840 17630 -7828
rect 17664 -7840 17707 -7806
rect 16603 -7846 17707 -7840
rect 17911 -7774 18290 -7740
rect 18324 -7774 18347 -7740
rect 17911 -7806 18347 -7774
rect 17911 -7840 18010 -7806
rect 18044 -7840 18082 -7806
rect 18116 -7812 18347 -7806
rect 18116 -7840 18290 -7812
rect 17911 -7846 18290 -7840
rect 18324 -7846 18347 -7812
rect 833 -7884 1269 -7846
rect 833 -7918 856 -7884
rect 890 -7918 1269 -7884
rect 4836 -7884 5626 -7846
rect 833 -7934 1269 -7918
rect 833 -7956 971 -7934
rect 833 -7990 856 -7956
rect 890 -7968 971 -7956
rect 1005 -7968 1229 -7934
rect 1263 -7968 1269 -7934
rect 890 -7990 1269 -7968
rect 833 -8006 1269 -7990
rect 833 -8028 971 -8006
rect 833 -8062 856 -8028
rect 890 -8040 971 -8028
rect 1005 -8040 1229 -8006
rect 1263 -8040 1269 -8006
rect 890 -8062 1269 -8040
rect 833 -8100 1269 -8062
rect 833 -8134 856 -8100
rect 890 -8134 1269 -8100
rect 833 -8172 1269 -8134
rect 833 -8206 856 -8172
rect 890 -8206 1269 -8172
rect 833 -8244 1269 -8206
rect 833 -8278 856 -8244
rect 890 -8278 1269 -8244
rect 833 -8316 1269 -8278
rect 833 -8350 856 -8316
rect 890 -8350 1269 -8316
rect 833 -8388 1269 -8350
rect 833 -8422 856 -8388
rect 890 -8422 1269 -8388
rect 833 -8460 1269 -8422
rect 833 -8494 856 -8460
rect 890 -8494 1269 -8460
rect 833 -8532 1269 -8494
rect 1417 -7934 1463 -7887
rect 1417 -7968 1423 -7934
rect 1457 -7968 1463 -7934
rect 1417 -8006 1463 -7968
rect 1417 -8040 1423 -8006
rect 1457 -8040 1463 -8006
rect 1417 -8521 1463 -8040
rect 1675 -7934 1721 -7887
rect 1675 -7968 1681 -7934
rect 1715 -7968 1721 -7934
rect 1675 -8006 1721 -7968
rect 1675 -8040 1681 -8006
rect 1715 -8040 1721 -8006
rect 1675 -8189 1721 -8040
rect 1933 -7934 1979 -7887
rect 1933 -7968 1939 -7934
rect 1973 -7968 1979 -7934
rect 1933 -8006 1979 -7968
rect 1933 -8040 1939 -8006
rect 1973 -8040 1979 -8006
rect 1598 -8199 1794 -8189
rect 1598 -8251 1607 -8199
rect 1659 -8251 1671 -8199
rect 1723 -8251 1735 -8199
rect 1787 -8251 1794 -8199
rect 1598 -8259 1794 -8251
rect 1933 -8521 1979 -8040
rect 2191 -7934 2237 -7887
rect 2191 -7968 2197 -7934
rect 2231 -7968 2237 -7934
rect 2191 -8006 2237 -7968
rect 2191 -8040 2197 -8006
rect 2231 -8040 2237 -8006
rect 2191 -8189 2237 -8040
rect 2449 -7934 2495 -7887
rect 2449 -7968 2455 -7934
rect 2489 -7968 2495 -7934
rect 2449 -8006 2495 -7968
rect 2449 -8040 2455 -8006
rect 2489 -8040 2495 -8006
rect 2116 -8199 2312 -8189
rect 2116 -8251 2125 -8199
rect 2177 -8251 2189 -8199
rect 2241 -8251 2253 -8199
rect 2305 -8251 2312 -8199
rect 2116 -8259 2312 -8251
rect 2449 -8521 2495 -8040
rect 2643 -7934 2689 -7887
rect 2643 -7968 2649 -7934
rect 2683 -7968 2689 -7934
rect 2643 -8006 2689 -7968
rect 2643 -8040 2649 -8006
rect 2683 -8040 2689 -8006
rect 2643 -8358 2689 -8040
rect 2901 -7934 2947 -7887
rect 2901 -7968 2907 -7934
rect 2941 -7968 2947 -7934
rect 2901 -8006 2947 -7968
rect 2901 -8040 2907 -8006
rect 2941 -8040 2947 -8006
rect 2570 -8368 2766 -8358
rect 2570 -8420 2577 -8368
rect 2629 -8420 2641 -8368
rect 2693 -8420 2705 -8368
rect 2757 -8420 2766 -8368
rect 2570 -8428 2766 -8420
rect 833 -8566 856 -8532
rect 890 -8566 1269 -8532
rect 833 -8604 1269 -8566
rect 1339 -8531 1535 -8521
rect 1339 -8583 1348 -8531
rect 1400 -8583 1412 -8531
rect 1464 -8583 1476 -8531
rect 1528 -8583 1535 -8531
rect 1339 -8591 1535 -8583
rect 1856 -8531 2052 -8521
rect 1856 -8583 1865 -8531
rect 1917 -8583 1929 -8531
rect 1981 -8583 1993 -8531
rect 2045 -8583 2052 -8531
rect 1856 -8591 2052 -8583
rect 2373 -8531 2569 -8521
rect 2373 -8583 2382 -8531
rect 2434 -8583 2446 -8531
rect 2498 -8583 2510 -8531
rect 2562 -8583 2569 -8531
rect 2373 -8591 2569 -8583
rect 833 -8638 856 -8604
rect 890 -8638 1269 -8604
rect 833 -8676 1269 -8638
rect 833 -8710 856 -8676
rect 890 -8710 1269 -8676
rect 2901 -8689 2947 -8040
rect 3159 -7934 3205 -7887
rect 3159 -7968 3165 -7934
rect 3199 -7968 3205 -7934
rect 3159 -8006 3205 -7968
rect 3159 -8040 3165 -8006
rect 3199 -8040 3205 -8006
rect 3159 -8358 3205 -8040
rect 3417 -7934 3463 -7887
rect 3417 -7968 3423 -7934
rect 3457 -7968 3463 -7934
rect 3417 -8006 3463 -7968
rect 3417 -8040 3423 -8006
rect 3457 -8040 3463 -8006
rect 3087 -8368 3283 -8358
rect 3087 -8420 3094 -8368
rect 3146 -8420 3158 -8368
rect 3210 -8420 3222 -8368
rect 3274 -8420 3283 -8368
rect 3087 -8428 3283 -8420
rect 3417 -8689 3463 -8040
rect 3611 -7934 3657 -7887
rect 3611 -7968 3617 -7934
rect 3651 -7968 3657 -7934
rect 3611 -8006 3657 -7968
rect 3611 -8040 3617 -8006
rect 3651 -8040 3657 -8006
rect 3611 -8521 3657 -8040
rect 3869 -7934 3915 -7887
rect 3869 -7968 3875 -7934
rect 3909 -7968 3915 -7934
rect 3869 -8006 3915 -7968
rect 3869 -8040 3875 -8006
rect 3909 -8040 3915 -8006
rect 3869 -8189 3915 -8040
rect 4127 -7934 4173 -7887
rect 4127 -7968 4133 -7934
rect 4167 -7968 4173 -7934
rect 4127 -8006 4173 -7968
rect 4127 -8040 4133 -8006
rect 4167 -8040 4173 -8006
rect 3793 -8199 3989 -8189
rect 3793 -8251 3802 -8199
rect 3854 -8251 3866 -8199
rect 3918 -8251 3930 -8199
rect 3982 -8251 3989 -8199
rect 3793 -8259 3989 -8251
rect 4127 -8521 4173 -8040
rect 4385 -7934 4431 -7887
rect 4385 -7968 4391 -7934
rect 4425 -7968 4431 -7934
rect 4385 -8006 4431 -7968
rect 4385 -8040 4391 -8006
rect 4425 -8040 4431 -8006
rect 4385 -8189 4431 -8040
rect 4643 -7934 4689 -7887
rect 4643 -7968 4649 -7934
rect 4683 -7968 4689 -7934
rect 4643 -8006 4689 -7968
rect 4643 -8040 4649 -8006
rect 4683 -8040 4689 -8006
rect 4310 -8199 4506 -8189
rect 4310 -8251 4319 -8199
rect 4371 -8251 4383 -8199
rect 4435 -8251 4447 -8199
rect 4499 -8251 4506 -8199
rect 4310 -8259 4506 -8251
rect 4643 -8521 4689 -8040
rect 4836 -7918 5214 -7884
rect 5248 -7918 5626 -7884
rect 9194 -7884 9986 -7846
rect 4836 -7934 5626 -7918
rect 4836 -7968 4842 -7934
rect 4876 -7968 5100 -7934
rect 5134 -7956 5328 -7934
rect 5134 -7968 5214 -7956
rect 4836 -7990 5214 -7968
rect 5248 -7968 5328 -7956
rect 5362 -7968 5586 -7934
rect 5620 -7968 5626 -7934
rect 5248 -7990 5626 -7968
rect 4836 -8006 5626 -7990
rect 4836 -8040 4842 -8006
rect 4876 -8040 5100 -8006
rect 5134 -8028 5328 -8006
rect 5134 -8040 5214 -8028
rect 4836 -8062 5214 -8040
rect 5248 -8040 5328 -8028
rect 5362 -8040 5586 -8006
rect 5620 -8040 5626 -8006
rect 5248 -8062 5626 -8040
rect 4836 -8100 5626 -8062
rect 4836 -8134 5214 -8100
rect 5248 -8134 5626 -8100
rect 4836 -8172 5626 -8134
rect 4836 -8206 5214 -8172
rect 5248 -8206 5626 -8172
rect 4836 -8244 5626 -8206
rect 4836 -8278 5214 -8244
rect 5248 -8278 5626 -8244
rect 4836 -8316 5626 -8278
rect 4836 -8350 5214 -8316
rect 5248 -8350 5626 -8316
rect 4836 -8388 5626 -8350
rect 4836 -8422 5214 -8388
rect 5248 -8422 5626 -8388
rect 4836 -8460 5626 -8422
rect 4836 -8494 5214 -8460
rect 5248 -8494 5626 -8460
rect 3534 -8531 3730 -8521
rect 3534 -8583 3543 -8531
rect 3595 -8583 3607 -8531
rect 3659 -8583 3671 -8531
rect 3723 -8583 3730 -8531
rect 3534 -8591 3730 -8583
rect 4051 -8531 4247 -8521
rect 4051 -8583 4060 -8531
rect 4112 -8583 4124 -8531
rect 4176 -8583 4188 -8531
rect 4240 -8583 4247 -8531
rect 4051 -8591 4247 -8583
rect 4566 -8531 4762 -8521
rect 4566 -8583 4575 -8531
rect 4627 -8583 4639 -8531
rect 4691 -8583 4703 -8531
rect 4755 -8583 4762 -8531
rect 4566 -8591 4762 -8583
rect 4836 -8532 5626 -8494
rect 5774 -7934 5820 -7887
rect 5774 -7968 5780 -7934
rect 5814 -7968 5820 -7934
rect 5774 -8006 5820 -7968
rect 5774 -8040 5780 -8006
rect 5814 -8040 5820 -8006
rect 5774 -8521 5820 -8040
rect 6032 -7934 6078 -7887
rect 6032 -7968 6038 -7934
rect 6072 -7968 6078 -7934
rect 6032 -8006 6078 -7968
rect 6032 -8040 6038 -8006
rect 6072 -8040 6078 -8006
rect 6032 -8189 6078 -8040
rect 6290 -7934 6336 -7887
rect 6290 -7968 6296 -7934
rect 6330 -7968 6336 -7934
rect 6290 -8006 6336 -7968
rect 6290 -8040 6296 -8006
rect 6330 -8040 6336 -8006
rect 5957 -8199 6153 -8189
rect 5957 -8251 5964 -8199
rect 6016 -8251 6028 -8199
rect 6080 -8251 6092 -8199
rect 6144 -8251 6153 -8199
rect 5957 -8259 6153 -8251
rect 6290 -8521 6336 -8040
rect 6548 -7934 6594 -7887
rect 6548 -7968 6554 -7934
rect 6588 -7968 6594 -7934
rect 6548 -8006 6594 -7968
rect 6548 -8040 6554 -8006
rect 6588 -8040 6594 -8006
rect 6548 -8189 6594 -8040
rect 6806 -7934 6852 -7887
rect 6806 -7968 6812 -7934
rect 6846 -7968 6852 -7934
rect 6806 -8006 6852 -7968
rect 6806 -8040 6812 -8006
rect 6846 -8040 6852 -8006
rect 6474 -8199 6670 -8189
rect 6474 -8251 6481 -8199
rect 6533 -8251 6545 -8199
rect 6597 -8251 6609 -8199
rect 6661 -8251 6670 -8199
rect 6474 -8259 6670 -8251
rect 6806 -8521 6852 -8040
rect 7000 -7934 7046 -7887
rect 7000 -7968 7006 -7934
rect 7040 -7968 7046 -7934
rect 7000 -8006 7046 -7968
rect 7000 -8040 7006 -8006
rect 7040 -8040 7046 -8006
rect 4836 -8566 5214 -8532
rect 5248 -8566 5626 -8532
rect 4836 -8604 5626 -8566
rect 5701 -8531 5897 -8521
rect 5701 -8583 5708 -8531
rect 5760 -8583 5772 -8531
rect 5824 -8583 5836 -8531
rect 5888 -8583 5897 -8531
rect 5701 -8591 5897 -8583
rect 6216 -8531 6412 -8521
rect 6216 -8583 6223 -8531
rect 6275 -8583 6287 -8531
rect 6339 -8583 6351 -8531
rect 6403 -8583 6412 -8531
rect 6216 -8591 6412 -8583
rect 6733 -8531 6929 -8521
rect 6733 -8583 6740 -8531
rect 6792 -8583 6804 -8531
rect 6856 -8583 6868 -8531
rect 6920 -8583 6929 -8531
rect 6733 -8591 6929 -8583
rect 4836 -8638 5214 -8604
rect 5248 -8638 5626 -8604
rect 4836 -8676 5626 -8638
rect 833 -8748 1269 -8710
rect 833 -8782 856 -8748
rect 890 -8782 1269 -8748
rect 2827 -8699 3023 -8689
rect 2827 -8751 2834 -8699
rect 2886 -8751 2898 -8699
rect 2950 -8751 2962 -8699
rect 3014 -8751 3023 -8699
rect 2827 -8759 3023 -8751
rect 3344 -8699 3540 -8689
rect 3344 -8751 3351 -8699
rect 3403 -8751 3415 -8699
rect 3467 -8751 3479 -8699
rect 3531 -8751 3540 -8699
rect 3344 -8759 3540 -8751
rect 4836 -8710 5214 -8676
rect 5248 -8710 5626 -8676
rect 7000 -8689 7046 -8040
rect 7258 -7934 7304 -7887
rect 7258 -7968 7264 -7934
rect 7298 -7968 7304 -7934
rect 7258 -8006 7304 -7968
rect 7258 -8040 7264 -8006
rect 7298 -8040 7304 -8006
rect 7258 -8358 7304 -8040
rect 7516 -7934 7562 -7887
rect 7516 -7968 7522 -7934
rect 7556 -7968 7562 -7934
rect 7516 -8006 7562 -7968
rect 7516 -8040 7522 -8006
rect 7556 -8040 7562 -8006
rect 7180 -8368 7376 -8358
rect 7180 -8420 7189 -8368
rect 7241 -8420 7253 -8368
rect 7305 -8420 7317 -8368
rect 7369 -8420 7376 -8368
rect 7180 -8428 7376 -8420
rect 7516 -8689 7562 -8040
rect 7774 -7934 7820 -7887
rect 7774 -7968 7780 -7934
rect 7814 -7968 7820 -7934
rect 7774 -8006 7820 -7968
rect 7774 -8040 7780 -8006
rect 7814 -8040 7820 -8006
rect 7774 -8358 7820 -8040
rect 7968 -7934 8014 -7887
rect 7968 -7968 7974 -7934
rect 8008 -7968 8014 -7934
rect 7968 -8006 8014 -7968
rect 7968 -8040 7974 -8006
rect 8008 -8040 8014 -8006
rect 7697 -8368 7893 -8358
rect 7697 -8420 7706 -8368
rect 7758 -8420 7770 -8368
rect 7822 -8420 7834 -8368
rect 7886 -8420 7893 -8368
rect 7697 -8428 7893 -8420
rect 7968 -8521 8014 -8040
rect 8226 -7934 8272 -7887
rect 8226 -7968 8232 -7934
rect 8266 -7968 8272 -7934
rect 8226 -8006 8272 -7968
rect 8226 -8040 8232 -8006
rect 8266 -8040 8272 -8006
rect 8226 -8189 8272 -8040
rect 8484 -7934 8530 -7887
rect 8484 -7968 8490 -7934
rect 8524 -7968 8530 -7934
rect 8484 -8006 8530 -7968
rect 8484 -8040 8490 -8006
rect 8524 -8040 8530 -8006
rect 8151 -8199 8347 -8189
rect 8151 -8251 8158 -8199
rect 8210 -8251 8222 -8199
rect 8274 -8251 8286 -8199
rect 8338 -8251 8347 -8199
rect 8151 -8259 8347 -8251
rect 8484 -8521 8530 -8040
rect 8742 -7934 8788 -7887
rect 8742 -7968 8748 -7934
rect 8782 -7968 8788 -7934
rect 8742 -8006 8788 -7968
rect 8742 -8040 8748 -8006
rect 8782 -8040 8788 -8006
rect 8742 -8189 8788 -8040
rect 9000 -7934 9046 -7887
rect 9000 -7968 9006 -7934
rect 9040 -7968 9046 -7934
rect 9000 -8006 9046 -7968
rect 9000 -8040 9006 -8006
rect 9040 -8040 9046 -8006
rect 8668 -8199 8864 -8189
rect 8668 -8251 8675 -8199
rect 8727 -8251 8739 -8199
rect 8791 -8251 8803 -8199
rect 8855 -8251 8864 -8199
rect 8668 -8259 8864 -8251
rect 9000 -8521 9046 -8040
rect 9194 -7918 9573 -7884
rect 9607 -7918 9986 -7884
rect 13554 -7884 14344 -7846
rect 9194 -7934 9986 -7918
rect 9194 -7968 9200 -7934
rect 9234 -7968 9458 -7934
rect 9492 -7956 9688 -7934
rect 9492 -7968 9573 -7956
rect 9194 -7990 9573 -7968
rect 9607 -7968 9688 -7956
rect 9722 -7968 9946 -7934
rect 9980 -7968 9986 -7934
rect 9607 -7990 9986 -7968
rect 9194 -8006 9986 -7990
rect 9194 -8040 9200 -8006
rect 9234 -8040 9458 -8006
rect 9492 -8028 9688 -8006
rect 9492 -8040 9573 -8028
rect 9194 -8062 9573 -8040
rect 9607 -8040 9688 -8028
rect 9722 -8040 9946 -8006
rect 9980 -8040 9986 -8006
rect 9607 -8062 9986 -8040
rect 9194 -8100 9986 -8062
rect 9194 -8134 9573 -8100
rect 9607 -8134 9986 -8100
rect 9194 -8172 9986 -8134
rect 9194 -8206 9573 -8172
rect 9607 -8206 9986 -8172
rect 9194 -8244 9986 -8206
rect 9194 -8278 9573 -8244
rect 9607 -8278 9986 -8244
rect 9194 -8316 9986 -8278
rect 9194 -8350 9573 -8316
rect 9607 -8350 9986 -8316
rect 9194 -8388 9986 -8350
rect 9194 -8422 9573 -8388
rect 9607 -8422 9986 -8388
rect 9194 -8460 9986 -8422
rect 9194 -8494 9573 -8460
rect 9607 -8494 9986 -8460
rect 7894 -8531 8090 -8521
rect 7894 -8583 7901 -8531
rect 7953 -8583 7965 -8531
rect 8017 -8583 8029 -8531
rect 8081 -8583 8090 -8531
rect 7894 -8591 8090 -8583
rect 8410 -8531 8606 -8521
rect 8410 -8583 8417 -8531
rect 8469 -8583 8481 -8531
rect 8533 -8583 8545 -8531
rect 8597 -8583 8606 -8531
rect 8410 -8591 8606 -8583
rect 8928 -8531 9124 -8521
rect 8928 -8583 8935 -8531
rect 8987 -8583 8999 -8531
rect 9051 -8583 9063 -8531
rect 9115 -8583 9124 -8531
rect 8928 -8591 9124 -8583
rect 9194 -8532 9986 -8494
rect 10134 -7934 10180 -7887
rect 10134 -7968 10140 -7934
rect 10174 -7968 10180 -7934
rect 10134 -8006 10180 -7968
rect 10134 -8040 10140 -8006
rect 10174 -8040 10180 -8006
rect 10134 -8521 10180 -8040
rect 10392 -7934 10438 -7887
rect 10392 -7968 10398 -7934
rect 10432 -7968 10438 -7934
rect 10392 -8006 10438 -7968
rect 10392 -8040 10398 -8006
rect 10432 -8040 10438 -8006
rect 10392 -8189 10438 -8040
rect 10650 -7934 10696 -7887
rect 10650 -7968 10656 -7934
rect 10690 -7968 10696 -7934
rect 10650 -8006 10696 -7968
rect 10650 -8040 10656 -8006
rect 10690 -8040 10696 -8006
rect 10316 -8199 10512 -8189
rect 10316 -8251 10325 -8199
rect 10377 -8251 10389 -8199
rect 10441 -8251 10453 -8199
rect 10505 -8251 10512 -8199
rect 10316 -8259 10512 -8251
rect 10650 -8521 10696 -8040
rect 10908 -7934 10954 -7887
rect 10908 -7968 10914 -7934
rect 10948 -7968 10954 -7934
rect 10908 -8006 10954 -7968
rect 10908 -8040 10914 -8006
rect 10948 -8040 10954 -8006
rect 10908 -8189 10954 -8040
rect 11166 -7934 11212 -7887
rect 11166 -7968 11172 -7934
rect 11206 -7968 11212 -7934
rect 11166 -8006 11212 -7968
rect 11166 -8040 11172 -8006
rect 11206 -8040 11212 -8006
rect 10833 -8199 11029 -8189
rect 10833 -8251 10842 -8199
rect 10894 -8251 10906 -8199
rect 10958 -8251 10970 -8199
rect 11022 -8251 11029 -8199
rect 10833 -8259 11029 -8251
rect 11166 -8521 11212 -8040
rect 11360 -7934 11406 -7887
rect 11360 -7968 11366 -7934
rect 11400 -7968 11406 -7934
rect 11360 -8006 11406 -7968
rect 11360 -8040 11366 -8006
rect 11400 -8040 11406 -8006
rect 11360 -8358 11406 -8040
rect 11618 -7934 11664 -7887
rect 11618 -7968 11624 -7934
rect 11658 -7968 11664 -7934
rect 11618 -8006 11664 -7968
rect 11618 -8040 11624 -8006
rect 11658 -8040 11664 -8006
rect 11287 -8368 11483 -8358
rect 11287 -8420 11294 -8368
rect 11346 -8420 11358 -8368
rect 11410 -8420 11422 -8368
rect 11474 -8420 11483 -8368
rect 11287 -8428 11483 -8420
rect 9194 -8566 9573 -8532
rect 9607 -8566 9986 -8532
rect 9194 -8604 9986 -8566
rect 10056 -8531 10252 -8521
rect 10056 -8583 10065 -8531
rect 10117 -8583 10129 -8531
rect 10181 -8583 10193 -8531
rect 10245 -8583 10252 -8531
rect 10056 -8591 10252 -8583
rect 10574 -8531 10770 -8521
rect 10574 -8583 10583 -8531
rect 10635 -8583 10647 -8531
rect 10699 -8583 10711 -8531
rect 10763 -8583 10770 -8531
rect 10574 -8591 10770 -8583
rect 11090 -8531 11286 -8521
rect 11090 -8583 11099 -8531
rect 11151 -8583 11163 -8531
rect 11215 -8583 11227 -8531
rect 11279 -8583 11286 -8531
rect 11090 -8591 11286 -8583
rect 9194 -8638 9573 -8604
rect 9607 -8638 9986 -8604
rect 9194 -8676 9986 -8638
rect 4836 -8748 5626 -8710
rect 833 -8820 1269 -8782
rect 833 -8854 856 -8820
rect 890 -8854 1269 -8820
rect 4836 -8782 5214 -8748
rect 5248 -8782 5626 -8748
rect 6922 -8699 7118 -8689
rect 6922 -8751 6931 -8699
rect 6983 -8751 6995 -8699
rect 7047 -8751 7059 -8699
rect 7111 -8751 7118 -8699
rect 6922 -8759 7118 -8751
rect 7440 -8699 7636 -8689
rect 7440 -8751 7449 -8699
rect 7501 -8751 7513 -8699
rect 7565 -8751 7577 -8699
rect 7629 -8751 7636 -8699
rect 7440 -8759 7636 -8751
rect 9194 -8710 9573 -8676
rect 9607 -8710 9986 -8676
rect 11618 -8689 11664 -8040
rect 11876 -7934 11922 -7887
rect 11876 -7968 11882 -7934
rect 11916 -7968 11922 -7934
rect 11876 -8006 11922 -7968
rect 11876 -8040 11882 -8006
rect 11916 -8040 11922 -8006
rect 11876 -8358 11922 -8040
rect 12134 -7934 12180 -7887
rect 12134 -7968 12140 -7934
rect 12174 -7968 12180 -7934
rect 12134 -8006 12180 -7968
rect 12134 -8040 12140 -8006
rect 12174 -8040 12180 -8006
rect 11804 -8368 12000 -8358
rect 11804 -8420 11811 -8368
rect 11863 -8420 11875 -8368
rect 11927 -8420 11939 -8368
rect 11991 -8420 12000 -8368
rect 11804 -8428 12000 -8420
rect 12134 -8689 12180 -8040
rect 12328 -7934 12374 -7887
rect 12328 -7968 12334 -7934
rect 12368 -7968 12374 -7934
rect 12328 -8006 12374 -7968
rect 12328 -8040 12334 -8006
rect 12368 -8040 12374 -8006
rect 12328 -8521 12374 -8040
rect 12586 -7934 12632 -7887
rect 12586 -7968 12592 -7934
rect 12626 -7968 12632 -7934
rect 12586 -8006 12632 -7968
rect 12586 -8040 12592 -8006
rect 12626 -8040 12632 -8006
rect 12586 -8189 12632 -8040
rect 12844 -7934 12890 -7887
rect 12844 -7968 12850 -7934
rect 12884 -7968 12890 -7934
rect 12844 -8006 12890 -7968
rect 12844 -8040 12850 -8006
rect 12884 -8040 12890 -8006
rect 12510 -8199 12706 -8189
rect 12510 -8251 12519 -8199
rect 12571 -8251 12583 -8199
rect 12635 -8251 12647 -8199
rect 12699 -8251 12706 -8199
rect 12510 -8259 12706 -8251
rect 12844 -8521 12890 -8040
rect 13102 -7934 13148 -7887
rect 13102 -7968 13108 -7934
rect 13142 -7968 13148 -7934
rect 13102 -8006 13148 -7968
rect 13102 -8040 13108 -8006
rect 13142 -8040 13148 -8006
rect 13102 -8189 13148 -8040
rect 13360 -7934 13406 -7887
rect 13360 -7968 13366 -7934
rect 13400 -7968 13406 -7934
rect 13360 -8006 13406 -7968
rect 13360 -8040 13366 -8006
rect 13400 -8040 13406 -8006
rect 13027 -8199 13223 -8189
rect 13027 -8251 13036 -8199
rect 13088 -8251 13100 -8199
rect 13152 -8251 13164 -8199
rect 13216 -8251 13223 -8199
rect 13027 -8259 13223 -8251
rect 13360 -8521 13406 -8040
rect 13554 -7918 13932 -7884
rect 13966 -7918 14344 -7884
rect 17911 -7884 18347 -7846
rect 13554 -7934 14344 -7918
rect 13554 -7968 13560 -7934
rect 13594 -7968 13818 -7934
rect 13852 -7956 14046 -7934
rect 13852 -7968 13932 -7956
rect 13554 -7990 13932 -7968
rect 13966 -7968 14046 -7956
rect 14080 -7968 14304 -7934
rect 14338 -7968 14344 -7934
rect 13966 -7990 14344 -7968
rect 13554 -8006 14344 -7990
rect 13554 -8040 13560 -8006
rect 13594 -8040 13818 -8006
rect 13852 -8028 14046 -8006
rect 13852 -8040 13932 -8028
rect 13554 -8062 13932 -8040
rect 13966 -8040 14046 -8028
rect 14080 -8040 14304 -8006
rect 14338 -8040 14344 -8006
rect 13966 -8062 14344 -8040
rect 13554 -8100 14344 -8062
rect 13554 -8134 13932 -8100
rect 13966 -8134 14344 -8100
rect 13554 -8172 14344 -8134
rect 13554 -8206 13932 -8172
rect 13966 -8206 14344 -8172
rect 13554 -8244 14344 -8206
rect 13554 -8278 13932 -8244
rect 13966 -8278 14344 -8244
rect 13554 -8316 14344 -8278
rect 13554 -8350 13932 -8316
rect 13966 -8350 14344 -8316
rect 13554 -8388 14344 -8350
rect 13554 -8422 13932 -8388
rect 13966 -8422 14344 -8388
rect 13554 -8460 14344 -8422
rect 13554 -8494 13932 -8460
rect 13966 -8494 14344 -8460
rect 12251 -8531 12447 -8521
rect 12251 -8583 12260 -8531
rect 12312 -8583 12324 -8531
rect 12376 -8583 12388 -8531
rect 12440 -8583 12447 -8531
rect 12251 -8591 12447 -8583
rect 12768 -8531 12964 -8521
rect 12768 -8583 12777 -8531
rect 12829 -8583 12841 -8531
rect 12893 -8583 12905 -8531
rect 12957 -8583 12964 -8531
rect 12768 -8591 12964 -8583
rect 13283 -8531 13479 -8521
rect 13283 -8583 13292 -8531
rect 13344 -8583 13356 -8531
rect 13408 -8583 13420 -8531
rect 13472 -8583 13479 -8531
rect 13283 -8591 13479 -8583
rect 13554 -8532 14344 -8494
rect 14491 -7934 14537 -7887
rect 14491 -7968 14497 -7934
rect 14531 -7968 14537 -7934
rect 14491 -8006 14537 -7968
rect 14491 -8040 14497 -8006
rect 14531 -8040 14537 -8006
rect 14491 -8521 14537 -8040
rect 14749 -7934 14795 -7887
rect 14749 -7968 14755 -7934
rect 14789 -7968 14795 -7934
rect 14749 -8006 14795 -7968
rect 14749 -8040 14755 -8006
rect 14789 -8040 14795 -8006
rect 14749 -8189 14795 -8040
rect 15007 -7934 15053 -7887
rect 15007 -7968 15013 -7934
rect 15047 -7968 15053 -7934
rect 15007 -8006 15053 -7968
rect 15007 -8040 15013 -8006
rect 15047 -8040 15053 -8006
rect 14674 -8199 14870 -8189
rect 14674 -8251 14681 -8199
rect 14733 -8251 14745 -8199
rect 14797 -8251 14809 -8199
rect 14861 -8251 14870 -8199
rect 14674 -8259 14870 -8251
rect 15007 -8521 15053 -8040
rect 15265 -7934 15311 -7887
rect 15265 -7968 15271 -7934
rect 15305 -7968 15311 -7934
rect 15265 -8006 15311 -7968
rect 15265 -8040 15271 -8006
rect 15305 -8040 15311 -8006
rect 15265 -8189 15311 -8040
rect 15523 -7934 15569 -7887
rect 15523 -7968 15529 -7934
rect 15563 -7968 15569 -7934
rect 15523 -8006 15569 -7968
rect 15523 -8040 15529 -8006
rect 15563 -8040 15569 -8006
rect 15191 -8199 15387 -8189
rect 15191 -8251 15198 -8199
rect 15250 -8251 15262 -8199
rect 15314 -8251 15326 -8199
rect 15378 -8251 15387 -8199
rect 15191 -8259 15387 -8251
rect 15523 -8521 15569 -8040
rect 15717 -7934 15763 -7887
rect 15717 -7968 15723 -7934
rect 15757 -7968 15763 -7934
rect 15717 -8006 15763 -7968
rect 15717 -8040 15723 -8006
rect 15757 -8040 15763 -8006
rect 13554 -8566 13932 -8532
rect 13966 -8566 14344 -8532
rect 13554 -8604 14344 -8566
rect 14418 -8531 14614 -8521
rect 14418 -8583 14425 -8531
rect 14477 -8583 14489 -8531
rect 14541 -8583 14553 -8531
rect 14605 -8583 14614 -8531
rect 14418 -8591 14614 -8583
rect 14933 -8531 15129 -8521
rect 14933 -8583 14940 -8531
rect 14992 -8583 15004 -8531
rect 15056 -8583 15068 -8531
rect 15120 -8583 15129 -8531
rect 14933 -8591 15129 -8583
rect 15450 -8531 15646 -8521
rect 15450 -8583 15457 -8531
rect 15509 -8583 15521 -8531
rect 15573 -8583 15585 -8531
rect 15637 -8583 15646 -8531
rect 15450 -8591 15646 -8583
rect 13554 -8638 13932 -8604
rect 13966 -8638 14344 -8604
rect 13554 -8676 14344 -8638
rect 9194 -8748 9986 -8710
rect 4836 -8820 5626 -8782
rect 833 -8878 1269 -8854
rect 833 -8892 971 -8878
rect 833 -8926 856 -8892
rect 890 -8912 971 -8892
rect 1005 -8912 1229 -8878
rect 1263 -8912 1269 -8878
rect 890 -8926 1269 -8912
rect 833 -8950 1269 -8926
rect 833 -8964 971 -8950
rect 833 -8998 856 -8964
rect 890 -8984 971 -8964
rect 1005 -8984 1229 -8950
rect 1263 -8984 1269 -8950
rect 890 -8998 1269 -8984
rect 833 -9036 1269 -8998
rect 833 -9070 856 -9036
rect 890 -9070 1269 -9036
rect 833 -9072 1269 -9070
rect 1417 -8878 1463 -8831
rect 1417 -8912 1423 -8878
rect 1457 -8912 1463 -8878
rect 1417 -8950 1463 -8912
rect 1417 -8984 1423 -8950
rect 1457 -8984 1463 -8950
rect 1417 -9072 1463 -8984
rect 1675 -8878 1721 -8831
rect 1675 -8912 1681 -8878
rect 1715 -8912 1721 -8878
rect 1675 -8950 1721 -8912
rect 1675 -8984 1681 -8950
rect 1715 -8984 1721 -8950
rect 1675 -9072 1721 -8984
rect 1933 -8878 1979 -8831
rect 1933 -8912 1939 -8878
rect 1973 -8912 1979 -8878
rect 1933 -8950 1979 -8912
rect 1933 -8984 1939 -8950
rect 1973 -8984 1979 -8950
rect 1933 -9072 1979 -8984
rect 2191 -8878 2237 -8831
rect 2191 -8912 2197 -8878
rect 2231 -8912 2237 -8878
rect 2191 -8950 2237 -8912
rect 2191 -8984 2197 -8950
rect 2231 -8984 2237 -8950
rect 2191 -9072 2237 -8984
rect 2449 -8878 2495 -8831
rect 2449 -8912 2455 -8878
rect 2489 -8912 2495 -8878
rect 2449 -8950 2495 -8912
rect 2449 -8984 2455 -8950
rect 2489 -8984 2495 -8950
rect 2449 -9072 2495 -8984
rect 2643 -8878 2689 -8831
rect 2643 -8912 2649 -8878
rect 2683 -8912 2689 -8878
rect 2643 -8950 2689 -8912
rect 2643 -8984 2649 -8950
rect 2683 -8984 2689 -8950
rect 2643 -9072 2689 -8984
rect 2901 -8878 2947 -8831
rect 2901 -8912 2907 -8878
rect 2941 -8912 2947 -8878
rect 2901 -8950 2947 -8912
rect 2901 -8984 2907 -8950
rect 2941 -8984 2947 -8950
rect 2901 -9072 2947 -8984
rect 3159 -8878 3205 -8831
rect 3159 -8912 3165 -8878
rect 3199 -8912 3205 -8878
rect 3159 -8950 3205 -8912
rect 3159 -8984 3165 -8950
rect 3199 -8984 3205 -8950
rect 3159 -9072 3205 -8984
rect 3417 -8878 3463 -8831
rect 3417 -8912 3423 -8878
rect 3457 -8912 3463 -8878
rect 3417 -8950 3463 -8912
rect 3417 -8984 3423 -8950
rect 3457 -8984 3463 -8950
rect 3417 -9072 3463 -8984
rect 3611 -8878 3657 -8831
rect 3611 -8912 3617 -8878
rect 3651 -8912 3657 -8878
rect 3611 -8950 3657 -8912
rect 3611 -8984 3617 -8950
rect 3651 -8984 3657 -8950
rect 3611 -9072 3657 -8984
rect 3869 -8878 3915 -8831
rect 3869 -8912 3875 -8878
rect 3909 -8912 3915 -8878
rect 3869 -8950 3915 -8912
rect 3869 -8984 3875 -8950
rect 3909 -8984 3915 -8950
rect 3869 -9072 3915 -8984
rect 4127 -8878 4173 -8831
rect 4127 -8912 4133 -8878
rect 4167 -8912 4173 -8878
rect 4127 -8950 4173 -8912
rect 4127 -8984 4133 -8950
rect 4167 -8984 4173 -8950
rect 4127 -9072 4173 -8984
rect 4385 -8878 4431 -8831
rect 4385 -8912 4391 -8878
rect 4425 -8912 4431 -8878
rect 4385 -8950 4431 -8912
rect 4385 -8984 4391 -8950
rect 4425 -8984 4431 -8950
rect 4385 -9072 4431 -8984
rect 4643 -8878 4689 -8831
rect 4643 -8912 4649 -8878
rect 4683 -8912 4689 -8878
rect 4643 -8950 4689 -8912
rect 4643 -8984 4649 -8950
rect 4683 -8984 4689 -8950
rect 4643 -9072 4689 -8984
rect 4836 -8854 5214 -8820
rect 5248 -8854 5626 -8820
rect 9194 -8782 9573 -8748
rect 9607 -8782 9986 -8748
rect 11544 -8699 11740 -8689
rect 11544 -8751 11551 -8699
rect 11603 -8751 11615 -8699
rect 11667 -8751 11679 -8699
rect 11731 -8751 11740 -8699
rect 11544 -8759 11740 -8751
rect 12062 -8699 12258 -8689
rect 12062 -8751 12069 -8699
rect 12121 -8751 12133 -8699
rect 12185 -8751 12197 -8699
rect 12249 -8751 12258 -8699
rect 12062 -8759 12258 -8751
rect 13554 -8710 13932 -8676
rect 13966 -8710 14344 -8676
rect 15717 -8689 15763 -8040
rect 15975 -7934 16021 -7887
rect 15975 -7968 15981 -7934
rect 16015 -7968 16021 -7934
rect 15975 -8006 16021 -7968
rect 15975 -8040 15981 -8006
rect 16015 -8040 16021 -8006
rect 15975 -8358 16021 -8040
rect 16233 -7934 16279 -7887
rect 16233 -7968 16239 -7934
rect 16273 -7968 16279 -7934
rect 16233 -8006 16279 -7968
rect 16233 -8040 16239 -8006
rect 16273 -8040 16279 -8006
rect 15897 -8368 16093 -8358
rect 15897 -8420 15906 -8368
rect 15958 -8420 15970 -8368
rect 16022 -8420 16034 -8368
rect 16086 -8420 16093 -8368
rect 15897 -8428 16093 -8420
rect 16233 -8689 16279 -8040
rect 16491 -7934 16537 -7887
rect 16491 -7968 16497 -7934
rect 16531 -7968 16537 -7934
rect 16491 -8006 16537 -7968
rect 16491 -8040 16497 -8006
rect 16531 -8040 16537 -8006
rect 16491 -8358 16537 -8040
rect 16685 -7934 16731 -7887
rect 16685 -7968 16691 -7934
rect 16725 -7968 16731 -7934
rect 16685 -8006 16731 -7968
rect 16685 -8040 16691 -8006
rect 16725 -8040 16731 -8006
rect 16414 -8368 16610 -8358
rect 16414 -8420 16423 -8368
rect 16475 -8420 16487 -8368
rect 16539 -8420 16551 -8368
rect 16603 -8420 16610 -8368
rect 16414 -8428 16610 -8420
rect 16685 -8521 16731 -8040
rect 16943 -7934 16989 -7887
rect 16943 -7968 16949 -7934
rect 16983 -7968 16989 -7934
rect 16943 -8006 16989 -7968
rect 16943 -8040 16949 -8006
rect 16983 -8040 16989 -8006
rect 16943 -8189 16989 -8040
rect 17201 -7934 17247 -7887
rect 17201 -7968 17207 -7934
rect 17241 -7968 17247 -7934
rect 17201 -8006 17247 -7968
rect 17201 -8040 17207 -8006
rect 17241 -8040 17247 -8006
rect 16868 -8199 17064 -8189
rect 16868 -8251 16875 -8199
rect 16927 -8251 16939 -8199
rect 16991 -8251 17003 -8199
rect 17055 -8251 17064 -8199
rect 16868 -8259 17064 -8251
rect 17201 -8521 17247 -8040
rect 17459 -7934 17505 -7887
rect 17459 -7968 17465 -7934
rect 17499 -7968 17505 -7934
rect 17459 -8006 17505 -7968
rect 17459 -8040 17465 -8006
rect 17499 -8040 17505 -8006
rect 17459 -8189 17505 -8040
rect 17717 -7934 17763 -7887
rect 17717 -7968 17723 -7934
rect 17757 -7968 17763 -7934
rect 17717 -8006 17763 -7968
rect 17717 -8040 17723 -8006
rect 17757 -8040 17763 -8006
rect 17386 -8199 17582 -8189
rect 17386 -8251 17393 -8199
rect 17445 -8251 17457 -8199
rect 17509 -8251 17521 -8199
rect 17573 -8251 17582 -8199
rect 17386 -8259 17582 -8251
rect 17717 -8521 17763 -8040
rect 17911 -7918 18290 -7884
rect 18324 -7918 18347 -7884
rect 17911 -7934 18347 -7918
rect 17911 -7968 17917 -7934
rect 17951 -7968 18175 -7934
rect 18209 -7956 18347 -7934
rect 18209 -7968 18290 -7956
rect 17911 -7990 18290 -7968
rect 18324 -7990 18347 -7956
rect 17911 -8006 18347 -7990
rect 17911 -8040 17917 -8006
rect 17951 -8040 18175 -8006
rect 18209 -8028 18347 -8006
rect 18209 -8040 18290 -8028
rect 17911 -8062 18290 -8040
rect 18324 -8062 18347 -8028
rect 17911 -8100 18347 -8062
rect 17911 -8134 18290 -8100
rect 18324 -8134 18347 -8100
rect 17911 -8172 18347 -8134
rect 17911 -8206 18290 -8172
rect 18324 -8206 18347 -8172
rect 17911 -8244 18347 -8206
rect 17911 -8278 18290 -8244
rect 18324 -8278 18347 -8244
rect 17911 -8316 18347 -8278
rect 17911 -8350 18290 -8316
rect 18324 -8350 18347 -8316
rect 17911 -8388 18347 -8350
rect 17911 -8422 18290 -8388
rect 18324 -8422 18347 -8388
rect 17911 -8460 18347 -8422
rect 17911 -8494 18290 -8460
rect 18324 -8494 18347 -8460
rect 16611 -8531 16807 -8521
rect 16611 -8583 16618 -8531
rect 16670 -8583 16682 -8531
rect 16734 -8583 16746 -8531
rect 16798 -8583 16807 -8531
rect 16611 -8591 16807 -8583
rect 17128 -8531 17324 -8521
rect 17128 -8583 17135 -8531
rect 17187 -8583 17199 -8531
rect 17251 -8583 17263 -8531
rect 17315 -8583 17324 -8531
rect 17128 -8591 17324 -8583
rect 17645 -8531 17841 -8521
rect 17645 -8583 17652 -8531
rect 17704 -8583 17716 -8531
rect 17768 -8583 17780 -8531
rect 17832 -8583 17841 -8531
rect 17645 -8591 17841 -8583
rect 17911 -8532 18347 -8494
rect 17911 -8566 18290 -8532
rect 18324 -8566 18347 -8532
rect 17911 -8604 18347 -8566
rect 17911 -8638 18290 -8604
rect 18324 -8638 18347 -8604
rect 17911 -8676 18347 -8638
rect 13554 -8748 14344 -8710
rect 9194 -8820 9986 -8782
rect 4836 -8878 5626 -8854
rect 4836 -8912 4842 -8878
rect 4876 -8912 5100 -8878
rect 5134 -8892 5328 -8878
rect 5134 -8912 5214 -8892
rect 4836 -8926 5214 -8912
rect 5248 -8912 5328 -8892
rect 5362 -8912 5586 -8878
rect 5620 -8912 5626 -8878
rect 5248 -8926 5626 -8912
rect 4836 -8950 5626 -8926
rect 4836 -8984 4842 -8950
rect 4876 -8984 5100 -8950
rect 5134 -8964 5328 -8950
rect 5134 -8984 5214 -8964
rect 4836 -8998 5214 -8984
rect 5248 -8984 5328 -8964
rect 5362 -8984 5586 -8950
rect 5620 -8984 5626 -8950
rect 5248 -8998 5626 -8984
rect 4836 -9036 5626 -8998
rect 4836 -9070 5214 -9036
rect 5248 -9070 5626 -9036
rect 4836 -9072 5626 -9070
rect 5774 -8878 5820 -8831
rect 5774 -8912 5780 -8878
rect 5814 -8912 5820 -8878
rect 5774 -8950 5820 -8912
rect 5774 -8984 5780 -8950
rect 5814 -8984 5820 -8950
rect 5774 -9072 5820 -8984
rect 6032 -8878 6078 -8831
rect 6032 -8912 6038 -8878
rect 6072 -8912 6078 -8878
rect 6032 -8950 6078 -8912
rect 6032 -8984 6038 -8950
rect 6072 -8984 6078 -8950
rect 6032 -9072 6078 -8984
rect 6290 -8878 6336 -8831
rect 6290 -8912 6296 -8878
rect 6330 -8912 6336 -8878
rect 6290 -8950 6336 -8912
rect 6290 -8984 6296 -8950
rect 6330 -8984 6336 -8950
rect 6290 -9072 6336 -8984
rect 6548 -8878 6594 -8831
rect 6548 -8912 6554 -8878
rect 6588 -8912 6594 -8878
rect 6548 -8950 6594 -8912
rect 6548 -8984 6554 -8950
rect 6588 -8984 6594 -8950
rect 6548 -9072 6594 -8984
rect 6806 -8878 6852 -8831
rect 6806 -8912 6812 -8878
rect 6846 -8912 6852 -8878
rect 6806 -8950 6852 -8912
rect 6806 -8984 6812 -8950
rect 6846 -8984 6852 -8950
rect 6806 -9072 6852 -8984
rect 7000 -8878 7046 -8831
rect 7000 -8912 7006 -8878
rect 7040 -8912 7046 -8878
rect 7000 -8950 7046 -8912
rect 7000 -8984 7006 -8950
rect 7040 -8984 7046 -8950
rect 7000 -9072 7046 -8984
rect 7258 -8878 7304 -8831
rect 7258 -8912 7264 -8878
rect 7298 -8912 7304 -8878
rect 7258 -8950 7304 -8912
rect 7258 -8984 7264 -8950
rect 7298 -8984 7304 -8950
rect 7258 -9072 7304 -8984
rect 7516 -8878 7562 -8831
rect 7516 -8912 7522 -8878
rect 7556 -8912 7562 -8878
rect 7516 -8950 7562 -8912
rect 7516 -8984 7522 -8950
rect 7556 -8984 7562 -8950
rect 7516 -9072 7562 -8984
rect 7774 -8878 7820 -8831
rect 7774 -8912 7780 -8878
rect 7814 -8912 7820 -8878
rect 7774 -8950 7820 -8912
rect 7774 -8984 7780 -8950
rect 7814 -8984 7820 -8950
rect 7774 -9072 7820 -8984
rect 7968 -8878 8014 -8831
rect 7968 -8912 7974 -8878
rect 8008 -8912 8014 -8878
rect 7968 -8950 8014 -8912
rect 7968 -8984 7974 -8950
rect 8008 -8984 8014 -8950
rect 7968 -9072 8014 -8984
rect 8226 -8878 8272 -8831
rect 8226 -8912 8232 -8878
rect 8266 -8912 8272 -8878
rect 8226 -8950 8272 -8912
rect 8226 -8984 8232 -8950
rect 8266 -8984 8272 -8950
rect 8226 -9072 8272 -8984
rect 8484 -8878 8530 -8831
rect 8484 -8912 8490 -8878
rect 8524 -8912 8530 -8878
rect 8484 -8950 8530 -8912
rect 8484 -8984 8490 -8950
rect 8524 -8984 8530 -8950
rect 8484 -9072 8530 -8984
rect 8742 -8878 8788 -8831
rect 8742 -8912 8748 -8878
rect 8782 -8912 8788 -8878
rect 8742 -8950 8788 -8912
rect 8742 -8984 8748 -8950
rect 8782 -8984 8788 -8950
rect 8742 -9072 8788 -8984
rect 9000 -8878 9046 -8831
rect 9000 -8912 9006 -8878
rect 9040 -8912 9046 -8878
rect 9000 -8950 9046 -8912
rect 9000 -8984 9006 -8950
rect 9040 -8984 9046 -8950
rect 9000 -9072 9046 -8984
rect 9194 -8854 9573 -8820
rect 9607 -8854 9986 -8820
rect 13554 -8782 13932 -8748
rect 13966 -8782 14344 -8748
rect 15640 -8699 15836 -8689
rect 15640 -8751 15649 -8699
rect 15701 -8751 15713 -8699
rect 15765 -8751 15777 -8699
rect 15829 -8751 15836 -8699
rect 15640 -8759 15836 -8751
rect 16157 -8699 16353 -8689
rect 16157 -8751 16166 -8699
rect 16218 -8751 16230 -8699
rect 16282 -8751 16294 -8699
rect 16346 -8751 16353 -8699
rect 16157 -8759 16353 -8751
rect 17911 -8710 18290 -8676
rect 18324 -8710 18347 -8676
rect 17911 -8748 18347 -8710
rect 13554 -8820 14344 -8782
rect 9194 -8878 9986 -8854
rect 9194 -8912 9200 -8878
rect 9234 -8912 9458 -8878
rect 9492 -8892 9688 -8878
rect 9492 -8912 9573 -8892
rect 9194 -8926 9573 -8912
rect 9607 -8912 9688 -8892
rect 9722 -8912 9946 -8878
rect 9980 -8912 9986 -8878
rect 9607 -8926 9986 -8912
rect 9194 -8950 9986 -8926
rect 9194 -8984 9200 -8950
rect 9234 -8984 9458 -8950
rect 9492 -8964 9688 -8950
rect 9492 -8984 9573 -8964
rect 9194 -8998 9573 -8984
rect 9607 -8984 9688 -8964
rect 9722 -8984 9946 -8950
rect 9980 -8984 9986 -8950
rect 9607 -8998 9986 -8984
rect 9194 -9036 9986 -8998
rect 9194 -9070 9573 -9036
rect 9607 -9070 9986 -9036
rect 9194 -9072 9986 -9070
rect 10134 -8878 10180 -8831
rect 10134 -8912 10140 -8878
rect 10174 -8912 10180 -8878
rect 10134 -8950 10180 -8912
rect 10134 -8984 10140 -8950
rect 10174 -8984 10180 -8950
rect 10134 -9072 10180 -8984
rect 10392 -8878 10438 -8831
rect 10392 -8912 10398 -8878
rect 10432 -8912 10438 -8878
rect 10392 -8950 10438 -8912
rect 10392 -8984 10398 -8950
rect 10432 -8984 10438 -8950
rect 10392 -9072 10438 -8984
rect 10650 -8878 10696 -8831
rect 10650 -8912 10656 -8878
rect 10690 -8912 10696 -8878
rect 10650 -8950 10696 -8912
rect 10650 -8984 10656 -8950
rect 10690 -8984 10696 -8950
rect 10650 -9072 10696 -8984
rect 10908 -8878 10954 -8831
rect 10908 -8912 10914 -8878
rect 10948 -8912 10954 -8878
rect 10908 -8950 10954 -8912
rect 10908 -8984 10914 -8950
rect 10948 -8984 10954 -8950
rect 10908 -9072 10954 -8984
rect 11166 -8878 11212 -8831
rect 11166 -8912 11172 -8878
rect 11206 -8912 11212 -8878
rect 11166 -8950 11212 -8912
rect 11166 -8984 11172 -8950
rect 11206 -8984 11212 -8950
rect 11166 -9072 11212 -8984
rect 11360 -8878 11406 -8831
rect 11360 -8912 11366 -8878
rect 11400 -8912 11406 -8878
rect 11360 -8950 11406 -8912
rect 11360 -8984 11366 -8950
rect 11400 -8984 11406 -8950
rect 11360 -9072 11406 -8984
rect 11618 -8878 11664 -8831
rect 11618 -8912 11624 -8878
rect 11658 -8912 11664 -8878
rect 11618 -8950 11664 -8912
rect 11618 -8984 11624 -8950
rect 11658 -8984 11664 -8950
rect 11618 -9072 11664 -8984
rect 11876 -8878 11922 -8831
rect 11876 -8912 11882 -8878
rect 11916 -8912 11922 -8878
rect 11876 -8950 11922 -8912
rect 11876 -8984 11882 -8950
rect 11916 -8984 11922 -8950
rect 11876 -9072 11922 -8984
rect 12134 -8878 12180 -8831
rect 12134 -8912 12140 -8878
rect 12174 -8912 12180 -8878
rect 12134 -8950 12180 -8912
rect 12134 -8984 12140 -8950
rect 12174 -8984 12180 -8950
rect 12134 -9072 12180 -8984
rect 12328 -8878 12374 -8831
rect 12328 -8912 12334 -8878
rect 12368 -8912 12374 -8878
rect 12328 -8950 12374 -8912
rect 12328 -8984 12334 -8950
rect 12368 -8984 12374 -8950
rect 12328 -9072 12374 -8984
rect 12586 -8878 12632 -8831
rect 12586 -8912 12592 -8878
rect 12626 -8912 12632 -8878
rect 12586 -8950 12632 -8912
rect 12586 -8984 12592 -8950
rect 12626 -8984 12632 -8950
rect 12586 -9072 12632 -8984
rect 12844 -8878 12890 -8831
rect 12844 -8912 12850 -8878
rect 12884 -8912 12890 -8878
rect 12844 -8950 12890 -8912
rect 12844 -8984 12850 -8950
rect 12884 -8984 12890 -8950
rect 12844 -9072 12890 -8984
rect 13102 -8878 13148 -8831
rect 13102 -8912 13108 -8878
rect 13142 -8912 13148 -8878
rect 13102 -8950 13148 -8912
rect 13102 -8984 13108 -8950
rect 13142 -8984 13148 -8950
rect 13102 -9072 13148 -8984
rect 13360 -8878 13406 -8831
rect 13360 -8912 13366 -8878
rect 13400 -8912 13406 -8878
rect 13360 -8950 13406 -8912
rect 13360 -8984 13366 -8950
rect 13400 -8984 13406 -8950
rect 13360 -9072 13406 -8984
rect 13554 -8854 13932 -8820
rect 13966 -8854 14344 -8820
rect 17911 -8782 18290 -8748
rect 18324 -8782 18347 -8748
rect 17911 -8820 18347 -8782
rect 13554 -8878 14344 -8854
rect 13554 -8912 13560 -8878
rect 13594 -8912 13818 -8878
rect 13852 -8892 14046 -8878
rect 13852 -8912 13932 -8892
rect 13554 -8926 13932 -8912
rect 13966 -8912 14046 -8892
rect 14080 -8912 14304 -8878
rect 14338 -8912 14344 -8878
rect 13966 -8926 14344 -8912
rect 13554 -8950 14344 -8926
rect 13554 -8984 13560 -8950
rect 13594 -8984 13818 -8950
rect 13852 -8964 14046 -8950
rect 13852 -8984 13932 -8964
rect 13554 -8998 13932 -8984
rect 13966 -8984 14046 -8964
rect 14080 -8984 14304 -8950
rect 14338 -8984 14344 -8950
rect 13966 -8998 14344 -8984
rect 13554 -9036 14344 -8998
rect 13554 -9070 13932 -9036
rect 13966 -9070 14344 -9036
rect 13554 -9072 14344 -9070
rect 14491 -8878 14537 -8831
rect 14491 -8912 14497 -8878
rect 14531 -8912 14537 -8878
rect 14491 -8950 14537 -8912
rect 14491 -8984 14497 -8950
rect 14531 -8984 14537 -8950
rect 14491 -9072 14537 -8984
rect 14749 -8878 14795 -8831
rect 14749 -8912 14755 -8878
rect 14789 -8912 14795 -8878
rect 14749 -8950 14795 -8912
rect 14749 -8984 14755 -8950
rect 14789 -8984 14795 -8950
rect 14749 -9072 14795 -8984
rect 15007 -8878 15053 -8831
rect 15007 -8912 15013 -8878
rect 15047 -8912 15053 -8878
rect 15007 -8950 15053 -8912
rect 15007 -8984 15013 -8950
rect 15047 -8984 15053 -8950
rect 15007 -9072 15053 -8984
rect 15265 -8878 15311 -8831
rect 15265 -8912 15271 -8878
rect 15305 -8912 15311 -8878
rect 15265 -8950 15311 -8912
rect 15265 -8984 15271 -8950
rect 15305 -8984 15311 -8950
rect 15265 -9072 15311 -8984
rect 15523 -8878 15569 -8831
rect 15523 -8912 15529 -8878
rect 15563 -8912 15569 -8878
rect 15523 -8950 15569 -8912
rect 15523 -8984 15529 -8950
rect 15563 -8984 15569 -8950
rect 15523 -9072 15569 -8984
rect 15717 -8878 15763 -8831
rect 15717 -8912 15723 -8878
rect 15757 -8912 15763 -8878
rect 15717 -8950 15763 -8912
rect 15717 -8984 15723 -8950
rect 15757 -8984 15763 -8950
rect 15717 -9072 15763 -8984
rect 15975 -8878 16021 -8831
rect 15975 -8912 15981 -8878
rect 16015 -8912 16021 -8878
rect 15975 -8950 16021 -8912
rect 15975 -8984 15981 -8950
rect 16015 -8984 16021 -8950
rect 15975 -9072 16021 -8984
rect 16233 -8878 16279 -8831
rect 16233 -8912 16239 -8878
rect 16273 -8912 16279 -8878
rect 16233 -8950 16279 -8912
rect 16233 -8984 16239 -8950
rect 16273 -8984 16279 -8950
rect 16233 -9072 16279 -8984
rect 16491 -8878 16537 -8831
rect 16491 -8912 16497 -8878
rect 16531 -8912 16537 -8878
rect 16491 -8950 16537 -8912
rect 16491 -8984 16497 -8950
rect 16531 -8984 16537 -8950
rect 16491 -9072 16537 -8984
rect 16685 -8878 16731 -8831
rect 16685 -8912 16691 -8878
rect 16725 -8912 16731 -8878
rect 16685 -8950 16731 -8912
rect 16685 -8984 16691 -8950
rect 16725 -8984 16731 -8950
rect 16685 -9072 16731 -8984
rect 16943 -8878 16989 -8831
rect 16943 -8912 16949 -8878
rect 16983 -8912 16989 -8878
rect 16943 -8950 16989 -8912
rect 16943 -8984 16949 -8950
rect 16983 -8984 16989 -8950
rect 16943 -9072 16989 -8984
rect 17201 -8878 17247 -8831
rect 17201 -8912 17207 -8878
rect 17241 -8912 17247 -8878
rect 17201 -8950 17247 -8912
rect 17201 -8984 17207 -8950
rect 17241 -8984 17247 -8950
rect 17201 -9072 17247 -8984
rect 17459 -8878 17505 -8831
rect 17459 -8912 17465 -8878
rect 17499 -8912 17505 -8878
rect 17459 -8950 17505 -8912
rect 17459 -8984 17465 -8950
rect 17499 -8984 17505 -8950
rect 17459 -9072 17505 -8984
rect 17717 -8878 17763 -8831
rect 17717 -8912 17723 -8878
rect 17757 -8912 17763 -8878
rect 17717 -8950 17763 -8912
rect 17717 -8984 17723 -8950
rect 17757 -8984 17763 -8950
rect 17717 -9072 17763 -8984
rect 17911 -8854 18290 -8820
rect 18324 -8854 18347 -8820
rect 17911 -8878 18347 -8854
rect 17911 -8912 17917 -8878
rect 17951 -8912 18175 -8878
rect 18209 -8892 18347 -8878
rect 18209 -8912 18290 -8892
rect 17911 -8926 18290 -8912
rect 18324 -8926 18347 -8892
rect 17911 -8950 18347 -8926
rect 17911 -8984 17917 -8950
rect 17951 -8984 18175 -8950
rect 18209 -8964 18347 -8950
rect 18209 -8984 18290 -8964
rect 17911 -8998 18290 -8984
rect 18324 -8998 18347 -8964
rect 17911 -9036 18347 -8998
rect 17911 -9070 18290 -9036
rect 18324 -9070 18347 -9036
rect 17911 -9072 18347 -9070
rect 831 -9078 18349 -9072
rect 831 -9112 1064 -9078
rect 1098 -9112 1136 -9078
rect 1170 -9112 1516 -9078
rect 1550 -9112 1588 -9078
rect 1622 -9112 1774 -9078
rect 1808 -9112 1846 -9078
rect 1880 -9112 2032 -9078
rect 2066 -9112 2104 -9078
rect 2138 -9112 2290 -9078
rect 2324 -9112 2362 -9078
rect 2396 -9112 2742 -9078
rect 2776 -9112 2814 -9078
rect 2848 -9112 3000 -9078
rect 3034 -9112 3072 -9078
rect 3106 -9112 3258 -9078
rect 3292 -9112 3330 -9078
rect 3364 -9112 3710 -9078
rect 3744 -9112 3782 -9078
rect 3816 -9112 3968 -9078
rect 4002 -9112 4040 -9078
rect 4074 -9112 4226 -9078
rect 4260 -9112 4298 -9078
rect 4332 -9112 4484 -9078
rect 4518 -9112 4556 -9078
rect 4590 -9112 4935 -9078
rect 4969 -9112 5007 -9078
rect 5041 -9112 5421 -9078
rect 5455 -9112 5493 -9078
rect 5527 -9112 5873 -9078
rect 5907 -9112 5945 -9078
rect 5979 -9112 6131 -9078
rect 6165 -9112 6203 -9078
rect 6237 -9112 6389 -9078
rect 6423 -9112 6461 -9078
rect 6495 -9112 6647 -9078
rect 6681 -9112 6719 -9078
rect 6753 -9112 7099 -9078
rect 7133 -9112 7171 -9078
rect 7205 -9112 7357 -9078
rect 7391 -9112 7429 -9078
rect 7463 -9112 7615 -9078
rect 7649 -9112 7687 -9078
rect 7721 -9112 8067 -9078
rect 8101 -9112 8139 -9078
rect 8173 -9112 8325 -9078
rect 8359 -9112 8397 -9078
rect 8431 -9112 8583 -9078
rect 8617 -9112 8655 -9078
rect 8689 -9112 8841 -9078
rect 8875 -9112 8913 -9078
rect 8947 -9112 9293 -9078
rect 9327 -9112 9365 -9078
rect 9399 -9112 9781 -9078
rect 9815 -9112 9853 -9078
rect 9887 -9112 10233 -9078
rect 10267 -9112 10305 -9078
rect 10339 -9112 10491 -9078
rect 10525 -9112 10563 -9078
rect 10597 -9112 10749 -9078
rect 10783 -9112 10821 -9078
rect 10855 -9112 11007 -9078
rect 11041 -9112 11079 -9078
rect 11113 -9112 11459 -9078
rect 11493 -9112 11531 -9078
rect 11565 -9112 11717 -9078
rect 11751 -9112 11789 -9078
rect 11823 -9112 11975 -9078
rect 12009 -9112 12047 -9078
rect 12081 -9112 12427 -9078
rect 12461 -9112 12499 -9078
rect 12533 -9112 12685 -9078
rect 12719 -9112 12757 -9078
rect 12791 -9112 12943 -9078
rect 12977 -9112 13015 -9078
rect 13049 -9112 13201 -9078
rect 13235 -9112 13273 -9078
rect 13307 -9112 13653 -9078
rect 13687 -9112 13725 -9078
rect 13759 -9112 14139 -9078
rect 14173 -9112 14211 -9078
rect 14245 -9112 14590 -9078
rect 14624 -9112 14662 -9078
rect 14696 -9112 14848 -9078
rect 14882 -9112 14920 -9078
rect 14954 -9112 15106 -9078
rect 15140 -9112 15178 -9078
rect 15212 -9112 15364 -9078
rect 15398 -9112 15436 -9078
rect 15470 -9112 15816 -9078
rect 15850 -9112 15888 -9078
rect 15922 -9112 16074 -9078
rect 16108 -9112 16146 -9078
rect 16180 -9112 16332 -9078
rect 16366 -9112 16404 -9078
rect 16438 -9112 16784 -9078
rect 16818 -9112 16856 -9078
rect 16890 -9112 17042 -9078
rect 17076 -9112 17114 -9078
rect 17148 -9112 17300 -9078
rect 17334 -9112 17372 -9078
rect 17406 -9112 17558 -9078
rect 17592 -9112 17630 -9078
rect 17664 -9112 18010 -9078
rect 18044 -9112 18082 -9078
rect 18116 -9112 18349 -9078
rect 831 -9192 18349 -9112
rect 831 -9226 930 -9192
rect 964 -9226 1002 -9192
rect 1036 -9226 1074 -9192
rect 1108 -9226 1146 -9192
rect 1180 -9226 1218 -9192
rect 1252 -9226 1290 -9192
rect 1324 -9226 1362 -9192
rect 1396 -9226 1434 -9192
rect 1468 -9226 1506 -9192
rect 1540 -9226 1578 -9192
rect 1612 -9226 1650 -9192
rect 1684 -9226 1722 -9192
rect 1756 -9226 1794 -9192
rect 1828 -9226 1866 -9192
rect 1900 -9226 1938 -9192
rect 1972 -9226 2010 -9192
rect 2044 -9226 2082 -9192
rect 2116 -9226 2154 -9192
rect 2188 -9226 2226 -9192
rect 2260 -9226 2298 -9192
rect 2332 -9226 2370 -9192
rect 2404 -9226 2442 -9192
rect 2476 -9226 2514 -9192
rect 2548 -9226 2586 -9192
rect 2620 -9226 2658 -9192
rect 2692 -9226 2730 -9192
rect 2764 -9226 2802 -9192
rect 2836 -9226 2874 -9192
rect 2908 -9226 2946 -9192
rect 2980 -9226 3018 -9192
rect 3052 -9226 3090 -9192
rect 3124 -9226 3162 -9192
rect 3196 -9226 3234 -9192
rect 3268 -9226 3306 -9192
rect 3340 -9226 3378 -9192
rect 3412 -9226 3450 -9192
rect 3484 -9226 3522 -9192
rect 3556 -9226 3594 -9192
rect 3628 -9226 3666 -9192
rect 3700 -9226 3738 -9192
rect 3772 -9226 3810 -9192
rect 3844 -9226 3882 -9192
rect 3916 -9226 3954 -9192
rect 3988 -9226 4026 -9192
rect 4060 -9226 4098 -9192
rect 4132 -9226 4170 -9192
rect 4204 -9226 4242 -9192
rect 4276 -9226 4314 -9192
rect 4348 -9226 4386 -9192
rect 4420 -9226 4458 -9192
rect 4492 -9226 4530 -9192
rect 4564 -9226 4602 -9192
rect 4636 -9226 4674 -9192
rect 4708 -9226 4746 -9192
rect 4780 -9226 4818 -9192
rect 4852 -9226 4890 -9192
rect 4924 -9226 4962 -9192
rect 4996 -9226 5034 -9192
rect 5068 -9226 5106 -9192
rect 5140 -9226 5323 -9192
rect 5357 -9226 5395 -9192
rect 5429 -9226 5467 -9192
rect 5501 -9226 5539 -9192
rect 5573 -9226 5611 -9192
rect 5645 -9226 5683 -9192
rect 5717 -9226 5755 -9192
rect 5789 -9226 5827 -9192
rect 5861 -9226 5899 -9192
rect 5933 -9226 5971 -9192
rect 6005 -9226 6043 -9192
rect 6077 -9226 6115 -9192
rect 6149 -9226 6187 -9192
rect 6221 -9226 6259 -9192
rect 6293 -9226 6331 -9192
rect 6365 -9226 6403 -9192
rect 6437 -9226 6475 -9192
rect 6509 -9226 6547 -9192
rect 6581 -9226 6619 -9192
rect 6653 -9226 6691 -9192
rect 6725 -9226 6763 -9192
rect 6797 -9226 6835 -9192
rect 6869 -9226 6907 -9192
rect 6941 -9226 6979 -9192
rect 7013 -9226 7051 -9192
rect 7085 -9226 7123 -9192
rect 7157 -9226 7195 -9192
rect 7229 -9226 7267 -9192
rect 7301 -9226 7339 -9192
rect 7373 -9226 7411 -9192
rect 7445 -9226 7483 -9192
rect 7517 -9226 7555 -9192
rect 7589 -9226 7627 -9192
rect 7661 -9226 7699 -9192
rect 7733 -9226 7771 -9192
rect 7805 -9226 7843 -9192
rect 7877 -9226 7915 -9192
rect 7949 -9226 7987 -9192
rect 8021 -9226 8059 -9192
rect 8093 -9226 8131 -9192
rect 8165 -9226 8203 -9192
rect 8237 -9226 8275 -9192
rect 8309 -9226 8347 -9192
rect 8381 -9226 8419 -9192
rect 8453 -9226 8491 -9192
rect 8525 -9226 8563 -9192
rect 8597 -9226 8635 -9192
rect 8669 -9226 8707 -9192
rect 8741 -9226 8779 -9192
rect 8813 -9226 8851 -9192
rect 8885 -9226 8923 -9192
rect 8957 -9226 8995 -9192
rect 9029 -9226 9067 -9192
rect 9101 -9226 9139 -9192
rect 9173 -9226 9211 -9192
rect 9245 -9226 9283 -9192
rect 9317 -9226 9355 -9192
rect 9389 -9226 9427 -9192
rect 9461 -9226 9499 -9192
rect 9533 -9226 9647 -9192
rect 9681 -9226 9719 -9192
rect 9753 -9226 9791 -9192
rect 9825 -9226 9863 -9192
rect 9897 -9226 9935 -9192
rect 9969 -9226 10007 -9192
rect 10041 -9226 10079 -9192
rect 10113 -9226 10151 -9192
rect 10185 -9226 10223 -9192
rect 10257 -9226 10295 -9192
rect 10329 -9226 10367 -9192
rect 10401 -9226 10439 -9192
rect 10473 -9226 10511 -9192
rect 10545 -9226 10583 -9192
rect 10617 -9226 10655 -9192
rect 10689 -9226 10727 -9192
rect 10761 -9226 10799 -9192
rect 10833 -9226 10871 -9192
rect 10905 -9226 10943 -9192
rect 10977 -9226 11015 -9192
rect 11049 -9226 11087 -9192
rect 11121 -9226 11159 -9192
rect 11193 -9226 11231 -9192
rect 11265 -9226 11303 -9192
rect 11337 -9226 11375 -9192
rect 11409 -9226 11447 -9192
rect 11481 -9226 11519 -9192
rect 11553 -9226 11591 -9192
rect 11625 -9226 11663 -9192
rect 11697 -9226 11735 -9192
rect 11769 -9226 11807 -9192
rect 11841 -9226 11879 -9192
rect 11913 -9226 11951 -9192
rect 11985 -9226 12023 -9192
rect 12057 -9226 12095 -9192
rect 12129 -9226 12167 -9192
rect 12201 -9226 12239 -9192
rect 12273 -9226 12311 -9192
rect 12345 -9226 12383 -9192
rect 12417 -9226 12455 -9192
rect 12489 -9226 12527 -9192
rect 12561 -9226 12599 -9192
rect 12633 -9226 12671 -9192
rect 12705 -9226 12743 -9192
rect 12777 -9226 12815 -9192
rect 12849 -9226 12887 -9192
rect 12921 -9226 12959 -9192
rect 12993 -9226 13031 -9192
rect 13065 -9226 13103 -9192
rect 13137 -9226 13175 -9192
rect 13209 -9226 13247 -9192
rect 13281 -9226 13319 -9192
rect 13353 -9226 13391 -9192
rect 13425 -9226 13463 -9192
rect 13497 -9226 13535 -9192
rect 13569 -9226 13607 -9192
rect 13641 -9226 13679 -9192
rect 13713 -9226 13751 -9192
rect 13785 -9226 13823 -9192
rect 13857 -9226 14040 -9192
rect 14074 -9226 14112 -9192
rect 14146 -9226 14184 -9192
rect 14218 -9226 14256 -9192
rect 14290 -9226 14328 -9192
rect 14362 -9226 14400 -9192
rect 14434 -9226 14472 -9192
rect 14506 -9226 14544 -9192
rect 14578 -9226 14616 -9192
rect 14650 -9226 14688 -9192
rect 14722 -9226 14760 -9192
rect 14794 -9226 14832 -9192
rect 14866 -9226 14904 -9192
rect 14938 -9226 14976 -9192
rect 15010 -9226 15048 -9192
rect 15082 -9226 15120 -9192
rect 15154 -9226 15192 -9192
rect 15226 -9226 15264 -9192
rect 15298 -9226 15336 -9192
rect 15370 -9226 15408 -9192
rect 15442 -9226 15480 -9192
rect 15514 -9226 15552 -9192
rect 15586 -9226 15624 -9192
rect 15658 -9226 15696 -9192
rect 15730 -9226 15768 -9192
rect 15802 -9226 15840 -9192
rect 15874 -9226 15912 -9192
rect 15946 -9226 15984 -9192
rect 16018 -9226 16056 -9192
rect 16090 -9226 16128 -9192
rect 16162 -9226 16200 -9192
rect 16234 -9226 16272 -9192
rect 16306 -9226 16344 -9192
rect 16378 -9226 16416 -9192
rect 16450 -9226 16488 -9192
rect 16522 -9226 16560 -9192
rect 16594 -9226 16632 -9192
rect 16666 -9226 16704 -9192
rect 16738 -9226 16776 -9192
rect 16810 -9226 16848 -9192
rect 16882 -9226 16920 -9192
rect 16954 -9226 16992 -9192
rect 17026 -9226 17064 -9192
rect 17098 -9226 17136 -9192
rect 17170 -9226 17208 -9192
rect 17242 -9226 17280 -9192
rect 17314 -9226 17352 -9192
rect 17386 -9226 17424 -9192
rect 17458 -9226 17496 -9192
rect 17530 -9226 17568 -9192
rect 17602 -9226 17640 -9192
rect 17674 -9226 17712 -9192
rect 17746 -9226 17784 -9192
rect 17818 -9226 17856 -9192
rect 17890 -9226 17928 -9192
rect 17962 -9226 18000 -9192
rect 18034 -9226 18072 -9192
rect 18106 -9226 18144 -9192
rect 18178 -9226 18216 -9192
rect 18250 -9226 18349 -9192
rect 831 -9251 18349 -9226
<< via1 >>
rect 2834 -64 2886 -12
rect 2898 -64 2950 -12
rect 2962 -64 3014 -12
rect 3351 -64 3403 -12
rect 3415 -64 3467 -12
rect 3479 -64 3531 -12
rect 1348 -233 1400 -181
rect 1412 -233 1464 -181
rect 1476 -233 1528 -181
rect 1865 -233 1917 -181
rect 1929 -233 1981 -181
rect 1993 -233 2045 -181
rect 2382 -233 2434 -181
rect 2446 -233 2498 -181
rect 2510 -233 2562 -181
rect 1607 -564 1659 -512
rect 1671 -564 1723 -512
rect 1735 -564 1787 -512
rect 2125 -564 2177 -512
rect 2189 -564 2241 -512
rect 2253 -564 2305 -512
rect 2577 -396 2629 -344
rect 2641 -396 2693 -344
rect 2705 -396 2757 -344
rect 3094 -396 3146 -344
rect 3158 -396 3210 -344
rect 3222 -396 3274 -344
rect 6931 -64 6983 -12
rect 6995 -64 7047 -12
rect 7059 -64 7111 -12
rect 7449 -64 7501 -12
rect 7513 -64 7565 -12
rect 7577 -64 7629 -12
rect 3543 -233 3595 -181
rect 3607 -233 3659 -181
rect 3671 -233 3723 -181
rect 4060 -233 4112 -181
rect 4124 -233 4176 -181
rect 4188 -233 4240 -181
rect 4575 -233 4627 -181
rect 4639 -233 4691 -181
rect 4703 -233 4755 -181
rect 3802 -564 3854 -512
rect 3866 -564 3918 -512
rect 3930 -564 3982 -512
rect 4319 -564 4371 -512
rect 4383 -564 4435 -512
rect 4447 -564 4499 -512
rect 5708 -233 5760 -181
rect 5772 -233 5824 -181
rect 5836 -233 5888 -181
rect 6223 -233 6275 -181
rect 6287 -233 6339 -181
rect 6351 -233 6403 -181
rect 6740 -233 6792 -181
rect 6804 -233 6856 -181
rect 6868 -233 6920 -181
rect 5964 -564 6016 -512
rect 6028 -564 6080 -512
rect 6092 -564 6144 -512
rect 6481 -564 6533 -512
rect 6545 -564 6597 -512
rect 6609 -564 6661 -512
rect 7189 -396 7241 -344
rect 7253 -396 7305 -344
rect 7317 -396 7369 -344
rect 11551 -64 11603 -12
rect 11615 -64 11667 -12
rect 11679 -64 11731 -12
rect 12069 -64 12121 -12
rect 12133 -64 12185 -12
rect 12197 -64 12249 -12
rect 7901 -233 7953 -181
rect 7965 -233 8017 -181
rect 8029 -233 8081 -181
rect 8417 -233 8469 -181
rect 8481 -233 8533 -181
rect 8545 -233 8597 -181
rect 8935 -233 8987 -181
rect 8999 -233 9051 -181
rect 9063 -233 9115 -181
rect 7706 -396 7758 -344
rect 7770 -396 7822 -344
rect 7834 -396 7886 -344
rect 8158 -564 8210 -512
rect 8222 -564 8274 -512
rect 8286 -564 8338 -512
rect 8675 -564 8727 -512
rect 8739 -564 8791 -512
rect 8803 -564 8855 -512
rect 10065 -233 10117 -181
rect 10129 -233 10181 -181
rect 10193 -233 10245 -181
rect 10583 -233 10635 -181
rect 10647 -233 10699 -181
rect 10711 -233 10763 -181
rect 11099 -233 11151 -181
rect 11163 -233 11215 -181
rect 11227 -233 11279 -181
rect 1523 -957 1550 -936
rect 1550 -957 1575 -936
rect 1523 -988 1575 -957
rect 1587 -957 1588 -936
rect 1588 -957 1622 -936
rect 1622 -957 1639 -936
rect 1587 -988 1639 -957
rect 1651 -988 1703 -936
rect 1719 -988 1771 -936
rect 1783 -957 1808 -936
rect 1808 -957 1835 -936
rect 1847 -957 1880 -936
rect 1880 -957 1899 -936
rect 1783 -988 1835 -957
rect 1847 -988 1899 -957
rect 2009 -957 2032 -936
rect 2032 -957 2061 -936
rect 2073 -957 2104 -936
rect 2104 -957 2125 -936
rect 2137 -957 2138 -936
rect 2138 -957 2189 -936
rect 2009 -988 2061 -957
rect 2073 -988 2125 -957
rect 2137 -988 2189 -957
rect 2205 -988 2257 -936
rect 2269 -957 2290 -936
rect 2290 -957 2321 -936
rect 2333 -957 2362 -936
rect 2362 -957 2385 -936
rect 2269 -988 2321 -957
rect 2333 -988 2385 -957
rect 1523 -1126 1575 -1074
rect 1587 -1126 1639 -1074
rect 1651 -1126 1703 -1074
rect 1719 -1126 1771 -1074
rect 1783 -1126 1835 -1074
rect 1847 -1126 1899 -1074
rect 2009 -1126 2061 -1074
rect 2073 -1126 2125 -1074
rect 2137 -1126 2189 -1074
rect 2205 -1126 2257 -1074
rect 2269 -1126 2321 -1074
rect 2333 -1126 2385 -1074
rect 1523 -1286 1575 -1252
rect 1523 -1304 1550 -1286
rect 1550 -1304 1575 -1286
rect 1587 -1286 1639 -1252
rect 1587 -1304 1588 -1286
rect 1588 -1304 1622 -1286
rect 1622 -1304 1639 -1286
rect 1651 -1304 1703 -1252
rect 1719 -1304 1771 -1252
rect 1783 -1286 1835 -1252
rect 1847 -1286 1899 -1252
rect 1783 -1304 1808 -1286
rect 1808 -1304 1835 -1286
rect 1847 -1304 1880 -1286
rect 1880 -1304 1899 -1286
rect 2009 -1286 2061 -1252
rect 2073 -1286 2125 -1252
rect 2137 -1286 2189 -1252
rect 2009 -1304 2032 -1286
rect 2032 -1304 2061 -1286
rect 2073 -1304 2104 -1286
rect 2104 -1304 2125 -1286
rect 2137 -1304 2138 -1286
rect 2138 -1304 2189 -1286
rect 2205 -1304 2257 -1252
rect 2269 -1286 2321 -1252
rect 2333 -1286 2385 -1252
rect 2269 -1304 2290 -1286
rect 2290 -1304 2321 -1286
rect 2333 -1304 2362 -1286
rect 2362 -1304 2385 -1286
rect 2733 -1126 2785 -1074
rect 2797 -1126 2849 -1074
rect 2861 -1126 2913 -1074
rect 2929 -1126 2981 -1074
rect 2993 -1126 3045 -1074
rect 3057 -1126 3109 -1074
rect 3121 -1126 3173 -1074
rect 3189 -1126 3241 -1074
rect 3253 -1126 3305 -1074
rect 3317 -1126 3369 -1074
rect 3721 -957 3744 -936
rect 3744 -957 3773 -936
rect 3785 -957 3816 -936
rect 3816 -957 3837 -936
rect 3721 -988 3773 -957
rect 3785 -988 3837 -957
rect 3849 -988 3901 -936
rect 3917 -957 3968 -936
rect 3968 -957 3969 -936
rect 3981 -957 4002 -936
rect 4002 -957 4033 -936
rect 4045 -957 4074 -936
rect 4074 -957 4097 -936
rect 3917 -988 3969 -957
rect 3981 -988 4033 -957
rect 4045 -988 4097 -957
rect 4207 -957 4226 -936
rect 4226 -957 4259 -936
rect 4271 -957 4298 -936
rect 4298 -957 4323 -936
rect 4207 -988 4259 -957
rect 4271 -988 4323 -957
rect 4335 -988 4387 -936
rect 4403 -988 4455 -936
rect 4467 -957 4484 -936
rect 4484 -957 4518 -936
rect 4518 -957 4519 -936
rect 4467 -988 4519 -957
rect 4531 -957 4556 -936
rect 4556 -957 4583 -936
rect 4531 -988 4583 -957
rect 10325 -564 10377 -512
rect 10389 -564 10441 -512
rect 10453 -564 10505 -512
rect 10842 -564 10894 -512
rect 10906 -564 10958 -512
rect 10970 -564 11022 -512
rect 11294 -396 11346 -344
rect 11358 -396 11410 -344
rect 11422 -396 11474 -344
rect 11811 -396 11863 -344
rect 11875 -396 11927 -344
rect 11939 -396 11991 -344
rect 15649 -64 15701 -12
rect 15713 -64 15765 -12
rect 15777 -64 15829 -12
rect 16166 -64 16218 -12
rect 16230 -64 16282 -12
rect 16294 -64 16346 -12
rect 12260 -233 12312 -181
rect 12324 -233 12376 -181
rect 12388 -233 12440 -181
rect 12777 -233 12829 -181
rect 12841 -233 12893 -181
rect 12905 -233 12957 -181
rect 13292 -233 13344 -181
rect 13356 -233 13408 -181
rect 13420 -233 13472 -181
rect 12519 -564 12571 -512
rect 12583 -564 12635 -512
rect 12647 -564 12699 -512
rect 13036 -564 13088 -512
rect 13100 -564 13152 -512
rect 13164 -564 13216 -512
rect 14425 -233 14477 -181
rect 14489 -233 14541 -181
rect 14553 -233 14605 -181
rect 14940 -233 14992 -181
rect 15004 -233 15056 -181
rect 15068 -233 15120 -181
rect 15457 -233 15509 -181
rect 15521 -233 15573 -181
rect 15585 -233 15637 -181
rect 5880 -957 5907 -936
rect 5907 -957 5932 -936
rect 5880 -988 5932 -957
rect 5944 -957 5945 -936
rect 5945 -957 5979 -936
rect 5979 -957 5996 -936
rect 5944 -988 5996 -957
rect 6008 -988 6060 -936
rect 6076 -988 6128 -936
rect 6140 -957 6165 -936
rect 6165 -957 6192 -936
rect 6204 -957 6237 -936
rect 6237 -957 6256 -936
rect 6140 -988 6192 -957
rect 6204 -988 6256 -957
rect 6366 -957 6389 -936
rect 6389 -957 6418 -936
rect 6430 -957 6461 -936
rect 6461 -957 6482 -936
rect 6494 -957 6495 -936
rect 6495 -957 6546 -936
rect 6366 -988 6418 -957
rect 6430 -988 6482 -957
rect 6494 -988 6546 -957
rect 6562 -988 6614 -936
rect 6626 -957 6647 -936
rect 6647 -957 6678 -936
rect 6690 -957 6719 -936
rect 6719 -957 6742 -936
rect 6626 -988 6678 -957
rect 6690 -988 6742 -957
rect 3721 -1126 3773 -1074
rect 3785 -1126 3837 -1074
rect 3849 -1126 3901 -1074
rect 3917 -1126 3969 -1074
rect 3981 -1126 4033 -1074
rect 4045 -1126 4097 -1074
rect 4207 -1126 4259 -1074
rect 4271 -1126 4323 -1074
rect 4335 -1126 4387 -1074
rect 4403 -1126 4455 -1074
rect 4467 -1126 4519 -1074
rect 4531 -1126 4583 -1074
rect 3721 -1286 3773 -1252
rect 3785 -1286 3837 -1252
rect 3721 -1304 3744 -1286
rect 3744 -1304 3773 -1286
rect 3785 -1304 3816 -1286
rect 3816 -1304 3837 -1286
rect 3849 -1304 3901 -1252
rect 3917 -1286 3969 -1252
rect 3981 -1286 4033 -1252
rect 4045 -1286 4097 -1252
rect 3917 -1304 3968 -1286
rect 3968 -1304 3969 -1286
rect 3981 -1304 4002 -1286
rect 4002 -1304 4033 -1286
rect 4045 -1304 4074 -1286
rect 4074 -1304 4097 -1286
rect 4207 -1286 4259 -1252
rect 4271 -1286 4323 -1252
rect 4207 -1304 4226 -1286
rect 4226 -1304 4259 -1286
rect 4271 -1304 4298 -1286
rect 4298 -1304 4323 -1286
rect 4335 -1304 4387 -1252
rect 4403 -1304 4455 -1252
rect 4467 -1286 4519 -1252
rect 4467 -1304 4484 -1286
rect 4484 -1304 4518 -1286
rect 4518 -1304 4519 -1286
rect 4531 -1286 4583 -1252
rect 4531 -1304 4556 -1286
rect 4556 -1304 4583 -1286
rect 5880 -1126 5932 -1074
rect 5944 -1126 5996 -1074
rect 6008 -1126 6060 -1074
rect 6076 -1126 6128 -1074
rect 6140 -1126 6192 -1074
rect 6204 -1126 6256 -1074
rect 6366 -1126 6418 -1074
rect 6430 -1126 6482 -1074
rect 6494 -1126 6546 -1074
rect 6562 -1126 6614 -1074
rect 6626 -1126 6678 -1074
rect 6690 -1126 6742 -1074
rect 5880 -1286 5932 -1252
rect 5880 -1304 5907 -1286
rect 5907 -1304 5932 -1286
rect 5944 -1286 5996 -1252
rect 5944 -1304 5945 -1286
rect 5945 -1304 5979 -1286
rect 5979 -1304 5996 -1286
rect 6008 -1304 6060 -1252
rect 6076 -1304 6128 -1252
rect 6140 -1286 6192 -1252
rect 6204 -1286 6256 -1252
rect 6140 -1304 6165 -1286
rect 6165 -1304 6192 -1286
rect 6204 -1304 6237 -1286
rect 6237 -1304 6256 -1286
rect 6366 -1286 6418 -1252
rect 6430 -1286 6482 -1252
rect 6494 -1286 6546 -1252
rect 6366 -1304 6389 -1286
rect 6389 -1304 6418 -1286
rect 6430 -1304 6461 -1286
rect 6461 -1304 6482 -1286
rect 6494 -1304 6495 -1286
rect 6495 -1304 6546 -1286
rect 6562 -1304 6614 -1252
rect 6626 -1286 6678 -1252
rect 6690 -1286 6742 -1252
rect 6626 -1304 6647 -1286
rect 6647 -1304 6678 -1286
rect 6690 -1304 6719 -1286
rect 6719 -1304 6742 -1286
rect 7094 -1126 7146 -1074
rect 7158 -1126 7210 -1074
rect 7222 -1126 7274 -1074
rect 7290 -1126 7342 -1074
rect 7354 -1126 7406 -1074
rect 7418 -1126 7470 -1074
rect 7482 -1126 7534 -1074
rect 7550 -1126 7602 -1074
rect 7614 -1126 7666 -1074
rect 7678 -1126 7730 -1074
rect 8078 -957 8101 -936
rect 8101 -957 8130 -936
rect 8142 -957 8173 -936
rect 8173 -957 8194 -936
rect 8078 -988 8130 -957
rect 8142 -988 8194 -957
rect 8206 -988 8258 -936
rect 8274 -957 8325 -936
rect 8325 -957 8326 -936
rect 8338 -957 8359 -936
rect 8359 -957 8390 -936
rect 8402 -957 8431 -936
rect 8431 -957 8454 -936
rect 8274 -988 8326 -957
rect 8338 -988 8390 -957
rect 8402 -988 8454 -957
rect 8564 -957 8583 -936
rect 8583 -957 8616 -936
rect 8628 -957 8655 -936
rect 8655 -957 8680 -936
rect 8564 -988 8616 -957
rect 8628 -988 8680 -957
rect 8692 -988 8744 -936
rect 8760 -988 8812 -936
rect 8824 -957 8841 -936
rect 8841 -957 8875 -936
rect 8875 -957 8876 -936
rect 8824 -988 8876 -957
rect 8888 -957 8913 -936
rect 8913 -957 8940 -936
rect 8888 -988 8940 -957
rect 14681 -564 14733 -512
rect 14745 -564 14797 -512
rect 14809 -564 14861 -512
rect 15198 -564 15250 -512
rect 15262 -564 15314 -512
rect 15326 -564 15378 -512
rect 15906 -396 15958 -344
rect 15970 -396 16022 -344
rect 16034 -396 16086 -344
rect 16618 -233 16670 -181
rect 16682 -233 16734 -181
rect 16746 -233 16798 -181
rect 17135 -233 17187 -181
rect 17199 -233 17251 -181
rect 17263 -233 17315 -181
rect 17652 -233 17704 -181
rect 17716 -233 17768 -181
rect 17780 -233 17832 -181
rect 16423 -396 16475 -344
rect 16487 -396 16539 -344
rect 16551 -396 16603 -344
rect 16875 -564 16927 -512
rect 16939 -564 16991 -512
rect 17003 -564 17055 -512
rect 17393 -564 17445 -512
rect 17457 -564 17509 -512
rect 17521 -564 17573 -512
rect 10240 -957 10267 -936
rect 10267 -957 10292 -936
rect 10240 -988 10292 -957
rect 10304 -957 10305 -936
rect 10305 -957 10339 -936
rect 10339 -957 10356 -936
rect 10304 -988 10356 -957
rect 10368 -988 10420 -936
rect 10436 -988 10488 -936
rect 10500 -957 10525 -936
rect 10525 -957 10552 -936
rect 10564 -957 10597 -936
rect 10597 -957 10616 -936
rect 10500 -988 10552 -957
rect 10564 -988 10616 -957
rect 10726 -957 10749 -936
rect 10749 -957 10778 -936
rect 10790 -957 10821 -936
rect 10821 -957 10842 -936
rect 10854 -957 10855 -936
rect 10855 -957 10906 -936
rect 10726 -988 10778 -957
rect 10790 -988 10842 -957
rect 10854 -988 10906 -957
rect 10922 -988 10974 -936
rect 10986 -957 11007 -936
rect 11007 -957 11038 -936
rect 11050 -957 11079 -936
rect 11079 -957 11102 -936
rect 10986 -988 11038 -957
rect 11050 -988 11102 -957
rect 8078 -1126 8130 -1074
rect 8142 -1126 8194 -1074
rect 8206 -1126 8258 -1074
rect 8274 -1126 8326 -1074
rect 8338 -1126 8390 -1074
rect 8402 -1126 8454 -1074
rect 8564 -1126 8616 -1074
rect 8628 -1126 8680 -1074
rect 8692 -1126 8744 -1074
rect 8760 -1126 8812 -1074
rect 8824 -1126 8876 -1074
rect 8888 -1126 8940 -1074
rect 8078 -1286 8130 -1252
rect 8142 -1286 8194 -1252
rect 8078 -1304 8101 -1286
rect 8101 -1304 8130 -1286
rect 8142 -1304 8173 -1286
rect 8173 -1304 8194 -1286
rect 8206 -1304 8258 -1252
rect 8274 -1286 8326 -1252
rect 8338 -1286 8390 -1252
rect 8402 -1286 8454 -1252
rect 8274 -1304 8325 -1286
rect 8325 -1304 8326 -1286
rect 8338 -1304 8359 -1286
rect 8359 -1304 8390 -1286
rect 8402 -1304 8431 -1286
rect 8431 -1304 8454 -1286
rect 8564 -1286 8616 -1252
rect 8628 -1286 8680 -1252
rect 8564 -1304 8583 -1286
rect 8583 -1304 8616 -1286
rect 8628 -1304 8655 -1286
rect 8655 -1304 8680 -1286
rect 8692 -1304 8744 -1252
rect 8760 -1304 8812 -1252
rect 8824 -1286 8876 -1252
rect 8824 -1304 8841 -1286
rect 8841 -1304 8875 -1286
rect 8875 -1304 8876 -1286
rect 8888 -1286 8940 -1252
rect 8888 -1304 8913 -1286
rect 8913 -1304 8940 -1286
rect 1350 -1754 1402 -1702
rect 1414 -1754 1466 -1702
rect 1478 -1754 1530 -1702
rect 1865 -1754 1917 -1702
rect 1929 -1754 1981 -1702
rect 1993 -1754 2045 -1702
rect 1608 -2055 1660 -2003
rect 1672 -2055 1724 -2003
rect 1736 -2055 1788 -2003
rect 2383 -1754 2435 -1702
rect 2447 -1754 2499 -1702
rect 2511 -1754 2563 -1702
rect 2126 -2055 2178 -2003
rect 2190 -2055 2242 -2003
rect 2254 -2055 2306 -2003
rect 2833 -1894 2885 -1842
rect 2897 -1894 2949 -1842
rect 2961 -1894 3013 -1842
rect 2575 -2199 2627 -2147
rect 2639 -2199 2691 -2147
rect 2703 -2199 2755 -2147
rect 3543 -1754 3595 -1702
rect 3607 -1754 3659 -1702
rect 3671 -1754 3723 -1702
rect 3350 -1894 3402 -1842
rect 3414 -1894 3466 -1842
rect 3478 -1894 3530 -1842
rect 3092 -2199 3144 -2147
rect 3156 -2199 3208 -2147
rect 3220 -2199 3272 -2147
rect 4060 -1754 4112 -1702
rect 4124 -1754 4176 -1702
rect 4188 -1754 4240 -1702
rect 3803 -2055 3855 -2003
rect 3867 -2055 3919 -2003
rect 3931 -2055 3983 -2003
rect 10240 -1126 10292 -1074
rect 10304 -1126 10356 -1074
rect 10368 -1126 10420 -1074
rect 10436 -1126 10488 -1074
rect 10500 -1126 10552 -1074
rect 10564 -1126 10616 -1074
rect 10726 -1126 10778 -1074
rect 10790 -1126 10842 -1074
rect 10854 -1126 10906 -1074
rect 10922 -1126 10974 -1074
rect 10986 -1126 11038 -1074
rect 11050 -1126 11102 -1074
rect 10240 -1286 10292 -1252
rect 10240 -1304 10267 -1286
rect 10267 -1304 10292 -1286
rect 10304 -1286 10356 -1252
rect 10304 -1304 10305 -1286
rect 10305 -1304 10339 -1286
rect 10339 -1304 10356 -1286
rect 10368 -1304 10420 -1252
rect 10436 -1304 10488 -1252
rect 10500 -1286 10552 -1252
rect 10564 -1286 10616 -1252
rect 10500 -1304 10525 -1286
rect 10525 -1304 10552 -1286
rect 10564 -1304 10597 -1286
rect 10597 -1304 10616 -1286
rect 10726 -1286 10778 -1252
rect 10790 -1286 10842 -1252
rect 10854 -1286 10906 -1252
rect 10726 -1304 10749 -1286
rect 10749 -1304 10778 -1286
rect 10790 -1304 10821 -1286
rect 10821 -1304 10842 -1286
rect 10854 -1304 10855 -1286
rect 10855 -1304 10906 -1286
rect 10922 -1304 10974 -1252
rect 10986 -1286 11038 -1252
rect 11050 -1286 11102 -1252
rect 10986 -1304 11007 -1286
rect 11007 -1304 11038 -1286
rect 11050 -1304 11079 -1286
rect 11079 -1304 11102 -1286
rect 11450 -1126 11502 -1074
rect 11514 -1126 11566 -1074
rect 11578 -1126 11630 -1074
rect 11646 -1126 11698 -1074
rect 11710 -1126 11762 -1074
rect 11774 -1126 11826 -1074
rect 11838 -1126 11890 -1074
rect 11906 -1126 11958 -1074
rect 11970 -1126 12022 -1074
rect 12034 -1126 12086 -1074
rect 12438 -957 12461 -936
rect 12461 -957 12490 -936
rect 12502 -957 12533 -936
rect 12533 -957 12554 -936
rect 12438 -988 12490 -957
rect 12502 -988 12554 -957
rect 12566 -988 12618 -936
rect 12634 -957 12685 -936
rect 12685 -957 12686 -936
rect 12698 -957 12719 -936
rect 12719 -957 12750 -936
rect 12762 -957 12791 -936
rect 12791 -957 12814 -936
rect 12634 -988 12686 -957
rect 12698 -988 12750 -957
rect 12762 -988 12814 -957
rect 12924 -957 12943 -936
rect 12943 -957 12976 -936
rect 12988 -957 13015 -936
rect 13015 -957 13040 -936
rect 12924 -988 12976 -957
rect 12988 -988 13040 -957
rect 13052 -988 13104 -936
rect 13120 -988 13172 -936
rect 13184 -957 13201 -936
rect 13201 -957 13235 -936
rect 13235 -957 13236 -936
rect 13184 -988 13236 -957
rect 13248 -957 13273 -936
rect 13273 -957 13300 -936
rect 13248 -988 13300 -957
rect 14597 -957 14624 -936
rect 14624 -957 14649 -936
rect 14597 -988 14649 -957
rect 14661 -957 14662 -936
rect 14662 -957 14696 -936
rect 14696 -957 14713 -936
rect 14661 -988 14713 -957
rect 14725 -988 14777 -936
rect 14793 -988 14845 -936
rect 14857 -957 14882 -936
rect 14882 -957 14909 -936
rect 14921 -957 14954 -936
rect 14954 -957 14973 -936
rect 14857 -988 14909 -957
rect 14921 -988 14973 -957
rect 15083 -957 15106 -936
rect 15106 -957 15135 -936
rect 15147 -957 15178 -936
rect 15178 -957 15199 -936
rect 15211 -957 15212 -936
rect 15212 -957 15263 -936
rect 15083 -988 15135 -957
rect 15147 -988 15199 -957
rect 15211 -988 15263 -957
rect 15279 -988 15331 -936
rect 15343 -957 15364 -936
rect 15364 -957 15395 -936
rect 15407 -957 15436 -936
rect 15436 -957 15459 -936
rect 15343 -988 15395 -957
rect 15407 -988 15459 -957
rect 12438 -1126 12490 -1074
rect 12502 -1126 12554 -1074
rect 12566 -1126 12618 -1074
rect 12634 -1126 12686 -1074
rect 12698 -1126 12750 -1074
rect 12762 -1126 12814 -1074
rect 12924 -1126 12976 -1074
rect 12988 -1126 13040 -1074
rect 13052 -1126 13104 -1074
rect 13120 -1126 13172 -1074
rect 13184 -1126 13236 -1074
rect 13248 -1126 13300 -1074
rect 12438 -1286 12490 -1252
rect 12502 -1286 12554 -1252
rect 12438 -1304 12461 -1286
rect 12461 -1304 12490 -1286
rect 12502 -1304 12533 -1286
rect 12533 -1304 12554 -1286
rect 12566 -1304 12618 -1252
rect 12634 -1286 12686 -1252
rect 12698 -1286 12750 -1252
rect 12762 -1286 12814 -1252
rect 12634 -1304 12685 -1286
rect 12685 -1304 12686 -1286
rect 12698 -1304 12719 -1286
rect 12719 -1304 12750 -1286
rect 12762 -1304 12791 -1286
rect 12791 -1304 12814 -1286
rect 12924 -1286 12976 -1252
rect 12988 -1286 13040 -1252
rect 12924 -1304 12943 -1286
rect 12943 -1304 12976 -1286
rect 12988 -1304 13015 -1286
rect 13015 -1304 13040 -1286
rect 13052 -1304 13104 -1252
rect 13120 -1304 13172 -1252
rect 13184 -1286 13236 -1252
rect 13184 -1304 13201 -1286
rect 13201 -1304 13235 -1286
rect 13235 -1304 13236 -1286
rect 13248 -1286 13300 -1252
rect 13248 -1304 13273 -1286
rect 13273 -1304 13300 -1286
rect 4577 -1754 4629 -1702
rect 4641 -1754 4693 -1702
rect 4705 -1754 4757 -1702
rect 4320 -2055 4372 -2003
rect 4384 -2055 4436 -2003
rect 4448 -2055 4500 -2003
rect 5706 -1754 5758 -1702
rect 5770 -1754 5822 -1702
rect 5834 -1754 5886 -1702
rect 6223 -1754 6275 -1702
rect 6287 -1754 6339 -1702
rect 6351 -1754 6403 -1702
rect 5963 -2055 6015 -2003
rect 6027 -2055 6079 -2003
rect 6091 -2055 6143 -2003
rect 6740 -1754 6792 -1702
rect 6804 -1754 6856 -1702
rect 6868 -1754 6920 -1702
rect 6480 -2055 6532 -2003
rect 6544 -2055 6596 -2003
rect 6608 -2055 6660 -2003
rect 6933 -1894 6985 -1842
rect 6997 -1894 7049 -1842
rect 7061 -1894 7113 -1842
rect 7450 -1894 7502 -1842
rect 7514 -1894 7566 -1842
rect 7578 -1894 7630 -1842
rect 7191 -2199 7243 -2147
rect 7255 -2199 7307 -2147
rect 7319 -2199 7371 -2147
rect 7900 -1754 7952 -1702
rect 7964 -1754 8016 -1702
rect 8028 -1754 8080 -1702
rect 7708 -2199 7760 -2147
rect 7772 -2199 7824 -2147
rect 7836 -2199 7888 -2147
rect 8417 -1754 8469 -1702
rect 8481 -1754 8533 -1702
rect 8545 -1754 8597 -1702
rect 8157 -2055 8209 -2003
rect 8221 -2055 8273 -2003
rect 8285 -2055 8337 -2003
rect 14597 -1126 14649 -1074
rect 14661 -1126 14713 -1074
rect 14725 -1126 14777 -1074
rect 14793 -1126 14845 -1074
rect 14857 -1126 14909 -1074
rect 14921 -1126 14973 -1074
rect 15083 -1126 15135 -1074
rect 15147 -1126 15199 -1074
rect 15211 -1126 15263 -1074
rect 15279 -1126 15331 -1074
rect 15343 -1126 15395 -1074
rect 15407 -1126 15459 -1074
rect 14597 -1286 14649 -1252
rect 14597 -1304 14624 -1286
rect 14624 -1304 14649 -1286
rect 14661 -1286 14713 -1252
rect 14661 -1304 14662 -1286
rect 14662 -1304 14696 -1286
rect 14696 -1304 14713 -1286
rect 14725 -1304 14777 -1252
rect 14793 -1304 14845 -1252
rect 14857 -1286 14909 -1252
rect 14921 -1286 14973 -1252
rect 14857 -1304 14882 -1286
rect 14882 -1304 14909 -1286
rect 14921 -1304 14954 -1286
rect 14954 -1304 14973 -1286
rect 15083 -1286 15135 -1252
rect 15147 -1286 15199 -1252
rect 15211 -1286 15263 -1252
rect 15083 -1304 15106 -1286
rect 15106 -1304 15135 -1286
rect 15147 -1304 15178 -1286
rect 15178 -1304 15199 -1286
rect 15211 -1304 15212 -1286
rect 15212 -1304 15263 -1286
rect 15279 -1304 15331 -1252
rect 15343 -1286 15395 -1252
rect 15407 -1286 15459 -1252
rect 15343 -1304 15364 -1286
rect 15364 -1304 15395 -1286
rect 15407 -1304 15436 -1286
rect 15436 -1304 15459 -1286
rect 15811 -1126 15863 -1074
rect 15875 -1126 15927 -1074
rect 15939 -1126 15991 -1074
rect 16007 -1126 16059 -1074
rect 16071 -1126 16123 -1074
rect 16135 -1126 16187 -1074
rect 16199 -1126 16251 -1074
rect 16267 -1126 16319 -1074
rect 16331 -1126 16383 -1074
rect 16395 -1126 16447 -1074
rect 16795 -957 16818 -936
rect 16818 -957 16847 -936
rect 16859 -957 16890 -936
rect 16890 -957 16911 -936
rect 16795 -988 16847 -957
rect 16859 -988 16911 -957
rect 16923 -988 16975 -936
rect 16991 -957 17042 -936
rect 17042 -957 17043 -936
rect 17055 -957 17076 -936
rect 17076 -957 17107 -936
rect 17119 -957 17148 -936
rect 17148 -957 17171 -936
rect 16991 -988 17043 -957
rect 17055 -988 17107 -957
rect 17119 -988 17171 -957
rect 17281 -957 17300 -936
rect 17300 -957 17333 -936
rect 17345 -957 17372 -936
rect 17372 -957 17397 -936
rect 17281 -988 17333 -957
rect 17345 -988 17397 -957
rect 17409 -988 17461 -936
rect 17477 -988 17529 -936
rect 17541 -957 17558 -936
rect 17558 -957 17592 -936
rect 17592 -957 17593 -936
rect 17541 -988 17593 -957
rect 17605 -957 17630 -936
rect 17630 -957 17657 -936
rect 17605 -988 17657 -957
rect 16795 -1126 16847 -1074
rect 16859 -1126 16911 -1074
rect 16923 -1126 16975 -1074
rect 16991 -1126 17043 -1074
rect 17055 -1126 17107 -1074
rect 17119 -1126 17171 -1074
rect 17281 -1126 17333 -1074
rect 17345 -1126 17397 -1074
rect 17409 -1126 17461 -1074
rect 17477 -1126 17529 -1074
rect 17541 -1126 17593 -1074
rect 17605 -1126 17657 -1074
rect 16795 -1286 16847 -1252
rect 16859 -1286 16911 -1252
rect 16795 -1304 16818 -1286
rect 16818 -1304 16847 -1286
rect 16859 -1304 16890 -1286
rect 16890 -1304 16911 -1286
rect 16923 -1304 16975 -1252
rect 16991 -1286 17043 -1252
rect 17055 -1286 17107 -1252
rect 17119 -1286 17171 -1252
rect 16991 -1304 17042 -1286
rect 17042 -1304 17043 -1286
rect 17055 -1304 17076 -1286
rect 17076 -1304 17107 -1286
rect 17119 -1304 17148 -1286
rect 17148 -1304 17171 -1286
rect 17281 -1286 17333 -1252
rect 17345 -1286 17397 -1252
rect 17281 -1304 17300 -1286
rect 17300 -1304 17333 -1286
rect 17345 -1304 17372 -1286
rect 17372 -1304 17397 -1286
rect 17409 -1304 17461 -1252
rect 17477 -1304 17529 -1252
rect 17541 -1286 17593 -1252
rect 17541 -1304 17558 -1286
rect 17558 -1304 17592 -1286
rect 17592 -1304 17593 -1286
rect 17605 -1286 17657 -1252
rect 17605 -1304 17630 -1286
rect 17630 -1304 17657 -1286
rect 8932 -1754 8984 -1702
rect 8996 -1754 9048 -1702
rect 9060 -1754 9112 -1702
rect 8674 -2055 8726 -2003
rect 8738 -2055 8790 -2003
rect 8802 -2055 8854 -2003
rect 10068 -1754 10120 -1702
rect 10132 -1754 10184 -1702
rect 10196 -1754 10248 -1702
rect 1523 -2604 1550 -2583
rect 1550 -2604 1575 -2583
rect 1523 -2635 1575 -2604
rect 1587 -2604 1588 -2583
rect 1588 -2604 1622 -2583
rect 1622 -2604 1639 -2583
rect 1587 -2635 1639 -2604
rect 1651 -2635 1703 -2583
rect 1719 -2635 1771 -2583
rect 1783 -2604 1808 -2583
rect 1808 -2604 1835 -2583
rect 1847 -2604 1880 -2583
rect 1880 -2604 1899 -2583
rect 1783 -2635 1835 -2604
rect 1847 -2635 1899 -2604
rect 2009 -2604 2032 -2583
rect 2032 -2604 2061 -2583
rect 2073 -2604 2104 -2583
rect 2104 -2604 2125 -2583
rect 2137 -2604 2138 -2583
rect 2138 -2604 2189 -2583
rect 2009 -2635 2061 -2604
rect 2073 -2635 2125 -2604
rect 2137 -2635 2189 -2604
rect 2205 -2635 2257 -2583
rect 2269 -2604 2290 -2583
rect 2290 -2604 2321 -2583
rect 2333 -2604 2362 -2583
rect 2362 -2604 2385 -2583
rect 2269 -2635 2321 -2604
rect 2333 -2635 2385 -2604
rect 1523 -2773 1575 -2721
rect 1587 -2773 1639 -2721
rect 1651 -2773 1703 -2721
rect 1719 -2773 1771 -2721
rect 1783 -2773 1835 -2721
rect 1847 -2773 1899 -2721
rect 2009 -2773 2061 -2721
rect 2073 -2773 2125 -2721
rect 2137 -2773 2189 -2721
rect 2205 -2773 2257 -2721
rect 2269 -2773 2321 -2721
rect 2333 -2773 2385 -2721
rect 1523 -2933 1575 -2899
rect 1523 -2951 1550 -2933
rect 1550 -2951 1575 -2933
rect 1587 -2933 1639 -2899
rect 1587 -2951 1588 -2933
rect 1588 -2951 1622 -2933
rect 1622 -2951 1639 -2933
rect 1651 -2951 1703 -2899
rect 1719 -2951 1771 -2899
rect 1783 -2933 1835 -2899
rect 1847 -2933 1899 -2899
rect 1783 -2951 1808 -2933
rect 1808 -2951 1835 -2933
rect 1847 -2951 1880 -2933
rect 1880 -2951 1899 -2933
rect 2009 -2933 2061 -2899
rect 2073 -2933 2125 -2899
rect 2137 -2933 2189 -2899
rect 2009 -2951 2032 -2933
rect 2032 -2951 2061 -2933
rect 2073 -2951 2104 -2933
rect 2104 -2951 2125 -2933
rect 2137 -2951 2138 -2933
rect 2138 -2951 2189 -2933
rect 2205 -2951 2257 -2899
rect 2269 -2933 2321 -2899
rect 2333 -2933 2385 -2899
rect 2269 -2951 2290 -2933
rect 2290 -2951 2321 -2933
rect 2333 -2951 2362 -2933
rect 2362 -2951 2385 -2933
rect 2733 -2773 2785 -2721
rect 2797 -2773 2849 -2721
rect 2861 -2773 2913 -2721
rect 2929 -2773 2981 -2721
rect 2993 -2773 3045 -2721
rect 3057 -2773 3109 -2721
rect 3121 -2773 3173 -2721
rect 3189 -2773 3241 -2721
rect 3253 -2773 3305 -2721
rect 3317 -2773 3369 -2721
rect 3721 -2604 3744 -2583
rect 3744 -2604 3773 -2583
rect 3785 -2604 3816 -2583
rect 3816 -2604 3837 -2583
rect 3721 -2635 3773 -2604
rect 3785 -2635 3837 -2604
rect 3849 -2635 3901 -2583
rect 3917 -2604 3968 -2583
rect 3968 -2604 3969 -2583
rect 3981 -2604 4002 -2583
rect 4002 -2604 4033 -2583
rect 4045 -2604 4074 -2583
rect 4074 -2604 4097 -2583
rect 3917 -2635 3969 -2604
rect 3981 -2635 4033 -2604
rect 4045 -2635 4097 -2604
rect 4207 -2604 4226 -2583
rect 4226 -2604 4259 -2583
rect 4271 -2604 4298 -2583
rect 4298 -2604 4323 -2583
rect 4207 -2635 4259 -2604
rect 4271 -2635 4323 -2604
rect 4335 -2635 4387 -2583
rect 4403 -2635 4455 -2583
rect 4467 -2604 4484 -2583
rect 4484 -2604 4518 -2583
rect 4518 -2604 4519 -2583
rect 4467 -2635 4519 -2604
rect 4531 -2604 4556 -2583
rect 4556 -2604 4583 -2583
rect 4531 -2635 4583 -2604
rect 10583 -1754 10635 -1702
rect 10647 -1754 10699 -1702
rect 10711 -1754 10763 -1702
rect 10326 -2055 10378 -2003
rect 10390 -2055 10442 -2003
rect 10454 -2055 10506 -2003
rect 11100 -1754 11152 -1702
rect 11164 -1754 11216 -1702
rect 11228 -1754 11280 -1702
rect 10843 -2055 10895 -2003
rect 10907 -2055 10959 -2003
rect 10971 -2055 11023 -2003
rect 11550 -1894 11602 -1842
rect 11614 -1894 11666 -1842
rect 11678 -1894 11730 -1842
rect 11292 -2199 11344 -2147
rect 11356 -2199 11408 -2147
rect 11420 -2199 11472 -2147
rect 12260 -1754 12312 -1702
rect 12324 -1754 12376 -1702
rect 12388 -1754 12440 -1702
rect 12067 -1894 12119 -1842
rect 12131 -1894 12183 -1842
rect 12195 -1894 12247 -1842
rect 11809 -2199 11861 -2147
rect 11873 -2199 11925 -2147
rect 11937 -2199 11989 -2147
rect 12777 -1754 12829 -1702
rect 12841 -1754 12893 -1702
rect 12905 -1754 12957 -1702
rect 12520 -2055 12572 -2003
rect 12584 -2055 12636 -2003
rect 12648 -2055 12700 -2003
rect 13294 -1754 13346 -1702
rect 13358 -1754 13410 -1702
rect 13422 -1754 13474 -1702
rect 13037 -2055 13089 -2003
rect 13101 -2055 13153 -2003
rect 13165 -2055 13217 -2003
rect 14423 -1754 14475 -1702
rect 14487 -1754 14539 -1702
rect 14551 -1754 14603 -1702
rect 5880 -2604 5907 -2583
rect 5907 -2604 5932 -2583
rect 5880 -2635 5932 -2604
rect 5944 -2604 5945 -2583
rect 5945 -2604 5979 -2583
rect 5979 -2604 5996 -2583
rect 5944 -2635 5996 -2604
rect 6008 -2635 6060 -2583
rect 6076 -2635 6128 -2583
rect 6140 -2604 6165 -2583
rect 6165 -2604 6192 -2583
rect 6204 -2604 6237 -2583
rect 6237 -2604 6256 -2583
rect 6140 -2635 6192 -2604
rect 6204 -2635 6256 -2604
rect 6366 -2604 6389 -2583
rect 6389 -2604 6418 -2583
rect 6430 -2604 6461 -2583
rect 6461 -2604 6482 -2583
rect 6494 -2604 6495 -2583
rect 6495 -2604 6546 -2583
rect 6366 -2635 6418 -2604
rect 6430 -2635 6482 -2604
rect 6494 -2635 6546 -2604
rect 6562 -2635 6614 -2583
rect 6626 -2604 6647 -2583
rect 6647 -2604 6678 -2583
rect 6690 -2604 6719 -2583
rect 6719 -2604 6742 -2583
rect 6626 -2635 6678 -2604
rect 6690 -2635 6742 -2604
rect 3721 -2773 3773 -2721
rect 3785 -2773 3837 -2721
rect 3849 -2773 3901 -2721
rect 3917 -2773 3969 -2721
rect 3981 -2773 4033 -2721
rect 4045 -2773 4097 -2721
rect 4207 -2773 4259 -2721
rect 4271 -2773 4323 -2721
rect 4335 -2773 4387 -2721
rect 4403 -2773 4455 -2721
rect 4467 -2773 4519 -2721
rect 4531 -2773 4583 -2721
rect 3721 -2933 3773 -2899
rect 3785 -2933 3837 -2899
rect 3721 -2951 3744 -2933
rect 3744 -2951 3773 -2933
rect 3785 -2951 3816 -2933
rect 3816 -2951 3837 -2933
rect 3849 -2951 3901 -2899
rect 3917 -2933 3969 -2899
rect 3981 -2933 4033 -2899
rect 4045 -2933 4097 -2899
rect 3917 -2951 3968 -2933
rect 3968 -2951 3969 -2933
rect 3981 -2951 4002 -2933
rect 4002 -2951 4033 -2933
rect 4045 -2951 4074 -2933
rect 4074 -2951 4097 -2933
rect 4207 -2933 4259 -2899
rect 4271 -2933 4323 -2899
rect 4207 -2951 4226 -2933
rect 4226 -2951 4259 -2933
rect 4271 -2951 4298 -2933
rect 4298 -2951 4323 -2933
rect 4335 -2951 4387 -2899
rect 4403 -2951 4455 -2899
rect 4467 -2933 4519 -2899
rect 4467 -2951 4484 -2933
rect 4484 -2951 4518 -2933
rect 4518 -2951 4519 -2933
rect 4531 -2933 4583 -2899
rect 4531 -2951 4556 -2933
rect 4556 -2951 4583 -2933
rect 5880 -2773 5932 -2721
rect 5944 -2773 5996 -2721
rect 6008 -2773 6060 -2721
rect 6076 -2773 6128 -2721
rect 6140 -2773 6192 -2721
rect 6204 -2773 6256 -2721
rect 6366 -2773 6418 -2721
rect 6430 -2773 6482 -2721
rect 6494 -2773 6546 -2721
rect 6562 -2773 6614 -2721
rect 6626 -2773 6678 -2721
rect 6690 -2773 6742 -2721
rect 5880 -2933 5932 -2899
rect 5880 -2951 5907 -2933
rect 5907 -2951 5932 -2933
rect 5944 -2933 5996 -2899
rect 5944 -2951 5945 -2933
rect 5945 -2951 5979 -2933
rect 5979 -2951 5996 -2933
rect 6008 -2951 6060 -2899
rect 6076 -2951 6128 -2899
rect 6140 -2933 6192 -2899
rect 6204 -2933 6256 -2899
rect 6140 -2951 6165 -2933
rect 6165 -2951 6192 -2933
rect 6204 -2951 6237 -2933
rect 6237 -2951 6256 -2933
rect 6366 -2933 6418 -2899
rect 6430 -2933 6482 -2899
rect 6494 -2933 6546 -2899
rect 6366 -2951 6389 -2933
rect 6389 -2951 6418 -2933
rect 6430 -2951 6461 -2933
rect 6461 -2951 6482 -2933
rect 6494 -2951 6495 -2933
rect 6495 -2951 6546 -2933
rect 6562 -2951 6614 -2899
rect 6626 -2933 6678 -2899
rect 6690 -2933 6742 -2899
rect 6626 -2951 6647 -2933
rect 6647 -2951 6678 -2933
rect 6690 -2951 6719 -2933
rect 6719 -2951 6742 -2933
rect 7094 -2773 7146 -2721
rect 7158 -2773 7210 -2721
rect 7222 -2773 7274 -2721
rect 7290 -2773 7342 -2721
rect 7354 -2773 7406 -2721
rect 7418 -2773 7470 -2721
rect 7482 -2773 7534 -2721
rect 7550 -2773 7602 -2721
rect 7614 -2773 7666 -2721
rect 7678 -2773 7730 -2721
rect 8078 -2604 8101 -2583
rect 8101 -2604 8130 -2583
rect 8142 -2604 8173 -2583
rect 8173 -2604 8194 -2583
rect 8078 -2635 8130 -2604
rect 8142 -2635 8194 -2604
rect 8206 -2635 8258 -2583
rect 8274 -2604 8325 -2583
rect 8325 -2604 8326 -2583
rect 8338 -2604 8359 -2583
rect 8359 -2604 8390 -2583
rect 8402 -2604 8431 -2583
rect 8431 -2604 8454 -2583
rect 8274 -2635 8326 -2604
rect 8338 -2635 8390 -2604
rect 8402 -2635 8454 -2604
rect 8564 -2604 8583 -2583
rect 8583 -2604 8616 -2583
rect 8628 -2604 8655 -2583
rect 8655 -2604 8680 -2583
rect 8564 -2635 8616 -2604
rect 8628 -2635 8680 -2604
rect 8692 -2635 8744 -2583
rect 8760 -2635 8812 -2583
rect 8824 -2604 8841 -2583
rect 8841 -2604 8875 -2583
rect 8875 -2604 8876 -2583
rect 8824 -2635 8876 -2604
rect 8888 -2604 8913 -2583
rect 8913 -2604 8940 -2583
rect 8888 -2635 8940 -2604
rect 14940 -1754 14992 -1702
rect 15004 -1754 15056 -1702
rect 15068 -1754 15120 -1702
rect 14680 -2055 14732 -2003
rect 14744 -2055 14796 -2003
rect 14808 -2055 14860 -2003
rect 15457 -1754 15509 -1702
rect 15521 -1754 15573 -1702
rect 15585 -1754 15637 -1702
rect 15197 -2055 15249 -2003
rect 15261 -2055 15313 -2003
rect 15325 -2055 15377 -2003
rect 15650 -1894 15702 -1842
rect 15714 -1894 15766 -1842
rect 15778 -1894 15830 -1842
rect 16167 -1894 16219 -1842
rect 16231 -1894 16283 -1842
rect 16295 -1894 16347 -1842
rect 15908 -2199 15960 -2147
rect 15972 -2199 16024 -2147
rect 16036 -2199 16088 -2147
rect 16617 -1754 16669 -1702
rect 16681 -1754 16733 -1702
rect 16745 -1754 16797 -1702
rect 16425 -2199 16477 -2147
rect 16489 -2199 16541 -2147
rect 16553 -2199 16605 -2147
rect 17135 -1754 17187 -1702
rect 17199 -1754 17251 -1702
rect 17263 -1754 17315 -1702
rect 16874 -2055 16926 -2003
rect 16938 -2055 16990 -2003
rect 17002 -2055 17054 -2003
rect 17650 -1754 17702 -1702
rect 17714 -1754 17766 -1702
rect 17778 -1754 17830 -1702
rect 17392 -2055 17444 -2003
rect 17456 -2055 17508 -2003
rect 17520 -2055 17572 -2003
rect 10240 -2604 10267 -2583
rect 10267 -2604 10292 -2583
rect 10240 -2635 10292 -2604
rect 10304 -2604 10305 -2583
rect 10305 -2604 10339 -2583
rect 10339 -2604 10356 -2583
rect 10304 -2635 10356 -2604
rect 10368 -2635 10420 -2583
rect 10436 -2635 10488 -2583
rect 10500 -2604 10525 -2583
rect 10525 -2604 10552 -2583
rect 10564 -2604 10597 -2583
rect 10597 -2604 10616 -2583
rect 10500 -2635 10552 -2604
rect 10564 -2635 10616 -2604
rect 10726 -2604 10749 -2583
rect 10749 -2604 10778 -2583
rect 10790 -2604 10821 -2583
rect 10821 -2604 10842 -2583
rect 10854 -2604 10855 -2583
rect 10855 -2604 10906 -2583
rect 10726 -2635 10778 -2604
rect 10790 -2635 10842 -2604
rect 10854 -2635 10906 -2604
rect 10922 -2635 10974 -2583
rect 10986 -2604 11007 -2583
rect 11007 -2604 11038 -2583
rect 11050 -2604 11079 -2583
rect 11079 -2604 11102 -2583
rect 10986 -2635 11038 -2604
rect 11050 -2635 11102 -2604
rect 8078 -2773 8130 -2721
rect 8142 -2773 8194 -2721
rect 8206 -2773 8258 -2721
rect 8274 -2773 8326 -2721
rect 8338 -2773 8390 -2721
rect 8402 -2773 8454 -2721
rect 8564 -2773 8616 -2721
rect 8628 -2773 8680 -2721
rect 8692 -2773 8744 -2721
rect 8760 -2773 8812 -2721
rect 8824 -2773 8876 -2721
rect 8888 -2773 8940 -2721
rect 8078 -2933 8130 -2899
rect 8142 -2933 8194 -2899
rect 8078 -2951 8101 -2933
rect 8101 -2951 8130 -2933
rect 8142 -2951 8173 -2933
rect 8173 -2951 8194 -2933
rect 8206 -2951 8258 -2899
rect 8274 -2933 8326 -2899
rect 8338 -2933 8390 -2899
rect 8402 -2933 8454 -2899
rect 8274 -2951 8325 -2933
rect 8325 -2951 8326 -2933
rect 8338 -2951 8359 -2933
rect 8359 -2951 8390 -2933
rect 8402 -2951 8431 -2933
rect 8431 -2951 8454 -2933
rect 8564 -2933 8616 -2899
rect 8628 -2933 8680 -2899
rect 8564 -2951 8583 -2933
rect 8583 -2951 8616 -2933
rect 8628 -2951 8655 -2933
rect 8655 -2951 8680 -2933
rect 8692 -2951 8744 -2899
rect 8760 -2951 8812 -2899
rect 8824 -2933 8876 -2899
rect 8824 -2951 8841 -2933
rect 8841 -2951 8875 -2933
rect 8875 -2951 8876 -2933
rect 8888 -2933 8940 -2899
rect 8888 -2951 8913 -2933
rect 8913 -2951 8940 -2933
rect 1607 -3378 1659 -3326
rect 1671 -3378 1723 -3326
rect 1735 -3378 1787 -3326
rect 2125 -3378 2177 -3326
rect 2189 -3378 2241 -3326
rect 2253 -3378 2305 -3326
rect 2577 -3547 2629 -3495
rect 2641 -3547 2693 -3495
rect 2705 -3547 2757 -3495
rect 1348 -3709 1400 -3657
rect 1412 -3709 1464 -3657
rect 1476 -3709 1528 -3657
rect 1865 -3709 1917 -3657
rect 1929 -3709 1981 -3657
rect 1993 -3709 2045 -3657
rect 2382 -3709 2434 -3657
rect 2446 -3709 2498 -3657
rect 2510 -3709 2562 -3657
rect 3094 -3547 3146 -3495
rect 3158 -3547 3210 -3495
rect 3222 -3547 3274 -3495
rect 3802 -3378 3854 -3326
rect 3866 -3378 3918 -3326
rect 3930 -3378 3982 -3326
rect 4319 -3378 4371 -3326
rect 4383 -3378 4435 -3326
rect 4447 -3378 4499 -3326
rect 10240 -2773 10292 -2721
rect 10304 -2773 10356 -2721
rect 10368 -2773 10420 -2721
rect 10436 -2773 10488 -2721
rect 10500 -2773 10552 -2721
rect 10564 -2773 10616 -2721
rect 10726 -2773 10778 -2721
rect 10790 -2773 10842 -2721
rect 10854 -2773 10906 -2721
rect 10922 -2773 10974 -2721
rect 10986 -2773 11038 -2721
rect 11050 -2773 11102 -2721
rect 10240 -2933 10292 -2899
rect 10240 -2951 10267 -2933
rect 10267 -2951 10292 -2933
rect 10304 -2933 10356 -2899
rect 10304 -2951 10305 -2933
rect 10305 -2951 10339 -2933
rect 10339 -2951 10356 -2933
rect 10368 -2951 10420 -2899
rect 10436 -2951 10488 -2899
rect 10500 -2933 10552 -2899
rect 10564 -2933 10616 -2899
rect 10500 -2951 10525 -2933
rect 10525 -2951 10552 -2933
rect 10564 -2951 10597 -2933
rect 10597 -2951 10616 -2933
rect 10726 -2933 10778 -2899
rect 10790 -2933 10842 -2899
rect 10854 -2933 10906 -2899
rect 10726 -2951 10749 -2933
rect 10749 -2951 10778 -2933
rect 10790 -2951 10821 -2933
rect 10821 -2951 10842 -2933
rect 10854 -2951 10855 -2933
rect 10855 -2951 10906 -2933
rect 10922 -2951 10974 -2899
rect 10986 -2933 11038 -2899
rect 11050 -2933 11102 -2899
rect 10986 -2951 11007 -2933
rect 11007 -2951 11038 -2933
rect 11050 -2951 11079 -2933
rect 11079 -2951 11102 -2933
rect 11450 -2773 11502 -2721
rect 11514 -2773 11566 -2721
rect 11578 -2773 11630 -2721
rect 11646 -2773 11698 -2721
rect 11710 -2773 11762 -2721
rect 11774 -2773 11826 -2721
rect 11838 -2773 11890 -2721
rect 11906 -2773 11958 -2721
rect 11970 -2773 12022 -2721
rect 12034 -2773 12086 -2721
rect 12438 -2604 12461 -2583
rect 12461 -2604 12490 -2583
rect 12502 -2604 12533 -2583
rect 12533 -2604 12554 -2583
rect 12438 -2635 12490 -2604
rect 12502 -2635 12554 -2604
rect 12566 -2635 12618 -2583
rect 12634 -2604 12685 -2583
rect 12685 -2604 12686 -2583
rect 12698 -2604 12719 -2583
rect 12719 -2604 12750 -2583
rect 12762 -2604 12791 -2583
rect 12791 -2604 12814 -2583
rect 12634 -2635 12686 -2604
rect 12698 -2635 12750 -2604
rect 12762 -2635 12814 -2604
rect 12924 -2604 12943 -2583
rect 12943 -2604 12976 -2583
rect 12988 -2604 13015 -2583
rect 13015 -2604 13040 -2583
rect 12924 -2635 12976 -2604
rect 12988 -2635 13040 -2604
rect 13052 -2635 13104 -2583
rect 13120 -2635 13172 -2583
rect 13184 -2604 13201 -2583
rect 13201 -2604 13235 -2583
rect 13235 -2604 13236 -2583
rect 13184 -2635 13236 -2604
rect 13248 -2604 13273 -2583
rect 13273 -2604 13300 -2583
rect 13248 -2635 13300 -2604
rect 14597 -2604 14624 -2583
rect 14624 -2604 14649 -2583
rect 14597 -2635 14649 -2604
rect 14661 -2604 14662 -2583
rect 14662 -2604 14696 -2583
rect 14696 -2604 14713 -2583
rect 14661 -2635 14713 -2604
rect 14725 -2635 14777 -2583
rect 14793 -2635 14845 -2583
rect 14857 -2604 14882 -2583
rect 14882 -2604 14909 -2583
rect 14921 -2604 14954 -2583
rect 14954 -2604 14973 -2583
rect 14857 -2635 14909 -2604
rect 14921 -2635 14973 -2604
rect 15083 -2604 15106 -2583
rect 15106 -2604 15135 -2583
rect 15147 -2604 15178 -2583
rect 15178 -2604 15199 -2583
rect 15211 -2604 15212 -2583
rect 15212 -2604 15263 -2583
rect 15083 -2635 15135 -2604
rect 15147 -2635 15199 -2604
rect 15211 -2635 15263 -2604
rect 15279 -2635 15331 -2583
rect 15343 -2604 15364 -2583
rect 15364 -2604 15395 -2583
rect 15407 -2604 15436 -2583
rect 15436 -2604 15459 -2583
rect 15343 -2635 15395 -2604
rect 15407 -2635 15459 -2604
rect 12438 -2773 12490 -2721
rect 12502 -2773 12554 -2721
rect 12566 -2773 12618 -2721
rect 12634 -2773 12686 -2721
rect 12698 -2773 12750 -2721
rect 12762 -2773 12814 -2721
rect 12924 -2773 12976 -2721
rect 12988 -2773 13040 -2721
rect 13052 -2773 13104 -2721
rect 13120 -2773 13172 -2721
rect 13184 -2773 13236 -2721
rect 13248 -2773 13300 -2721
rect 12438 -2933 12490 -2899
rect 12502 -2933 12554 -2899
rect 12438 -2951 12461 -2933
rect 12461 -2951 12490 -2933
rect 12502 -2951 12533 -2933
rect 12533 -2951 12554 -2933
rect 12566 -2951 12618 -2899
rect 12634 -2933 12686 -2899
rect 12698 -2933 12750 -2899
rect 12762 -2933 12814 -2899
rect 12634 -2951 12685 -2933
rect 12685 -2951 12686 -2933
rect 12698 -2951 12719 -2933
rect 12719 -2951 12750 -2933
rect 12762 -2951 12791 -2933
rect 12791 -2951 12814 -2933
rect 12924 -2933 12976 -2899
rect 12988 -2933 13040 -2899
rect 12924 -2951 12943 -2933
rect 12943 -2951 12976 -2933
rect 12988 -2951 13015 -2933
rect 13015 -2951 13040 -2933
rect 13052 -2951 13104 -2899
rect 13120 -2951 13172 -2899
rect 13184 -2933 13236 -2899
rect 13184 -2951 13201 -2933
rect 13201 -2951 13235 -2933
rect 13235 -2951 13236 -2933
rect 13248 -2933 13300 -2899
rect 13248 -2951 13273 -2933
rect 13273 -2951 13300 -2933
rect 3543 -3709 3595 -3657
rect 3607 -3709 3659 -3657
rect 3671 -3709 3723 -3657
rect 4060 -3709 4112 -3657
rect 4124 -3709 4176 -3657
rect 4188 -3709 4240 -3657
rect 4575 -3709 4627 -3657
rect 4639 -3709 4691 -3657
rect 4703 -3709 4755 -3657
rect 5964 -3378 6016 -3326
rect 6028 -3378 6080 -3326
rect 6092 -3378 6144 -3326
rect 6481 -3378 6533 -3326
rect 6545 -3378 6597 -3326
rect 6609 -3378 6661 -3326
rect 5708 -3709 5760 -3657
rect 5772 -3709 5824 -3657
rect 5836 -3709 5888 -3657
rect 6223 -3709 6275 -3657
rect 6287 -3709 6339 -3657
rect 6351 -3709 6403 -3657
rect 6740 -3709 6792 -3657
rect 6804 -3709 6856 -3657
rect 6868 -3709 6920 -3657
rect 2834 -3878 2886 -3826
rect 2898 -3878 2950 -3826
rect 2962 -3878 3014 -3826
rect 3351 -3878 3403 -3826
rect 3415 -3878 3467 -3826
rect 3479 -3878 3531 -3826
rect 7189 -3547 7241 -3495
rect 7253 -3547 7305 -3495
rect 7317 -3547 7369 -3495
rect 7706 -3547 7758 -3495
rect 7770 -3547 7822 -3495
rect 7834 -3547 7886 -3495
rect 8158 -3378 8210 -3326
rect 8222 -3378 8274 -3326
rect 8286 -3378 8338 -3326
rect 8675 -3378 8727 -3326
rect 8739 -3378 8791 -3326
rect 8803 -3378 8855 -3326
rect 14597 -2773 14649 -2721
rect 14661 -2773 14713 -2721
rect 14725 -2773 14777 -2721
rect 14793 -2773 14845 -2721
rect 14857 -2773 14909 -2721
rect 14921 -2773 14973 -2721
rect 15083 -2773 15135 -2721
rect 15147 -2773 15199 -2721
rect 15211 -2773 15263 -2721
rect 15279 -2773 15331 -2721
rect 15343 -2773 15395 -2721
rect 15407 -2773 15459 -2721
rect 14597 -2933 14649 -2899
rect 14597 -2951 14624 -2933
rect 14624 -2951 14649 -2933
rect 14661 -2933 14713 -2899
rect 14661 -2951 14662 -2933
rect 14662 -2951 14696 -2933
rect 14696 -2951 14713 -2933
rect 14725 -2951 14777 -2899
rect 14793 -2951 14845 -2899
rect 14857 -2933 14909 -2899
rect 14921 -2933 14973 -2899
rect 14857 -2951 14882 -2933
rect 14882 -2951 14909 -2933
rect 14921 -2951 14954 -2933
rect 14954 -2951 14973 -2933
rect 15083 -2933 15135 -2899
rect 15147 -2933 15199 -2899
rect 15211 -2933 15263 -2899
rect 15083 -2951 15106 -2933
rect 15106 -2951 15135 -2933
rect 15147 -2951 15178 -2933
rect 15178 -2951 15199 -2933
rect 15211 -2951 15212 -2933
rect 15212 -2951 15263 -2933
rect 15279 -2951 15331 -2899
rect 15343 -2933 15395 -2899
rect 15407 -2933 15459 -2899
rect 15343 -2951 15364 -2933
rect 15364 -2951 15395 -2933
rect 15407 -2951 15436 -2933
rect 15436 -2951 15459 -2933
rect 15811 -2773 15863 -2721
rect 15875 -2773 15927 -2721
rect 15939 -2773 15991 -2721
rect 16007 -2773 16059 -2721
rect 16071 -2773 16123 -2721
rect 16135 -2773 16187 -2721
rect 16199 -2773 16251 -2721
rect 16267 -2773 16319 -2721
rect 16331 -2773 16383 -2721
rect 16395 -2773 16447 -2721
rect 16795 -2604 16818 -2583
rect 16818 -2604 16847 -2583
rect 16859 -2604 16890 -2583
rect 16890 -2604 16911 -2583
rect 16795 -2635 16847 -2604
rect 16859 -2635 16911 -2604
rect 16923 -2635 16975 -2583
rect 16991 -2604 17042 -2583
rect 17042 -2604 17043 -2583
rect 17055 -2604 17076 -2583
rect 17076 -2604 17107 -2583
rect 17119 -2604 17148 -2583
rect 17148 -2604 17171 -2583
rect 16991 -2635 17043 -2604
rect 17055 -2635 17107 -2604
rect 17119 -2635 17171 -2604
rect 17281 -2604 17300 -2583
rect 17300 -2604 17333 -2583
rect 17345 -2604 17372 -2583
rect 17372 -2604 17397 -2583
rect 17281 -2635 17333 -2604
rect 17345 -2635 17397 -2604
rect 17409 -2635 17461 -2583
rect 17477 -2635 17529 -2583
rect 17541 -2604 17558 -2583
rect 17558 -2604 17592 -2583
rect 17592 -2604 17593 -2583
rect 17541 -2635 17593 -2604
rect 17605 -2604 17630 -2583
rect 17630 -2604 17657 -2583
rect 17605 -2635 17657 -2604
rect 16795 -2773 16847 -2721
rect 16859 -2773 16911 -2721
rect 16923 -2773 16975 -2721
rect 16991 -2773 17043 -2721
rect 17055 -2773 17107 -2721
rect 17119 -2773 17171 -2721
rect 17281 -2773 17333 -2721
rect 17345 -2773 17397 -2721
rect 17409 -2773 17461 -2721
rect 17477 -2773 17529 -2721
rect 17541 -2773 17593 -2721
rect 17605 -2773 17657 -2721
rect 16795 -2933 16847 -2899
rect 16859 -2933 16911 -2899
rect 16795 -2951 16818 -2933
rect 16818 -2951 16847 -2933
rect 16859 -2951 16890 -2933
rect 16890 -2951 16911 -2933
rect 16923 -2951 16975 -2899
rect 16991 -2933 17043 -2899
rect 17055 -2933 17107 -2899
rect 17119 -2933 17171 -2899
rect 16991 -2951 17042 -2933
rect 17042 -2951 17043 -2933
rect 17055 -2951 17076 -2933
rect 17076 -2951 17107 -2933
rect 17119 -2951 17148 -2933
rect 17148 -2951 17171 -2933
rect 17281 -2933 17333 -2899
rect 17345 -2933 17397 -2899
rect 17281 -2951 17300 -2933
rect 17300 -2951 17333 -2933
rect 17345 -2951 17372 -2933
rect 17372 -2951 17397 -2933
rect 17409 -2951 17461 -2899
rect 17477 -2951 17529 -2899
rect 17541 -2933 17593 -2899
rect 17541 -2951 17558 -2933
rect 17558 -2951 17592 -2933
rect 17592 -2951 17593 -2933
rect 17605 -2933 17657 -2899
rect 17605 -2951 17630 -2933
rect 17630 -2951 17657 -2933
rect 7901 -3709 7953 -3657
rect 7965 -3709 8017 -3657
rect 8029 -3709 8081 -3657
rect 8417 -3709 8469 -3657
rect 8481 -3709 8533 -3657
rect 8545 -3709 8597 -3657
rect 8935 -3709 8987 -3657
rect 8999 -3709 9051 -3657
rect 9063 -3709 9115 -3657
rect 10325 -3378 10377 -3326
rect 10389 -3378 10441 -3326
rect 10453 -3378 10505 -3326
rect 10842 -3378 10894 -3326
rect 10906 -3378 10958 -3326
rect 10970 -3378 11022 -3326
rect 11294 -3547 11346 -3495
rect 11358 -3547 11410 -3495
rect 11422 -3547 11474 -3495
rect 10065 -3709 10117 -3657
rect 10129 -3709 10181 -3657
rect 10193 -3709 10245 -3657
rect 10583 -3709 10635 -3657
rect 10647 -3709 10699 -3657
rect 10711 -3709 10763 -3657
rect 11099 -3709 11151 -3657
rect 11163 -3709 11215 -3657
rect 11227 -3709 11279 -3657
rect 6931 -3878 6983 -3826
rect 6995 -3878 7047 -3826
rect 7059 -3878 7111 -3826
rect 7449 -3878 7501 -3826
rect 7513 -3878 7565 -3826
rect 7577 -3878 7629 -3826
rect 11811 -3547 11863 -3495
rect 11875 -3547 11927 -3495
rect 11939 -3547 11991 -3495
rect 12519 -3378 12571 -3326
rect 12583 -3378 12635 -3326
rect 12647 -3378 12699 -3326
rect 13036 -3378 13088 -3326
rect 13100 -3378 13152 -3326
rect 13164 -3378 13216 -3326
rect 12260 -3709 12312 -3657
rect 12324 -3709 12376 -3657
rect 12388 -3709 12440 -3657
rect 12777 -3709 12829 -3657
rect 12841 -3709 12893 -3657
rect 12905 -3709 12957 -3657
rect 13292 -3709 13344 -3657
rect 13356 -3709 13408 -3657
rect 13420 -3709 13472 -3657
rect 14681 -3378 14733 -3326
rect 14745 -3378 14797 -3326
rect 14809 -3378 14861 -3326
rect 15198 -3378 15250 -3326
rect 15262 -3378 15314 -3326
rect 15326 -3378 15378 -3326
rect 14425 -3709 14477 -3657
rect 14489 -3709 14541 -3657
rect 14553 -3709 14605 -3657
rect 14940 -3709 14992 -3657
rect 15004 -3709 15056 -3657
rect 15068 -3709 15120 -3657
rect 15457 -3709 15509 -3657
rect 15521 -3709 15573 -3657
rect 15585 -3709 15637 -3657
rect 11551 -3878 11603 -3826
rect 11615 -3878 11667 -3826
rect 11679 -3878 11731 -3826
rect 12069 -3878 12121 -3826
rect 12133 -3878 12185 -3826
rect 12197 -3878 12249 -3826
rect 15906 -3547 15958 -3495
rect 15970 -3547 16022 -3495
rect 16034 -3547 16086 -3495
rect 16423 -3547 16475 -3495
rect 16487 -3547 16539 -3495
rect 16551 -3547 16603 -3495
rect 16875 -3378 16927 -3326
rect 16939 -3378 16991 -3326
rect 17003 -3378 17055 -3326
rect 17393 -3378 17445 -3326
rect 17457 -3378 17509 -3326
rect 17521 -3378 17573 -3326
rect 16618 -3709 16670 -3657
rect 16682 -3709 16734 -3657
rect 16746 -3709 16798 -3657
rect 17135 -3709 17187 -3657
rect 17199 -3709 17251 -3657
rect 17263 -3709 17315 -3657
rect 17652 -3709 17704 -3657
rect 17716 -3709 17768 -3657
rect 17780 -3709 17832 -3657
rect 15649 -3878 15701 -3826
rect 15713 -3878 15765 -3826
rect 15777 -3878 15829 -3826
rect 16166 -3878 16218 -3826
rect 16230 -3878 16282 -3826
rect 16294 -3878 16346 -3826
rect 2834 -4937 2886 -4885
rect 2898 -4937 2950 -4885
rect 2962 -4937 3014 -4885
rect 3351 -4937 3403 -4885
rect 3415 -4937 3467 -4885
rect 3479 -4937 3531 -4885
rect 1348 -5106 1400 -5054
rect 1412 -5106 1464 -5054
rect 1476 -5106 1528 -5054
rect 1865 -5106 1917 -5054
rect 1929 -5106 1981 -5054
rect 1993 -5106 2045 -5054
rect 2382 -5106 2434 -5054
rect 2446 -5106 2498 -5054
rect 2510 -5106 2562 -5054
rect 1607 -5438 1659 -5386
rect 1671 -5438 1723 -5386
rect 1735 -5438 1787 -5386
rect 2125 -5438 2177 -5386
rect 2189 -5438 2241 -5386
rect 2253 -5438 2305 -5386
rect 2577 -5269 2629 -5217
rect 2641 -5269 2693 -5217
rect 2705 -5269 2757 -5217
rect 3094 -5269 3146 -5217
rect 3158 -5269 3210 -5217
rect 3222 -5269 3274 -5217
rect 6931 -4937 6983 -4885
rect 6995 -4937 7047 -4885
rect 7059 -4937 7111 -4885
rect 7449 -4937 7501 -4885
rect 7513 -4937 7565 -4885
rect 7577 -4937 7629 -4885
rect 3543 -5106 3595 -5054
rect 3607 -5106 3659 -5054
rect 3671 -5106 3723 -5054
rect 4060 -5106 4112 -5054
rect 4124 -5106 4176 -5054
rect 4188 -5106 4240 -5054
rect 4575 -5106 4627 -5054
rect 4639 -5106 4691 -5054
rect 4703 -5106 4755 -5054
rect 3802 -5438 3854 -5386
rect 3866 -5438 3918 -5386
rect 3930 -5438 3982 -5386
rect 4319 -5438 4371 -5386
rect 4383 -5438 4435 -5386
rect 4447 -5438 4499 -5386
rect 5708 -5106 5760 -5054
rect 5772 -5106 5824 -5054
rect 5836 -5106 5888 -5054
rect 6223 -5106 6275 -5054
rect 6287 -5106 6339 -5054
rect 6351 -5106 6403 -5054
rect 6740 -5106 6792 -5054
rect 6804 -5106 6856 -5054
rect 6868 -5106 6920 -5054
rect 5964 -5438 6016 -5386
rect 6028 -5438 6080 -5386
rect 6092 -5438 6144 -5386
rect 6481 -5438 6533 -5386
rect 6545 -5438 6597 -5386
rect 6609 -5438 6661 -5386
rect 7189 -5269 7241 -5217
rect 7253 -5269 7305 -5217
rect 7317 -5269 7369 -5217
rect 11551 -4937 11603 -4885
rect 11615 -4937 11667 -4885
rect 11679 -4937 11731 -4885
rect 12069 -4937 12121 -4885
rect 12133 -4937 12185 -4885
rect 12197 -4937 12249 -4885
rect 7901 -5106 7953 -5054
rect 7965 -5106 8017 -5054
rect 8029 -5106 8081 -5054
rect 8417 -5106 8469 -5054
rect 8481 -5106 8533 -5054
rect 8545 -5106 8597 -5054
rect 8935 -5106 8987 -5054
rect 8999 -5106 9051 -5054
rect 9063 -5106 9115 -5054
rect 7706 -5269 7758 -5217
rect 7770 -5269 7822 -5217
rect 7834 -5269 7886 -5217
rect 8158 -5438 8210 -5386
rect 8222 -5438 8274 -5386
rect 8286 -5438 8338 -5386
rect 8675 -5438 8727 -5386
rect 8739 -5438 8791 -5386
rect 8803 -5438 8855 -5386
rect 10065 -5106 10117 -5054
rect 10129 -5106 10181 -5054
rect 10193 -5106 10245 -5054
rect 10583 -5106 10635 -5054
rect 10647 -5106 10699 -5054
rect 10711 -5106 10763 -5054
rect 11099 -5106 11151 -5054
rect 11163 -5106 11215 -5054
rect 11227 -5106 11279 -5054
rect 1523 -5831 1550 -5812
rect 1550 -5831 1575 -5812
rect 1523 -5864 1575 -5831
rect 1587 -5831 1588 -5812
rect 1588 -5831 1622 -5812
rect 1622 -5831 1639 -5812
rect 1587 -5864 1639 -5831
rect 1651 -5864 1703 -5812
rect 1719 -5864 1771 -5812
rect 1783 -5831 1808 -5812
rect 1808 -5831 1835 -5812
rect 1847 -5831 1880 -5812
rect 1880 -5831 1899 -5812
rect 1783 -5864 1835 -5831
rect 1847 -5864 1899 -5831
rect 2009 -5831 2032 -5812
rect 2032 -5831 2061 -5812
rect 2073 -5831 2104 -5812
rect 2104 -5831 2125 -5812
rect 2137 -5831 2138 -5812
rect 2138 -5831 2189 -5812
rect 2009 -5864 2061 -5831
rect 2073 -5864 2125 -5831
rect 2137 -5864 2189 -5831
rect 2205 -5864 2257 -5812
rect 2269 -5831 2290 -5812
rect 2290 -5831 2321 -5812
rect 2333 -5831 2362 -5812
rect 2362 -5831 2385 -5812
rect 2269 -5864 2321 -5831
rect 2333 -5864 2385 -5831
rect 1523 -6042 1575 -5990
rect 1587 -6042 1639 -5990
rect 1651 -6042 1703 -5990
rect 1719 -6042 1771 -5990
rect 1783 -6042 1835 -5990
rect 1847 -6042 1899 -5990
rect 2009 -6042 2061 -5990
rect 2073 -6042 2125 -5990
rect 2137 -6042 2189 -5990
rect 2205 -6042 2257 -5990
rect 2269 -6042 2321 -5990
rect 2333 -6042 2385 -5990
rect 1523 -6159 1575 -6129
rect 1523 -6181 1550 -6159
rect 1550 -6181 1575 -6159
rect 1587 -6159 1639 -6129
rect 1587 -6181 1588 -6159
rect 1588 -6181 1622 -6159
rect 1622 -6181 1639 -6159
rect 1651 -6181 1703 -6129
rect 1719 -6181 1771 -6129
rect 1783 -6159 1835 -6129
rect 1847 -6159 1899 -6129
rect 1783 -6181 1808 -6159
rect 1808 -6181 1835 -6159
rect 1847 -6181 1880 -6159
rect 1880 -6181 1899 -6159
rect 2009 -6159 2061 -6129
rect 2073 -6159 2125 -6129
rect 2137 -6159 2189 -6129
rect 2009 -6181 2032 -6159
rect 2032 -6181 2061 -6159
rect 2073 -6181 2104 -6159
rect 2104 -6181 2125 -6159
rect 2137 -6181 2138 -6159
rect 2138 -6181 2189 -6159
rect 2205 -6181 2257 -6129
rect 2269 -6159 2321 -6129
rect 2333 -6159 2385 -6129
rect 2269 -6181 2290 -6159
rect 2290 -6181 2321 -6159
rect 2333 -6181 2362 -6159
rect 2362 -6181 2385 -6159
rect 2733 -6042 2785 -5990
rect 2797 -6042 2849 -5990
rect 2861 -6042 2913 -5990
rect 2929 -6042 2981 -5990
rect 2993 -6042 3045 -5990
rect 3057 -6042 3109 -5990
rect 3121 -6042 3173 -5990
rect 3189 -6042 3241 -5990
rect 3253 -6042 3305 -5990
rect 3317 -6042 3369 -5990
rect 3721 -5831 3744 -5812
rect 3744 -5831 3773 -5812
rect 3785 -5831 3816 -5812
rect 3816 -5831 3837 -5812
rect 3721 -5864 3773 -5831
rect 3785 -5864 3837 -5831
rect 3849 -5864 3901 -5812
rect 3917 -5831 3968 -5812
rect 3968 -5831 3969 -5812
rect 3981 -5831 4002 -5812
rect 4002 -5831 4033 -5812
rect 4045 -5831 4074 -5812
rect 4074 -5831 4097 -5812
rect 3917 -5864 3969 -5831
rect 3981 -5864 4033 -5831
rect 4045 -5864 4097 -5831
rect 4207 -5831 4226 -5812
rect 4226 -5831 4259 -5812
rect 4271 -5831 4298 -5812
rect 4298 -5831 4323 -5812
rect 4207 -5864 4259 -5831
rect 4271 -5864 4323 -5831
rect 4335 -5864 4387 -5812
rect 4403 -5864 4455 -5812
rect 4467 -5831 4484 -5812
rect 4484 -5831 4518 -5812
rect 4518 -5831 4519 -5812
rect 4467 -5864 4519 -5831
rect 4531 -5831 4556 -5812
rect 4556 -5831 4583 -5812
rect 4531 -5864 4583 -5831
rect 3721 -6042 3773 -5990
rect 3785 -6042 3837 -5990
rect 3849 -6042 3901 -5990
rect 3917 -6042 3969 -5990
rect 3981 -6042 4033 -5990
rect 4045 -6042 4097 -5990
rect 4207 -6042 4259 -5990
rect 4271 -6042 4323 -5990
rect 4335 -6042 4387 -5990
rect 4403 -6042 4455 -5990
rect 4467 -6042 4519 -5990
rect 4531 -6042 4583 -5990
rect 10325 -5438 10377 -5386
rect 10389 -5438 10441 -5386
rect 10453 -5438 10505 -5386
rect 10842 -5438 10894 -5386
rect 10906 -5438 10958 -5386
rect 10970 -5438 11022 -5386
rect 11294 -5269 11346 -5217
rect 11358 -5269 11410 -5217
rect 11422 -5269 11474 -5217
rect 11811 -5269 11863 -5217
rect 11875 -5269 11927 -5217
rect 11939 -5269 11991 -5217
rect 15649 -4937 15701 -4885
rect 15713 -4937 15765 -4885
rect 15777 -4937 15829 -4885
rect 16166 -4937 16218 -4885
rect 16230 -4937 16282 -4885
rect 16294 -4937 16346 -4885
rect 12260 -5106 12312 -5054
rect 12324 -5106 12376 -5054
rect 12388 -5106 12440 -5054
rect 12777 -5106 12829 -5054
rect 12841 -5106 12893 -5054
rect 12905 -5106 12957 -5054
rect 13292 -5106 13344 -5054
rect 13356 -5106 13408 -5054
rect 13420 -5106 13472 -5054
rect 12519 -5438 12571 -5386
rect 12583 -5438 12635 -5386
rect 12647 -5438 12699 -5386
rect 13036 -5438 13088 -5386
rect 13100 -5438 13152 -5386
rect 13164 -5438 13216 -5386
rect 14425 -5106 14477 -5054
rect 14489 -5106 14541 -5054
rect 14553 -5106 14605 -5054
rect 14940 -5106 14992 -5054
rect 15004 -5106 15056 -5054
rect 15068 -5106 15120 -5054
rect 15457 -5106 15509 -5054
rect 15521 -5106 15573 -5054
rect 15585 -5106 15637 -5054
rect 5880 -5831 5907 -5812
rect 5907 -5831 5932 -5812
rect 5880 -5864 5932 -5831
rect 5944 -5831 5945 -5812
rect 5945 -5831 5979 -5812
rect 5979 -5831 5996 -5812
rect 5944 -5864 5996 -5831
rect 6008 -5864 6060 -5812
rect 6076 -5864 6128 -5812
rect 6140 -5831 6165 -5812
rect 6165 -5831 6192 -5812
rect 6204 -5831 6237 -5812
rect 6237 -5831 6256 -5812
rect 6140 -5864 6192 -5831
rect 6204 -5864 6256 -5831
rect 6366 -5831 6389 -5812
rect 6389 -5831 6418 -5812
rect 6430 -5831 6461 -5812
rect 6461 -5831 6482 -5812
rect 6494 -5831 6495 -5812
rect 6495 -5831 6546 -5812
rect 6366 -5864 6418 -5831
rect 6430 -5864 6482 -5831
rect 6494 -5864 6546 -5831
rect 6562 -5864 6614 -5812
rect 6626 -5831 6647 -5812
rect 6647 -5831 6678 -5812
rect 6690 -5831 6719 -5812
rect 6719 -5831 6742 -5812
rect 6626 -5864 6678 -5831
rect 6690 -5864 6742 -5831
rect 5880 -6042 5932 -5990
rect 5944 -6042 5996 -5990
rect 6008 -6042 6060 -5990
rect 6076 -6042 6128 -5990
rect 6140 -6042 6192 -5990
rect 6204 -6042 6256 -5990
rect 6366 -6042 6418 -5990
rect 6430 -6042 6482 -5990
rect 6494 -6042 6546 -5990
rect 6562 -6042 6614 -5990
rect 6626 -6042 6678 -5990
rect 6690 -6042 6742 -5990
rect 3721 -6159 3773 -6129
rect 3785 -6159 3837 -6129
rect 3721 -6181 3744 -6159
rect 3744 -6181 3773 -6159
rect 3785 -6181 3816 -6159
rect 3816 -6181 3837 -6159
rect 3849 -6181 3901 -6129
rect 3917 -6159 3969 -6129
rect 3981 -6159 4033 -6129
rect 4045 -6159 4097 -6129
rect 3917 -6181 3968 -6159
rect 3968 -6181 3969 -6159
rect 3981 -6181 4002 -6159
rect 4002 -6181 4033 -6159
rect 4045 -6181 4074 -6159
rect 4074 -6181 4097 -6159
rect 4207 -6159 4259 -6129
rect 4271 -6159 4323 -6129
rect 4207 -6181 4226 -6159
rect 4226 -6181 4259 -6159
rect 4271 -6181 4298 -6159
rect 4298 -6181 4323 -6159
rect 4335 -6181 4387 -6129
rect 4403 -6181 4455 -6129
rect 4467 -6159 4519 -6129
rect 4467 -6181 4484 -6159
rect 4484 -6181 4518 -6159
rect 4518 -6181 4519 -6159
rect 4531 -6159 4583 -6129
rect 4531 -6181 4556 -6159
rect 4556 -6181 4583 -6159
rect 5880 -6159 5932 -6129
rect 5880 -6181 5907 -6159
rect 5907 -6181 5932 -6159
rect 5944 -6159 5996 -6129
rect 5944 -6181 5945 -6159
rect 5945 -6181 5979 -6159
rect 5979 -6181 5996 -6159
rect 6008 -6181 6060 -6129
rect 6076 -6181 6128 -6129
rect 6140 -6159 6192 -6129
rect 6204 -6159 6256 -6129
rect 6140 -6181 6165 -6159
rect 6165 -6181 6192 -6159
rect 6204 -6181 6237 -6159
rect 6237 -6181 6256 -6159
rect 6366 -6159 6418 -6129
rect 6430 -6159 6482 -6129
rect 6494 -6159 6546 -6129
rect 6366 -6181 6389 -6159
rect 6389 -6181 6418 -6159
rect 6430 -6181 6461 -6159
rect 6461 -6181 6482 -6159
rect 6494 -6181 6495 -6159
rect 6495 -6181 6546 -6159
rect 6562 -6181 6614 -6129
rect 6626 -6159 6678 -6129
rect 6690 -6159 6742 -6129
rect 6626 -6181 6647 -6159
rect 6647 -6181 6678 -6159
rect 6690 -6181 6719 -6159
rect 6719 -6181 6742 -6159
rect 7094 -6042 7146 -5990
rect 7158 -6042 7210 -5990
rect 7222 -6042 7274 -5990
rect 7290 -6042 7342 -5990
rect 7354 -6042 7406 -5990
rect 7418 -6042 7470 -5990
rect 7482 -6042 7534 -5990
rect 7550 -6042 7602 -5990
rect 7614 -6042 7666 -5990
rect 7678 -6042 7730 -5990
rect 8078 -5831 8101 -5812
rect 8101 -5831 8130 -5812
rect 8142 -5831 8173 -5812
rect 8173 -5831 8194 -5812
rect 8078 -5864 8130 -5831
rect 8142 -5864 8194 -5831
rect 8206 -5864 8258 -5812
rect 8274 -5831 8325 -5812
rect 8325 -5831 8326 -5812
rect 8338 -5831 8359 -5812
rect 8359 -5831 8390 -5812
rect 8402 -5831 8431 -5812
rect 8431 -5831 8454 -5812
rect 8274 -5864 8326 -5831
rect 8338 -5864 8390 -5831
rect 8402 -5864 8454 -5831
rect 8564 -5831 8583 -5812
rect 8583 -5831 8616 -5812
rect 8628 -5831 8655 -5812
rect 8655 -5831 8680 -5812
rect 8564 -5864 8616 -5831
rect 8628 -5864 8680 -5831
rect 8692 -5864 8744 -5812
rect 8760 -5864 8812 -5812
rect 8824 -5831 8841 -5812
rect 8841 -5831 8875 -5812
rect 8875 -5831 8876 -5812
rect 8824 -5864 8876 -5831
rect 8888 -5831 8913 -5812
rect 8913 -5831 8940 -5812
rect 8888 -5864 8940 -5831
rect 8078 -6042 8130 -5990
rect 8142 -6042 8194 -5990
rect 8206 -6042 8258 -5990
rect 8274 -6042 8326 -5990
rect 8338 -6042 8390 -5990
rect 8402 -6042 8454 -5990
rect 8564 -6042 8616 -5990
rect 8628 -6042 8680 -5990
rect 8692 -6042 8744 -5990
rect 8760 -6042 8812 -5990
rect 8824 -6042 8876 -5990
rect 8888 -6042 8940 -5990
rect 14681 -5438 14733 -5386
rect 14745 -5438 14797 -5386
rect 14809 -5438 14861 -5386
rect 15198 -5438 15250 -5386
rect 15262 -5438 15314 -5386
rect 15326 -5438 15378 -5386
rect 15906 -5269 15958 -5217
rect 15970 -5269 16022 -5217
rect 16034 -5269 16086 -5217
rect 16618 -5106 16670 -5054
rect 16682 -5106 16734 -5054
rect 16746 -5106 16798 -5054
rect 17135 -5106 17187 -5054
rect 17199 -5106 17251 -5054
rect 17263 -5106 17315 -5054
rect 17652 -5106 17704 -5054
rect 17716 -5106 17768 -5054
rect 17780 -5106 17832 -5054
rect 16423 -5269 16475 -5217
rect 16487 -5269 16539 -5217
rect 16551 -5269 16603 -5217
rect 16875 -5438 16927 -5386
rect 16939 -5438 16991 -5386
rect 17003 -5438 17055 -5386
rect 17393 -5438 17445 -5386
rect 17457 -5438 17509 -5386
rect 17521 -5438 17573 -5386
rect 10240 -5831 10267 -5812
rect 10267 -5831 10292 -5812
rect 10240 -5864 10292 -5831
rect 10304 -5831 10305 -5812
rect 10305 -5831 10339 -5812
rect 10339 -5831 10356 -5812
rect 10304 -5864 10356 -5831
rect 10368 -5864 10420 -5812
rect 10436 -5864 10488 -5812
rect 10500 -5831 10525 -5812
rect 10525 -5831 10552 -5812
rect 10564 -5831 10597 -5812
rect 10597 -5831 10616 -5812
rect 10500 -5864 10552 -5831
rect 10564 -5864 10616 -5831
rect 10726 -5831 10749 -5812
rect 10749 -5831 10778 -5812
rect 10790 -5831 10821 -5812
rect 10821 -5831 10842 -5812
rect 10854 -5831 10855 -5812
rect 10855 -5831 10906 -5812
rect 10726 -5864 10778 -5831
rect 10790 -5864 10842 -5831
rect 10854 -5864 10906 -5831
rect 10922 -5864 10974 -5812
rect 10986 -5831 11007 -5812
rect 11007 -5831 11038 -5812
rect 11050 -5831 11079 -5812
rect 11079 -5831 11102 -5812
rect 10986 -5864 11038 -5831
rect 11050 -5864 11102 -5831
rect 10240 -6042 10292 -5990
rect 10304 -6042 10356 -5990
rect 10368 -6042 10420 -5990
rect 10436 -6042 10488 -5990
rect 10500 -6042 10552 -5990
rect 10564 -6042 10616 -5990
rect 10726 -6042 10778 -5990
rect 10790 -6042 10842 -5990
rect 10854 -6042 10906 -5990
rect 10922 -6042 10974 -5990
rect 10986 -6042 11038 -5990
rect 11050 -6042 11102 -5990
rect 8078 -6159 8130 -6129
rect 8142 -6159 8194 -6129
rect 8078 -6181 8101 -6159
rect 8101 -6181 8130 -6159
rect 8142 -6181 8173 -6159
rect 8173 -6181 8194 -6159
rect 8206 -6181 8258 -6129
rect 8274 -6159 8326 -6129
rect 8338 -6159 8390 -6129
rect 8402 -6159 8454 -6129
rect 8274 -6181 8325 -6159
rect 8325 -6181 8326 -6159
rect 8338 -6181 8359 -6159
rect 8359 -6181 8390 -6159
rect 8402 -6181 8431 -6159
rect 8431 -6181 8454 -6159
rect 8564 -6159 8616 -6129
rect 8628 -6159 8680 -6129
rect 8564 -6181 8583 -6159
rect 8583 -6181 8616 -6159
rect 8628 -6181 8655 -6159
rect 8655 -6181 8680 -6159
rect 8692 -6181 8744 -6129
rect 8760 -6181 8812 -6129
rect 8824 -6159 8876 -6129
rect 8824 -6181 8841 -6159
rect 8841 -6181 8875 -6159
rect 8875 -6181 8876 -6159
rect 8888 -6159 8940 -6129
rect 8888 -6181 8913 -6159
rect 8913 -6181 8940 -6159
rect 1608 -6761 1660 -6709
rect 1672 -6761 1724 -6709
rect 1736 -6761 1788 -6709
rect 1350 -7062 1402 -7010
rect 1414 -7062 1466 -7010
rect 1478 -7062 1530 -7010
rect 2126 -6761 2178 -6709
rect 2190 -6761 2242 -6709
rect 2254 -6761 2306 -6709
rect 1865 -7062 1917 -7010
rect 1929 -7062 1981 -7010
rect 1993 -7062 2045 -7010
rect 2575 -6616 2627 -6564
rect 2639 -6616 2691 -6564
rect 2703 -6616 2755 -6564
rect 2383 -7062 2435 -7010
rect 2447 -7062 2499 -7010
rect 2511 -7062 2563 -7010
rect 3092 -6616 3144 -6564
rect 3156 -6616 3208 -6564
rect 3220 -6616 3272 -6564
rect 2833 -6922 2885 -6870
rect 2897 -6922 2949 -6870
rect 2961 -6922 3013 -6870
rect 3350 -6922 3402 -6870
rect 3414 -6922 3466 -6870
rect 3478 -6922 3530 -6870
rect 3803 -6761 3855 -6709
rect 3867 -6761 3919 -6709
rect 3931 -6761 3983 -6709
rect 3543 -7062 3595 -7010
rect 3607 -7062 3659 -7010
rect 3671 -7062 3723 -7010
rect 4320 -6761 4372 -6709
rect 4384 -6761 4436 -6709
rect 4448 -6761 4500 -6709
rect 4060 -7062 4112 -7010
rect 4124 -7062 4176 -7010
rect 4188 -7062 4240 -7010
rect 10240 -6159 10292 -6129
rect 10240 -6181 10267 -6159
rect 10267 -6181 10292 -6159
rect 10304 -6159 10356 -6129
rect 10304 -6181 10305 -6159
rect 10305 -6181 10339 -6159
rect 10339 -6181 10356 -6159
rect 10368 -6181 10420 -6129
rect 10436 -6181 10488 -6129
rect 10500 -6159 10552 -6129
rect 10564 -6159 10616 -6129
rect 10500 -6181 10525 -6159
rect 10525 -6181 10552 -6159
rect 10564 -6181 10597 -6159
rect 10597 -6181 10616 -6159
rect 10726 -6159 10778 -6129
rect 10790 -6159 10842 -6129
rect 10854 -6159 10906 -6129
rect 10726 -6181 10749 -6159
rect 10749 -6181 10778 -6159
rect 10790 -6181 10821 -6159
rect 10821 -6181 10842 -6159
rect 10854 -6181 10855 -6159
rect 10855 -6181 10906 -6159
rect 10922 -6181 10974 -6129
rect 10986 -6159 11038 -6129
rect 11050 -6159 11102 -6129
rect 10986 -6181 11007 -6159
rect 11007 -6181 11038 -6159
rect 11050 -6181 11079 -6159
rect 11079 -6181 11102 -6159
rect 11450 -6042 11502 -5990
rect 11514 -6042 11566 -5990
rect 11578 -6042 11630 -5990
rect 11646 -6042 11698 -5990
rect 11710 -6042 11762 -5990
rect 11774 -6042 11826 -5990
rect 11838 -6042 11890 -5990
rect 11906 -6042 11958 -5990
rect 11970 -6042 12022 -5990
rect 12034 -6042 12086 -5990
rect 12438 -5831 12461 -5812
rect 12461 -5831 12490 -5812
rect 12502 -5831 12533 -5812
rect 12533 -5831 12554 -5812
rect 12438 -5864 12490 -5831
rect 12502 -5864 12554 -5831
rect 12566 -5864 12618 -5812
rect 12634 -5831 12685 -5812
rect 12685 -5831 12686 -5812
rect 12698 -5831 12719 -5812
rect 12719 -5831 12750 -5812
rect 12762 -5831 12791 -5812
rect 12791 -5831 12814 -5812
rect 12634 -5864 12686 -5831
rect 12698 -5864 12750 -5831
rect 12762 -5864 12814 -5831
rect 12924 -5831 12943 -5812
rect 12943 -5831 12976 -5812
rect 12988 -5831 13015 -5812
rect 13015 -5831 13040 -5812
rect 12924 -5864 12976 -5831
rect 12988 -5864 13040 -5831
rect 13052 -5864 13104 -5812
rect 13120 -5864 13172 -5812
rect 13184 -5831 13201 -5812
rect 13201 -5831 13235 -5812
rect 13235 -5831 13236 -5812
rect 13184 -5864 13236 -5831
rect 13248 -5831 13273 -5812
rect 13273 -5831 13300 -5812
rect 13248 -5864 13300 -5831
rect 12438 -6042 12490 -5990
rect 12502 -6042 12554 -5990
rect 12566 -6042 12618 -5990
rect 12634 -6042 12686 -5990
rect 12698 -6042 12750 -5990
rect 12762 -6042 12814 -5990
rect 12924 -6042 12976 -5990
rect 12988 -6042 13040 -5990
rect 13052 -6042 13104 -5990
rect 13120 -6042 13172 -5990
rect 13184 -6042 13236 -5990
rect 13248 -6042 13300 -5990
rect 14597 -5831 14624 -5812
rect 14624 -5831 14649 -5812
rect 14597 -5864 14649 -5831
rect 14661 -5831 14662 -5812
rect 14662 -5831 14696 -5812
rect 14696 -5831 14713 -5812
rect 14661 -5864 14713 -5831
rect 14725 -5864 14777 -5812
rect 14793 -5864 14845 -5812
rect 14857 -5831 14882 -5812
rect 14882 -5831 14909 -5812
rect 14921 -5831 14954 -5812
rect 14954 -5831 14973 -5812
rect 14857 -5864 14909 -5831
rect 14921 -5864 14973 -5831
rect 15083 -5831 15106 -5812
rect 15106 -5831 15135 -5812
rect 15147 -5831 15178 -5812
rect 15178 -5831 15199 -5812
rect 15211 -5831 15212 -5812
rect 15212 -5831 15263 -5812
rect 15083 -5864 15135 -5831
rect 15147 -5864 15199 -5831
rect 15211 -5864 15263 -5831
rect 15279 -5864 15331 -5812
rect 15343 -5831 15364 -5812
rect 15364 -5831 15395 -5812
rect 15407 -5831 15436 -5812
rect 15436 -5831 15459 -5812
rect 15343 -5864 15395 -5831
rect 15407 -5864 15459 -5831
rect 14597 -6042 14649 -5990
rect 14661 -6042 14713 -5990
rect 14725 -6042 14777 -5990
rect 14793 -6042 14845 -5990
rect 14857 -6042 14909 -5990
rect 14921 -6042 14973 -5990
rect 15083 -6042 15135 -5990
rect 15147 -6042 15199 -5990
rect 15211 -6042 15263 -5990
rect 15279 -6042 15331 -5990
rect 15343 -6042 15395 -5990
rect 15407 -6042 15459 -5990
rect 12438 -6159 12490 -6129
rect 12502 -6159 12554 -6129
rect 12438 -6181 12461 -6159
rect 12461 -6181 12490 -6159
rect 12502 -6181 12533 -6159
rect 12533 -6181 12554 -6159
rect 12566 -6181 12618 -6129
rect 12634 -6159 12686 -6129
rect 12698 -6159 12750 -6129
rect 12762 -6159 12814 -6129
rect 12634 -6181 12685 -6159
rect 12685 -6181 12686 -6159
rect 12698 -6181 12719 -6159
rect 12719 -6181 12750 -6159
rect 12762 -6181 12791 -6159
rect 12791 -6181 12814 -6159
rect 12924 -6159 12976 -6129
rect 12988 -6159 13040 -6129
rect 12924 -6181 12943 -6159
rect 12943 -6181 12976 -6159
rect 12988 -6181 13015 -6159
rect 13015 -6181 13040 -6159
rect 13052 -6181 13104 -6129
rect 13120 -6181 13172 -6129
rect 13184 -6159 13236 -6129
rect 13184 -6181 13201 -6159
rect 13201 -6181 13235 -6159
rect 13235 -6181 13236 -6159
rect 13248 -6159 13300 -6129
rect 13248 -6181 13273 -6159
rect 13273 -6181 13300 -6159
rect 4577 -7062 4629 -7010
rect 4641 -7062 4693 -7010
rect 4705 -7062 4757 -7010
rect 5963 -6761 6015 -6709
rect 6027 -6761 6079 -6709
rect 6091 -6761 6143 -6709
rect 5706 -7062 5758 -7010
rect 5770 -7062 5822 -7010
rect 5834 -7062 5886 -7010
rect 6480 -6761 6532 -6709
rect 6544 -6761 6596 -6709
rect 6608 -6761 6660 -6709
rect 6223 -7062 6275 -7010
rect 6287 -7062 6339 -7010
rect 6351 -7062 6403 -7010
rect 7191 -6616 7243 -6564
rect 7255 -6616 7307 -6564
rect 7319 -6616 7371 -6564
rect 6933 -6922 6985 -6870
rect 6997 -6922 7049 -6870
rect 7061 -6922 7113 -6870
rect 6740 -7062 6792 -7010
rect 6804 -7062 6856 -7010
rect 6868 -7062 6920 -7010
rect 7708 -6616 7760 -6564
rect 7772 -6616 7824 -6564
rect 7836 -6616 7888 -6564
rect 7450 -6922 7502 -6870
rect 7514 -6922 7566 -6870
rect 7578 -6922 7630 -6870
rect 8157 -6761 8209 -6709
rect 8221 -6761 8273 -6709
rect 8285 -6761 8337 -6709
rect 7900 -7062 7952 -7010
rect 7964 -7062 8016 -7010
rect 8028 -7062 8080 -7010
rect 8674 -6761 8726 -6709
rect 8738 -6761 8790 -6709
rect 8802 -6761 8854 -6709
rect 8417 -7062 8469 -7010
rect 8481 -7062 8533 -7010
rect 8545 -7062 8597 -7010
rect 14597 -6159 14649 -6129
rect 14597 -6181 14624 -6159
rect 14624 -6181 14649 -6159
rect 14661 -6159 14713 -6129
rect 14661 -6181 14662 -6159
rect 14662 -6181 14696 -6159
rect 14696 -6181 14713 -6159
rect 14725 -6181 14777 -6129
rect 14793 -6181 14845 -6129
rect 14857 -6159 14909 -6129
rect 14921 -6159 14973 -6129
rect 14857 -6181 14882 -6159
rect 14882 -6181 14909 -6159
rect 14921 -6181 14954 -6159
rect 14954 -6181 14973 -6159
rect 15083 -6159 15135 -6129
rect 15147 -6159 15199 -6129
rect 15211 -6159 15263 -6129
rect 15083 -6181 15106 -6159
rect 15106 -6181 15135 -6159
rect 15147 -6181 15178 -6159
rect 15178 -6181 15199 -6159
rect 15211 -6181 15212 -6159
rect 15212 -6181 15263 -6159
rect 15279 -6181 15331 -6129
rect 15343 -6159 15395 -6129
rect 15407 -6159 15459 -6129
rect 15343 -6181 15364 -6159
rect 15364 -6181 15395 -6159
rect 15407 -6181 15436 -6159
rect 15436 -6181 15459 -6159
rect 15811 -6042 15863 -5990
rect 15875 -6042 15927 -5990
rect 15939 -6042 15991 -5990
rect 16007 -6042 16059 -5990
rect 16071 -6042 16123 -5990
rect 16135 -6042 16187 -5990
rect 16199 -6042 16251 -5990
rect 16267 -6042 16319 -5990
rect 16331 -6042 16383 -5990
rect 16395 -6042 16447 -5990
rect 16795 -5831 16818 -5812
rect 16818 -5831 16847 -5812
rect 16859 -5831 16890 -5812
rect 16890 -5831 16911 -5812
rect 16795 -5864 16847 -5831
rect 16859 -5864 16911 -5831
rect 16923 -5864 16975 -5812
rect 16991 -5831 17042 -5812
rect 17042 -5831 17043 -5812
rect 17055 -5831 17076 -5812
rect 17076 -5831 17107 -5812
rect 17119 -5831 17148 -5812
rect 17148 -5831 17171 -5812
rect 16991 -5864 17043 -5831
rect 17055 -5864 17107 -5831
rect 17119 -5864 17171 -5831
rect 17281 -5831 17300 -5812
rect 17300 -5831 17333 -5812
rect 17345 -5831 17372 -5812
rect 17372 -5831 17397 -5812
rect 17281 -5864 17333 -5831
rect 17345 -5864 17397 -5831
rect 17409 -5864 17461 -5812
rect 17477 -5864 17529 -5812
rect 17541 -5831 17558 -5812
rect 17558 -5831 17592 -5812
rect 17592 -5831 17593 -5812
rect 17541 -5864 17593 -5831
rect 17605 -5831 17630 -5812
rect 17630 -5831 17657 -5812
rect 17605 -5864 17657 -5831
rect 16795 -6042 16847 -5990
rect 16859 -6042 16911 -5990
rect 16923 -6042 16975 -5990
rect 16991 -6042 17043 -5990
rect 17055 -6042 17107 -5990
rect 17119 -6042 17171 -5990
rect 17281 -6042 17333 -5990
rect 17345 -6042 17397 -5990
rect 17409 -6042 17461 -5990
rect 17477 -6042 17529 -5990
rect 17541 -6042 17593 -5990
rect 17605 -6042 17657 -5990
rect 16795 -6159 16847 -6129
rect 16859 -6159 16911 -6129
rect 16795 -6181 16818 -6159
rect 16818 -6181 16847 -6159
rect 16859 -6181 16890 -6159
rect 16890 -6181 16911 -6159
rect 16923 -6181 16975 -6129
rect 16991 -6159 17043 -6129
rect 17055 -6159 17107 -6129
rect 17119 -6159 17171 -6129
rect 16991 -6181 17042 -6159
rect 17042 -6181 17043 -6159
rect 17055 -6181 17076 -6159
rect 17076 -6181 17107 -6159
rect 17119 -6181 17148 -6159
rect 17148 -6181 17171 -6159
rect 17281 -6159 17333 -6129
rect 17345 -6159 17397 -6129
rect 17281 -6181 17300 -6159
rect 17300 -6181 17333 -6159
rect 17345 -6181 17372 -6159
rect 17372 -6181 17397 -6159
rect 17409 -6181 17461 -6129
rect 17477 -6181 17529 -6129
rect 17541 -6159 17593 -6129
rect 17541 -6181 17558 -6159
rect 17558 -6181 17592 -6159
rect 17592 -6181 17593 -6159
rect 17605 -6159 17657 -6129
rect 17605 -6181 17630 -6159
rect 17630 -6181 17657 -6159
rect 8932 -7062 8984 -7010
rect 8996 -7062 9048 -7010
rect 9060 -7062 9112 -7010
rect 10326 -6761 10378 -6709
rect 10390 -6761 10442 -6709
rect 10454 -6761 10506 -6709
rect 10068 -7062 10120 -7010
rect 10132 -7062 10184 -7010
rect 10196 -7062 10248 -7010
rect 1523 -7478 1550 -7459
rect 1550 -7478 1575 -7459
rect 1523 -7511 1575 -7478
rect 1587 -7478 1588 -7459
rect 1588 -7478 1622 -7459
rect 1622 -7478 1639 -7459
rect 1587 -7511 1639 -7478
rect 1651 -7511 1703 -7459
rect 1719 -7511 1771 -7459
rect 1783 -7478 1808 -7459
rect 1808 -7478 1835 -7459
rect 1847 -7478 1880 -7459
rect 1880 -7478 1899 -7459
rect 1783 -7511 1835 -7478
rect 1847 -7511 1899 -7478
rect 2009 -7478 2032 -7459
rect 2032 -7478 2061 -7459
rect 2073 -7478 2104 -7459
rect 2104 -7478 2125 -7459
rect 2137 -7478 2138 -7459
rect 2138 -7478 2189 -7459
rect 2009 -7511 2061 -7478
rect 2073 -7511 2125 -7478
rect 2137 -7511 2189 -7478
rect 2205 -7511 2257 -7459
rect 2269 -7478 2290 -7459
rect 2290 -7478 2321 -7459
rect 2333 -7478 2362 -7459
rect 2362 -7478 2385 -7459
rect 2269 -7511 2321 -7478
rect 2333 -7511 2385 -7478
rect 1523 -7689 1575 -7637
rect 1587 -7689 1639 -7637
rect 1651 -7689 1703 -7637
rect 1719 -7689 1771 -7637
rect 1783 -7689 1835 -7637
rect 1847 -7689 1899 -7637
rect 2009 -7689 2061 -7637
rect 2073 -7689 2125 -7637
rect 2137 -7689 2189 -7637
rect 2205 -7689 2257 -7637
rect 2269 -7689 2321 -7637
rect 2333 -7689 2385 -7637
rect 1523 -7806 1575 -7776
rect 1523 -7828 1550 -7806
rect 1550 -7828 1575 -7806
rect 1587 -7806 1639 -7776
rect 1587 -7828 1588 -7806
rect 1588 -7828 1622 -7806
rect 1622 -7828 1639 -7806
rect 1651 -7828 1703 -7776
rect 1719 -7828 1771 -7776
rect 1783 -7806 1835 -7776
rect 1847 -7806 1899 -7776
rect 1783 -7828 1808 -7806
rect 1808 -7828 1835 -7806
rect 1847 -7828 1880 -7806
rect 1880 -7828 1899 -7806
rect 2009 -7806 2061 -7776
rect 2073 -7806 2125 -7776
rect 2137 -7806 2189 -7776
rect 2009 -7828 2032 -7806
rect 2032 -7828 2061 -7806
rect 2073 -7828 2104 -7806
rect 2104 -7828 2125 -7806
rect 2137 -7828 2138 -7806
rect 2138 -7828 2189 -7806
rect 2205 -7828 2257 -7776
rect 2269 -7806 2321 -7776
rect 2333 -7806 2385 -7776
rect 2269 -7828 2290 -7806
rect 2290 -7828 2321 -7806
rect 2333 -7828 2362 -7806
rect 2362 -7828 2385 -7806
rect 2733 -7689 2785 -7637
rect 2797 -7689 2849 -7637
rect 2861 -7689 2913 -7637
rect 2929 -7689 2981 -7637
rect 2993 -7689 3045 -7637
rect 3057 -7689 3109 -7637
rect 3121 -7689 3173 -7637
rect 3189 -7689 3241 -7637
rect 3253 -7689 3305 -7637
rect 3317 -7689 3369 -7637
rect 3721 -7478 3744 -7459
rect 3744 -7478 3773 -7459
rect 3785 -7478 3816 -7459
rect 3816 -7478 3837 -7459
rect 3721 -7511 3773 -7478
rect 3785 -7511 3837 -7478
rect 3849 -7511 3901 -7459
rect 3917 -7478 3968 -7459
rect 3968 -7478 3969 -7459
rect 3981 -7478 4002 -7459
rect 4002 -7478 4033 -7459
rect 4045 -7478 4074 -7459
rect 4074 -7478 4097 -7459
rect 3917 -7511 3969 -7478
rect 3981 -7511 4033 -7478
rect 4045 -7511 4097 -7478
rect 4207 -7478 4226 -7459
rect 4226 -7478 4259 -7459
rect 4271 -7478 4298 -7459
rect 4298 -7478 4323 -7459
rect 4207 -7511 4259 -7478
rect 4271 -7511 4323 -7478
rect 4335 -7511 4387 -7459
rect 4403 -7511 4455 -7459
rect 4467 -7478 4484 -7459
rect 4484 -7478 4518 -7459
rect 4518 -7478 4519 -7459
rect 4467 -7511 4519 -7478
rect 4531 -7478 4556 -7459
rect 4556 -7478 4583 -7459
rect 4531 -7511 4583 -7478
rect 3721 -7689 3773 -7637
rect 3785 -7689 3837 -7637
rect 3849 -7689 3901 -7637
rect 3917 -7689 3969 -7637
rect 3981 -7689 4033 -7637
rect 4045 -7689 4097 -7637
rect 4207 -7689 4259 -7637
rect 4271 -7689 4323 -7637
rect 4335 -7689 4387 -7637
rect 4403 -7689 4455 -7637
rect 4467 -7689 4519 -7637
rect 4531 -7689 4583 -7637
rect 10843 -6761 10895 -6709
rect 10907 -6761 10959 -6709
rect 10971 -6761 11023 -6709
rect 10583 -7062 10635 -7010
rect 10647 -7062 10699 -7010
rect 10711 -7062 10763 -7010
rect 11292 -6616 11344 -6564
rect 11356 -6616 11408 -6564
rect 11420 -6616 11472 -6564
rect 11100 -7062 11152 -7010
rect 11164 -7062 11216 -7010
rect 11228 -7062 11280 -7010
rect 11809 -6616 11861 -6564
rect 11873 -6616 11925 -6564
rect 11937 -6616 11989 -6564
rect 11550 -6922 11602 -6870
rect 11614 -6922 11666 -6870
rect 11678 -6922 11730 -6870
rect 12067 -6922 12119 -6870
rect 12131 -6922 12183 -6870
rect 12195 -6922 12247 -6870
rect 12520 -6761 12572 -6709
rect 12584 -6761 12636 -6709
rect 12648 -6761 12700 -6709
rect 12260 -7062 12312 -7010
rect 12324 -7062 12376 -7010
rect 12388 -7062 12440 -7010
rect 13037 -6761 13089 -6709
rect 13101 -6761 13153 -6709
rect 13165 -6761 13217 -6709
rect 12777 -7062 12829 -7010
rect 12841 -7062 12893 -7010
rect 12905 -7062 12957 -7010
rect 13294 -7062 13346 -7010
rect 13358 -7062 13410 -7010
rect 13422 -7062 13474 -7010
rect 14680 -6761 14732 -6709
rect 14744 -6761 14796 -6709
rect 14808 -6761 14860 -6709
rect 14423 -7062 14475 -7010
rect 14487 -7062 14539 -7010
rect 14551 -7062 14603 -7010
rect 5880 -7478 5907 -7459
rect 5907 -7478 5932 -7459
rect 5880 -7511 5932 -7478
rect 5944 -7478 5945 -7459
rect 5945 -7478 5979 -7459
rect 5979 -7478 5996 -7459
rect 5944 -7511 5996 -7478
rect 6008 -7511 6060 -7459
rect 6076 -7511 6128 -7459
rect 6140 -7478 6165 -7459
rect 6165 -7478 6192 -7459
rect 6204 -7478 6237 -7459
rect 6237 -7478 6256 -7459
rect 6140 -7511 6192 -7478
rect 6204 -7511 6256 -7478
rect 6366 -7478 6389 -7459
rect 6389 -7478 6418 -7459
rect 6430 -7478 6461 -7459
rect 6461 -7478 6482 -7459
rect 6494 -7478 6495 -7459
rect 6495 -7478 6546 -7459
rect 6366 -7511 6418 -7478
rect 6430 -7511 6482 -7478
rect 6494 -7511 6546 -7478
rect 6562 -7511 6614 -7459
rect 6626 -7478 6647 -7459
rect 6647 -7478 6678 -7459
rect 6690 -7478 6719 -7459
rect 6719 -7478 6742 -7459
rect 6626 -7511 6678 -7478
rect 6690 -7511 6742 -7478
rect 5880 -7689 5932 -7637
rect 5944 -7689 5996 -7637
rect 6008 -7689 6060 -7637
rect 6076 -7689 6128 -7637
rect 6140 -7689 6192 -7637
rect 6204 -7689 6256 -7637
rect 6366 -7689 6418 -7637
rect 6430 -7689 6482 -7637
rect 6494 -7689 6546 -7637
rect 6562 -7689 6614 -7637
rect 6626 -7689 6678 -7637
rect 6690 -7689 6742 -7637
rect 3721 -7806 3773 -7776
rect 3785 -7806 3837 -7776
rect 3721 -7828 3744 -7806
rect 3744 -7828 3773 -7806
rect 3785 -7828 3816 -7806
rect 3816 -7828 3837 -7806
rect 3849 -7828 3901 -7776
rect 3917 -7806 3969 -7776
rect 3981 -7806 4033 -7776
rect 4045 -7806 4097 -7776
rect 3917 -7828 3968 -7806
rect 3968 -7828 3969 -7806
rect 3981 -7828 4002 -7806
rect 4002 -7828 4033 -7806
rect 4045 -7828 4074 -7806
rect 4074 -7828 4097 -7806
rect 4207 -7806 4259 -7776
rect 4271 -7806 4323 -7776
rect 4207 -7828 4226 -7806
rect 4226 -7828 4259 -7806
rect 4271 -7828 4298 -7806
rect 4298 -7828 4323 -7806
rect 4335 -7828 4387 -7776
rect 4403 -7828 4455 -7776
rect 4467 -7806 4519 -7776
rect 4467 -7828 4484 -7806
rect 4484 -7828 4518 -7806
rect 4518 -7828 4519 -7806
rect 4531 -7806 4583 -7776
rect 4531 -7828 4556 -7806
rect 4556 -7828 4583 -7806
rect 5880 -7806 5932 -7776
rect 5880 -7828 5907 -7806
rect 5907 -7828 5932 -7806
rect 5944 -7806 5996 -7776
rect 5944 -7828 5945 -7806
rect 5945 -7828 5979 -7806
rect 5979 -7828 5996 -7806
rect 6008 -7828 6060 -7776
rect 6076 -7828 6128 -7776
rect 6140 -7806 6192 -7776
rect 6204 -7806 6256 -7776
rect 6140 -7828 6165 -7806
rect 6165 -7828 6192 -7806
rect 6204 -7828 6237 -7806
rect 6237 -7828 6256 -7806
rect 6366 -7806 6418 -7776
rect 6430 -7806 6482 -7776
rect 6494 -7806 6546 -7776
rect 6366 -7828 6389 -7806
rect 6389 -7828 6418 -7806
rect 6430 -7828 6461 -7806
rect 6461 -7828 6482 -7806
rect 6494 -7828 6495 -7806
rect 6495 -7828 6546 -7806
rect 6562 -7828 6614 -7776
rect 6626 -7806 6678 -7776
rect 6690 -7806 6742 -7776
rect 6626 -7828 6647 -7806
rect 6647 -7828 6678 -7806
rect 6690 -7828 6719 -7806
rect 6719 -7828 6742 -7806
rect 7094 -7689 7146 -7637
rect 7158 -7689 7210 -7637
rect 7222 -7689 7274 -7637
rect 7290 -7689 7342 -7637
rect 7354 -7689 7406 -7637
rect 7418 -7689 7470 -7637
rect 7482 -7689 7534 -7637
rect 7550 -7689 7602 -7637
rect 7614 -7689 7666 -7637
rect 7678 -7689 7730 -7637
rect 8078 -7478 8101 -7459
rect 8101 -7478 8130 -7459
rect 8142 -7478 8173 -7459
rect 8173 -7478 8194 -7459
rect 8078 -7511 8130 -7478
rect 8142 -7511 8194 -7478
rect 8206 -7511 8258 -7459
rect 8274 -7478 8325 -7459
rect 8325 -7478 8326 -7459
rect 8338 -7478 8359 -7459
rect 8359 -7478 8390 -7459
rect 8402 -7478 8431 -7459
rect 8431 -7478 8454 -7459
rect 8274 -7511 8326 -7478
rect 8338 -7511 8390 -7478
rect 8402 -7511 8454 -7478
rect 8564 -7478 8583 -7459
rect 8583 -7478 8616 -7459
rect 8628 -7478 8655 -7459
rect 8655 -7478 8680 -7459
rect 8564 -7511 8616 -7478
rect 8628 -7511 8680 -7478
rect 8692 -7511 8744 -7459
rect 8760 -7511 8812 -7459
rect 8824 -7478 8841 -7459
rect 8841 -7478 8875 -7459
rect 8875 -7478 8876 -7459
rect 8824 -7511 8876 -7478
rect 8888 -7478 8913 -7459
rect 8913 -7478 8940 -7459
rect 8888 -7511 8940 -7478
rect 8078 -7689 8130 -7637
rect 8142 -7689 8194 -7637
rect 8206 -7689 8258 -7637
rect 8274 -7689 8326 -7637
rect 8338 -7689 8390 -7637
rect 8402 -7689 8454 -7637
rect 8564 -7689 8616 -7637
rect 8628 -7689 8680 -7637
rect 8692 -7689 8744 -7637
rect 8760 -7689 8812 -7637
rect 8824 -7689 8876 -7637
rect 8888 -7689 8940 -7637
rect 15197 -6761 15249 -6709
rect 15261 -6761 15313 -6709
rect 15325 -6761 15377 -6709
rect 14940 -7062 14992 -7010
rect 15004 -7062 15056 -7010
rect 15068 -7062 15120 -7010
rect 15908 -6616 15960 -6564
rect 15972 -6616 16024 -6564
rect 16036 -6616 16088 -6564
rect 15650 -6922 15702 -6870
rect 15714 -6922 15766 -6870
rect 15778 -6922 15830 -6870
rect 15457 -7062 15509 -7010
rect 15521 -7062 15573 -7010
rect 15585 -7062 15637 -7010
rect 16425 -6616 16477 -6564
rect 16489 -6616 16541 -6564
rect 16553 -6616 16605 -6564
rect 16167 -6922 16219 -6870
rect 16231 -6922 16283 -6870
rect 16295 -6922 16347 -6870
rect 16874 -6761 16926 -6709
rect 16938 -6761 16990 -6709
rect 17002 -6761 17054 -6709
rect 16617 -7062 16669 -7010
rect 16681 -7062 16733 -7010
rect 16745 -7062 16797 -7010
rect 17392 -6761 17444 -6709
rect 17456 -6761 17508 -6709
rect 17520 -6761 17572 -6709
rect 17135 -7062 17187 -7010
rect 17199 -7062 17251 -7010
rect 17263 -7062 17315 -7010
rect 17650 -7062 17702 -7010
rect 17714 -7062 17766 -7010
rect 17778 -7062 17830 -7010
rect 10240 -7478 10267 -7459
rect 10267 -7478 10292 -7459
rect 10240 -7511 10292 -7478
rect 10304 -7478 10305 -7459
rect 10305 -7478 10339 -7459
rect 10339 -7478 10356 -7459
rect 10304 -7511 10356 -7478
rect 10368 -7511 10420 -7459
rect 10436 -7511 10488 -7459
rect 10500 -7478 10525 -7459
rect 10525 -7478 10552 -7459
rect 10564 -7478 10597 -7459
rect 10597 -7478 10616 -7459
rect 10500 -7511 10552 -7478
rect 10564 -7511 10616 -7478
rect 10726 -7478 10749 -7459
rect 10749 -7478 10778 -7459
rect 10790 -7478 10821 -7459
rect 10821 -7478 10842 -7459
rect 10854 -7478 10855 -7459
rect 10855 -7478 10906 -7459
rect 10726 -7511 10778 -7478
rect 10790 -7511 10842 -7478
rect 10854 -7511 10906 -7478
rect 10922 -7511 10974 -7459
rect 10986 -7478 11007 -7459
rect 11007 -7478 11038 -7459
rect 11050 -7478 11079 -7459
rect 11079 -7478 11102 -7459
rect 10986 -7511 11038 -7478
rect 11050 -7511 11102 -7478
rect 10240 -7689 10292 -7637
rect 10304 -7689 10356 -7637
rect 10368 -7689 10420 -7637
rect 10436 -7689 10488 -7637
rect 10500 -7689 10552 -7637
rect 10564 -7689 10616 -7637
rect 10726 -7689 10778 -7637
rect 10790 -7689 10842 -7637
rect 10854 -7689 10906 -7637
rect 10922 -7689 10974 -7637
rect 10986 -7689 11038 -7637
rect 11050 -7689 11102 -7637
rect 8078 -7806 8130 -7776
rect 8142 -7806 8194 -7776
rect 8078 -7828 8101 -7806
rect 8101 -7828 8130 -7806
rect 8142 -7828 8173 -7806
rect 8173 -7828 8194 -7806
rect 8206 -7828 8258 -7776
rect 8274 -7806 8326 -7776
rect 8338 -7806 8390 -7776
rect 8402 -7806 8454 -7776
rect 8274 -7828 8325 -7806
rect 8325 -7828 8326 -7806
rect 8338 -7828 8359 -7806
rect 8359 -7828 8390 -7806
rect 8402 -7828 8431 -7806
rect 8431 -7828 8454 -7806
rect 8564 -7806 8616 -7776
rect 8628 -7806 8680 -7776
rect 8564 -7828 8583 -7806
rect 8583 -7828 8616 -7806
rect 8628 -7828 8655 -7806
rect 8655 -7828 8680 -7806
rect 8692 -7828 8744 -7776
rect 8760 -7828 8812 -7776
rect 8824 -7806 8876 -7776
rect 8824 -7828 8841 -7806
rect 8841 -7828 8875 -7806
rect 8875 -7828 8876 -7806
rect 8888 -7806 8940 -7776
rect 8888 -7828 8913 -7806
rect 8913 -7828 8940 -7806
rect 10240 -7806 10292 -7776
rect 10240 -7828 10267 -7806
rect 10267 -7828 10292 -7806
rect 10304 -7806 10356 -7776
rect 10304 -7828 10305 -7806
rect 10305 -7828 10339 -7806
rect 10339 -7828 10356 -7806
rect 10368 -7828 10420 -7776
rect 10436 -7828 10488 -7776
rect 10500 -7806 10552 -7776
rect 10564 -7806 10616 -7776
rect 10500 -7828 10525 -7806
rect 10525 -7828 10552 -7806
rect 10564 -7828 10597 -7806
rect 10597 -7828 10616 -7806
rect 10726 -7806 10778 -7776
rect 10790 -7806 10842 -7776
rect 10854 -7806 10906 -7776
rect 10726 -7828 10749 -7806
rect 10749 -7828 10778 -7806
rect 10790 -7828 10821 -7806
rect 10821 -7828 10842 -7806
rect 10854 -7828 10855 -7806
rect 10855 -7828 10906 -7806
rect 10922 -7828 10974 -7776
rect 10986 -7806 11038 -7776
rect 11050 -7806 11102 -7776
rect 10986 -7828 11007 -7806
rect 11007 -7828 11038 -7806
rect 11050 -7828 11079 -7806
rect 11079 -7828 11102 -7806
rect 11450 -7689 11502 -7637
rect 11514 -7689 11566 -7637
rect 11578 -7689 11630 -7637
rect 11646 -7689 11698 -7637
rect 11710 -7689 11762 -7637
rect 11774 -7689 11826 -7637
rect 11838 -7689 11890 -7637
rect 11906 -7689 11958 -7637
rect 11970 -7689 12022 -7637
rect 12034 -7689 12086 -7637
rect 12438 -7478 12461 -7459
rect 12461 -7478 12490 -7459
rect 12502 -7478 12533 -7459
rect 12533 -7478 12554 -7459
rect 12438 -7511 12490 -7478
rect 12502 -7511 12554 -7478
rect 12566 -7511 12618 -7459
rect 12634 -7478 12685 -7459
rect 12685 -7478 12686 -7459
rect 12698 -7478 12719 -7459
rect 12719 -7478 12750 -7459
rect 12762 -7478 12791 -7459
rect 12791 -7478 12814 -7459
rect 12634 -7511 12686 -7478
rect 12698 -7511 12750 -7478
rect 12762 -7511 12814 -7478
rect 12924 -7478 12943 -7459
rect 12943 -7478 12976 -7459
rect 12988 -7478 13015 -7459
rect 13015 -7478 13040 -7459
rect 12924 -7511 12976 -7478
rect 12988 -7511 13040 -7478
rect 13052 -7511 13104 -7459
rect 13120 -7511 13172 -7459
rect 13184 -7478 13201 -7459
rect 13201 -7478 13235 -7459
rect 13235 -7478 13236 -7459
rect 13184 -7511 13236 -7478
rect 13248 -7478 13273 -7459
rect 13273 -7478 13300 -7459
rect 13248 -7511 13300 -7478
rect 12438 -7689 12490 -7637
rect 12502 -7689 12554 -7637
rect 12566 -7689 12618 -7637
rect 12634 -7689 12686 -7637
rect 12698 -7689 12750 -7637
rect 12762 -7689 12814 -7637
rect 12924 -7689 12976 -7637
rect 12988 -7689 13040 -7637
rect 13052 -7689 13104 -7637
rect 13120 -7689 13172 -7637
rect 13184 -7689 13236 -7637
rect 13248 -7689 13300 -7637
rect 14597 -7478 14624 -7459
rect 14624 -7478 14649 -7459
rect 14597 -7511 14649 -7478
rect 14661 -7478 14662 -7459
rect 14662 -7478 14696 -7459
rect 14696 -7478 14713 -7459
rect 14661 -7511 14713 -7478
rect 14725 -7511 14777 -7459
rect 14793 -7511 14845 -7459
rect 14857 -7478 14882 -7459
rect 14882 -7478 14909 -7459
rect 14921 -7478 14954 -7459
rect 14954 -7478 14973 -7459
rect 14857 -7511 14909 -7478
rect 14921 -7511 14973 -7478
rect 15083 -7478 15106 -7459
rect 15106 -7478 15135 -7459
rect 15147 -7478 15178 -7459
rect 15178 -7478 15199 -7459
rect 15211 -7478 15212 -7459
rect 15212 -7478 15263 -7459
rect 15083 -7511 15135 -7478
rect 15147 -7511 15199 -7478
rect 15211 -7511 15263 -7478
rect 15279 -7511 15331 -7459
rect 15343 -7478 15364 -7459
rect 15364 -7478 15395 -7459
rect 15407 -7478 15436 -7459
rect 15436 -7478 15459 -7459
rect 15343 -7511 15395 -7478
rect 15407 -7511 15459 -7478
rect 14597 -7689 14649 -7637
rect 14661 -7689 14713 -7637
rect 14725 -7689 14777 -7637
rect 14793 -7689 14845 -7637
rect 14857 -7689 14909 -7637
rect 14921 -7689 14973 -7637
rect 15083 -7689 15135 -7637
rect 15147 -7689 15199 -7637
rect 15211 -7689 15263 -7637
rect 15279 -7689 15331 -7637
rect 15343 -7689 15395 -7637
rect 15407 -7689 15459 -7637
rect 12438 -7806 12490 -7776
rect 12502 -7806 12554 -7776
rect 12438 -7828 12461 -7806
rect 12461 -7828 12490 -7806
rect 12502 -7828 12533 -7806
rect 12533 -7828 12554 -7806
rect 12566 -7828 12618 -7776
rect 12634 -7806 12686 -7776
rect 12698 -7806 12750 -7776
rect 12762 -7806 12814 -7776
rect 12634 -7828 12685 -7806
rect 12685 -7828 12686 -7806
rect 12698 -7828 12719 -7806
rect 12719 -7828 12750 -7806
rect 12762 -7828 12791 -7806
rect 12791 -7828 12814 -7806
rect 12924 -7806 12976 -7776
rect 12988 -7806 13040 -7776
rect 12924 -7828 12943 -7806
rect 12943 -7828 12976 -7806
rect 12988 -7828 13015 -7806
rect 13015 -7828 13040 -7806
rect 13052 -7828 13104 -7776
rect 13120 -7828 13172 -7776
rect 13184 -7806 13236 -7776
rect 13184 -7828 13201 -7806
rect 13201 -7828 13235 -7806
rect 13235 -7828 13236 -7806
rect 13248 -7806 13300 -7776
rect 13248 -7828 13273 -7806
rect 13273 -7828 13300 -7806
rect 14597 -7806 14649 -7776
rect 14597 -7828 14624 -7806
rect 14624 -7828 14649 -7806
rect 14661 -7806 14713 -7776
rect 14661 -7828 14662 -7806
rect 14662 -7828 14696 -7806
rect 14696 -7828 14713 -7806
rect 14725 -7828 14777 -7776
rect 14793 -7828 14845 -7776
rect 14857 -7806 14909 -7776
rect 14921 -7806 14973 -7776
rect 14857 -7828 14882 -7806
rect 14882 -7828 14909 -7806
rect 14921 -7828 14954 -7806
rect 14954 -7828 14973 -7806
rect 15083 -7806 15135 -7776
rect 15147 -7806 15199 -7776
rect 15211 -7806 15263 -7776
rect 15083 -7828 15106 -7806
rect 15106 -7828 15135 -7806
rect 15147 -7828 15178 -7806
rect 15178 -7828 15199 -7806
rect 15211 -7828 15212 -7806
rect 15212 -7828 15263 -7806
rect 15279 -7828 15331 -7776
rect 15343 -7806 15395 -7776
rect 15407 -7806 15459 -7776
rect 15343 -7828 15364 -7806
rect 15364 -7828 15395 -7806
rect 15407 -7828 15436 -7806
rect 15436 -7828 15459 -7806
rect 15811 -7689 15863 -7637
rect 15875 -7689 15927 -7637
rect 15939 -7689 15991 -7637
rect 16007 -7689 16059 -7637
rect 16071 -7689 16123 -7637
rect 16135 -7689 16187 -7637
rect 16199 -7689 16251 -7637
rect 16267 -7689 16319 -7637
rect 16331 -7689 16383 -7637
rect 16395 -7689 16447 -7637
rect 16795 -7478 16818 -7459
rect 16818 -7478 16847 -7459
rect 16859 -7478 16890 -7459
rect 16890 -7478 16911 -7459
rect 16795 -7511 16847 -7478
rect 16859 -7511 16911 -7478
rect 16923 -7511 16975 -7459
rect 16991 -7478 17042 -7459
rect 17042 -7478 17043 -7459
rect 17055 -7478 17076 -7459
rect 17076 -7478 17107 -7459
rect 17119 -7478 17148 -7459
rect 17148 -7478 17171 -7459
rect 16991 -7511 17043 -7478
rect 17055 -7511 17107 -7478
rect 17119 -7511 17171 -7478
rect 17281 -7478 17300 -7459
rect 17300 -7478 17333 -7459
rect 17345 -7478 17372 -7459
rect 17372 -7478 17397 -7459
rect 17281 -7511 17333 -7478
rect 17345 -7511 17397 -7478
rect 17409 -7511 17461 -7459
rect 17477 -7511 17529 -7459
rect 17541 -7478 17558 -7459
rect 17558 -7478 17592 -7459
rect 17592 -7478 17593 -7459
rect 17541 -7511 17593 -7478
rect 17605 -7478 17630 -7459
rect 17630 -7478 17657 -7459
rect 17605 -7511 17657 -7478
rect 16795 -7689 16847 -7637
rect 16859 -7689 16911 -7637
rect 16923 -7689 16975 -7637
rect 16991 -7689 17043 -7637
rect 17055 -7689 17107 -7637
rect 17119 -7689 17171 -7637
rect 17281 -7689 17333 -7637
rect 17345 -7689 17397 -7637
rect 17409 -7689 17461 -7637
rect 17477 -7689 17529 -7637
rect 17541 -7689 17593 -7637
rect 17605 -7689 17657 -7637
rect 16795 -7806 16847 -7776
rect 16859 -7806 16911 -7776
rect 16795 -7828 16818 -7806
rect 16818 -7828 16847 -7806
rect 16859 -7828 16890 -7806
rect 16890 -7828 16911 -7806
rect 16923 -7828 16975 -7776
rect 16991 -7806 17043 -7776
rect 17055 -7806 17107 -7776
rect 17119 -7806 17171 -7776
rect 16991 -7828 17042 -7806
rect 17042 -7828 17043 -7806
rect 17055 -7828 17076 -7806
rect 17076 -7828 17107 -7806
rect 17119 -7828 17148 -7806
rect 17148 -7828 17171 -7806
rect 17281 -7806 17333 -7776
rect 17345 -7806 17397 -7776
rect 17281 -7828 17300 -7806
rect 17300 -7828 17333 -7806
rect 17345 -7828 17372 -7806
rect 17372 -7828 17397 -7806
rect 17409 -7828 17461 -7776
rect 17477 -7828 17529 -7776
rect 17541 -7806 17593 -7776
rect 17541 -7828 17558 -7806
rect 17558 -7828 17592 -7806
rect 17592 -7828 17593 -7806
rect 17605 -7806 17657 -7776
rect 17605 -7828 17630 -7806
rect 17630 -7828 17657 -7806
rect 1607 -8251 1659 -8199
rect 1671 -8251 1723 -8199
rect 1735 -8251 1787 -8199
rect 2125 -8251 2177 -8199
rect 2189 -8251 2241 -8199
rect 2253 -8251 2305 -8199
rect 2577 -8420 2629 -8368
rect 2641 -8420 2693 -8368
rect 2705 -8420 2757 -8368
rect 1348 -8583 1400 -8531
rect 1412 -8583 1464 -8531
rect 1476 -8583 1528 -8531
rect 1865 -8583 1917 -8531
rect 1929 -8583 1981 -8531
rect 1993 -8583 2045 -8531
rect 2382 -8583 2434 -8531
rect 2446 -8583 2498 -8531
rect 2510 -8583 2562 -8531
rect 3094 -8420 3146 -8368
rect 3158 -8420 3210 -8368
rect 3222 -8420 3274 -8368
rect 3802 -8251 3854 -8199
rect 3866 -8251 3918 -8199
rect 3930 -8251 3982 -8199
rect 4319 -8251 4371 -8199
rect 4383 -8251 4435 -8199
rect 4447 -8251 4499 -8199
rect 3543 -8583 3595 -8531
rect 3607 -8583 3659 -8531
rect 3671 -8583 3723 -8531
rect 4060 -8583 4112 -8531
rect 4124 -8583 4176 -8531
rect 4188 -8583 4240 -8531
rect 4575 -8583 4627 -8531
rect 4639 -8583 4691 -8531
rect 4703 -8583 4755 -8531
rect 5964 -8251 6016 -8199
rect 6028 -8251 6080 -8199
rect 6092 -8251 6144 -8199
rect 6481 -8251 6533 -8199
rect 6545 -8251 6597 -8199
rect 6609 -8251 6661 -8199
rect 5708 -8583 5760 -8531
rect 5772 -8583 5824 -8531
rect 5836 -8583 5888 -8531
rect 6223 -8583 6275 -8531
rect 6287 -8583 6339 -8531
rect 6351 -8583 6403 -8531
rect 6740 -8583 6792 -8531
rect 6804 -8583 6856 -8531
rect 6868 -8583 6920 -8531
rect 2834 -8751 2886 -8699
rect 2898 -8751 2950 -8699
rect 2962 -8751 3014 -8699
rect 3351 -8751 3403 -8699
rect 3415 -8751 3467 -8699
rect 3479 -8751 3531 -8699
rect 7189 -8420 7241 -8368
rect 7253 -8420 7305 -8368
rect 7317 -8420 7369 -8368
rect 7706 -8420 7758 -8368
rect 7770 -8420 7822 -8368
rect 7834 -8420 7886 -8368
rect 8158 -8251 8210 -8199
rect 8222 -8251 8274 -8199
rect 8286 -8251 8338 -8199
rect 8675 -8251 8727 -8199
rect 8739 -8251 8791 -8199
rect 8803 -8251 8855 -8199
rect 7901 -8583 7953 -8531
rect 7965 -8583 8017 -8531
rect 8029 -8583 8081 -8531
rect 8417 -8583 8469 -8531
rect 8481 -8583 8533 -8531
rect 8545 -8583 8597 -8531
rect 8935 -8583 8987 -8531
rect 8999 -8583 9051 -8531
rect 9063 -8583 9115 -8531
rect 10325 -8251 10377 -8199
rect 10389 -8251 10441 -8199
rect 10453 -8251 10505 -8199
rect 10842 -8251 10894 -8199
rect 10906 -8251 10958 -8199
rect 10970 -8251 11022 -8199
rect 11294 -8420 11346 -8368
rect 11358 -8420 11410 -8368
rect 11422 -8420 11474 -8368
rect 10065 -8583 10117 -8531
rect 10129 -8583 10181 -8531
rect 10193 -8583 10245 -8531
rect 10583 -8583 10635 -8531
rect 10647 -8583 10699 -8531
rect 10711 -8583 10763 -8531
rect 11099 -8583 11151 -8531
rect 11163 -8583 11215 -8531
rect 11227 -8583 11279 -8531
rect 6931 -8751 6983 -8699
rect 6995 -8751 7047 -8699
rect 7059 -8751 7111 -8699
rect 7449 -8751 7501 -8699
rect 7513 -8751 7565 -8699
rect 7577 -8751 7629 -8699
rect 11811 -8420 11863 -8368
rect 11875 -8420 11927 -8368
rect 11939 -8420 11991 -8368
rect 12519 -8251 12571 -8199
rect 12583 -8251 12635 -8199
rect 12647 -8251 12699 -8199
rect 13036 -8251 13088 -8199
rect 13100 -8251 13152 -8199
rect 13164 -8251 13216 -8199
rect 12260 -8583 12312 -8531
rect 12324 -8583 12376 -8531
rect 12388 -8583 12440 -8531
rect 12777 -8583 12829 -8531
rect 12841 -8583 12893 -8531
rect 12905 -8583 12957 -8531
rect 13292 -8583 13344 -8531
rect 13356 -8583 13408 -8531
rect 13420 -8583 13472 -8531
rect 14681 -8251 14733 -8199
rect 14745 -8251 14797 -8199
rect 14809 -8251 14861 -8199
rect 15198 -8251 15250 -8199
rect 15262 -8251 15314 -8199
rect 15326 -8251 15378 -8199
rect 14425 -8583 14477 -8531
rect 14489 -8583 14541 -8531
rect 14553 -8583 14605 -8531
rect 14940 -8583 14992 -8531
rect 15004 -8583 15056 -8531
rect 15068 -8583 15120 -8531
rect 15457 -8583 15509 -8531
rect 15521 -8583 15573 -8531
rect 15585 -8583 15637 -8531
rect 11551 -8751 11603 -8699
rect 11615 -8751 11667 -8699
rect 11679 -8751 11731 -8699
rect 12069 -8751 12121 -8699
rect 12133 -8751 12185 -8699
rect 12197 -8751 12249 -8699
rect 15906 -8420 15958 -8368
rect 15970 -8420 16022 -8368
rect 16034 -8420 16086 -8368
rect 16423 -8420 16475 -8368
rect 16487 -8420 16539 -8368
rect 16551 -8420 16603 -8368
rect 16875 -8251 16927 -8199
rect 16939 -8251 16991 -8199
rect 17003 -8251 17055 -8199
rect 17393 -8251 17445 -8199
rect 17457 -8251 17509 -8199
rect 17521 -8251 17573 -8199
rect 16618 -8583 16670 -8531
rect 16682 -8583 16734 -8531
rect 16746 -8583 16798 -8531
rect 17135 -8583 17187 -8531
rect 17199 -8583 17251 -8531
rect 17263 -8583 17315 -8531
rect 17652 -8583 17704 -8531
rect 17716 -8583 17768 -8531
rect 17780 -8583 17832 -8531
rect 15649 -8751 15701 -8699
rect 15713 -8751 15765 -8699
rect 15777 -8751 15829 -8699
rect 16166 -8751 16218 -8699
rect 16230 -8751 16282 -8699
rect 16294 -8751 16346 -8699
<< metal2 >>
rect 2827 4 16353 26
rect 2827 -12 4985 4
rect 2827 -64 2834 -12
rect 2886 -64 2898 -12
rect 2950 -64 2962 -12
rect 3014 -64 3351 -12
rect 3403 -64 3415 -12
rect 3467 -64 3479 -12
rect 3531 -52 4985 -12
rect 5041 -52 5065 4
rect 5121 -52 5145 4
rect 5201 -52 5262 4
rect 5318 -52 5342 4
rect 5398 -52 5422 4
rect 5478 -12 13702 4
rect 5478 -52 6931 -12
rect 3531 -64 6931 -52
rect 6983 -64 6995 -12
rect 7047 -64 7059 -12
rect 7111 -64 7449 -12
rect 7501 -64 7513 -12
rect 7565 -64 7577 -12
rect 7629 -64 11551 -12
rect 11603 -64 11615 -12
rect 11667 -64 11679 -12
rect 11731 -64 12069 -12
rect 12121 -64 12133 -12
rect 12185 -64 12197 -12
rect 12249 -52 13702 -12
rect 13758 -52 13782 4
rect 13838 -52 13862 4
rect 13918 -52 13979 4
rect 14035 -52 14059 4
rect 14115 -52 14139 4
rect 14195 -12 16353 4
rect 14195 -52 15649 -12
rect 12249 -64 15649 -52
rect 15701 -64 15713 -12
rect 15765 -64 15777 -12
rect 15829 -64 16166 -12
rect 16218 -64 16230 -12
rect 16282 -64 16294 -12
rect 16346 -64 16353 -12
rect 2827 -74 16353 -64
rect 876 -165 18304 -143
rect 876 -221 916 -165
rect 972 -221 996 -165
rect 1052 -221 1076 -165
rect 1132 -181 9331 -165
rect 1132 -221 1348 -181
rect 876 -233 1348 -221
rect 1400 -233 1412 -181
rect 1464 -233 1476 -181
rect 1528 -233 1865 -181
rect 1917 -233 1929 -181
rect 1981 -233 1993 -181
rect 2045 -233 2382 -181
rect 2434 -233 2446 -181
rect 2498 -233 2510 -181
rect 2562 -233 3543 -181
rect 3595 -233 3607 -181
rect 3659 -233 3671 -181
rect 3723 -233 4060 -181
rect 4112 -233 4124 -181
rect 4176 -233 4188 -181
rect 4240 -233 4575 -181
rect 4627 -233 4639 -181
rect 4691 -233 4703 -181
rect 4755 -233 5708 -181
rect 5760 -233 5772 -181
rect 5824 -233 5836 -181
rect 5888 -233 6223 -181
rect 6275 -233 6287 -181
rect 6339 -233 6351 -181
rect 6403 -233 6740 -181
rect 6792 -233 6804 -181
rect 6856 -233 6868 -181
rect 6920 -233 7901 -181
rect 7953 -233 7965 -181
rect 8017 -233 8029 -181
rect 8081 -233 8417 -181
rect 8469 -233 8481 -181
rect 8533 -233 8545 -181
rect 8597 -233 8935 -181
rect 8987 -233 8999 -181
rect 9051 -233 9063 -181
rect 9115 -221 9331 -181
rect 9387 -221 9411 -165
rect 9467 -221 9491 -165
rect 9547 -221 9633 -165
rect 9689 -221 9713 -165
rect 9769 -221 9793 -165
rect 9849 -181 18048 -165
rect 9849 -221 10065 -181
rect 9115 -233 10065 -221
rect 10117 -233 10129 -181
rect 10181 -233 10193 -181
rect 10245 -233 10583 -181
rect 10635 -233 10647 -181
rect 10699 -233 10711 -181
rect 10763 -233 11099 -181
rect 11151 -233 11163 -181
rect 11215 -233 11227 -181
rect 11279 -233 12260 -181
rect 12312 -233 12324 -181
rect 12376 -233 12388 -181
rect 12440 -233 12777 -181
rect 12829 -233 12841 -181
rect 12893 -233 12905 -181
rect 12957 -233 13292 -181
rect 13344 -233 13356 -181
rect 13408 -233 13420 -181
rect 13472 -233 14425 -181
rect 14477 -233 14489 -181
rect 14541 -233 14553 -181
rect 14605 -233 14940 -181
rect 14992 -233 15004 -181
rect 15056 -233 15068 -181
rect 15120 -233 15457 -181
rect 15509 -233 15521 -181
rect 15573 -233 15585 -181
rect 15637 -233 16618 -181
rect 16670 -233 16682 -181
rect 16734 -233 16746 -181
rect 16798 -233 17135 -181
rect 17187 -233 17199 -181
rect 17251 -233 17263 -181
rect 17315 -233 17652 -181
rect 17704 -233 17716 -181
rect 17768 -233 17780 -181
rect 17832 -221 18048 -181
rect 18104 -221 18128 -165
rect 18184 -221 18208 -165
rect 18264 -221 18304 -165
rect 17832 -233 18304 -221
rect 876 -243 18304 -233
rect 2570 -328 16610 -306
rect 2570 -344 4550 -328
rect 2570 -396 2577 -344
rect 2629 -396 2641 -344
rect 2693 -396 2705 -344
rect 2757 -396 3094 -344
rect 3146 -396 3158 -344
rect 3210 -396 3222 -344
rect 3274 -384 4550 -344
rect 4606 -384 4630 -328
rect 4686 -384 4710 -328
rect 4766 -384 5697 -328
rect 5753 -384 5777 -328
rect 5833 -384 5857 -328
rect 5913 -344 13267 -328
rect 5913 -384 7189 -344
rect 3274 -396 7189 -384
rect 7241 -396 7253 -344
rect 7305 -396 7317 -344
rect 7369 -396 7706 -344
rect 7758 -396 7770 -344
rect 7822 -396 7834 -344
rect 7886 -396 11294 -344
rect 11346 -396 11358 -344
rect 11410 -396 11422 -344
rect 11474 -396 11811 -344
rect 11863 -396 11875 -344
rect 11927 -396 11939 -344
rect 11991 -384 13267 -344
rect 13323 -384 13347 -328
rect 13403 -384 13427 -328
rect 13483 -384 14414 -328
rect 14470 -384 14494 -328
rect 14550 -384 14574 -328
rect 14630 -344 16610 -328
rect 14630 -384 15906 -344
rect 11991 -396 15906 -384
rect 15958 -396 15970 -344
rect 16022 -396 16034 -344
rect 16086 -396 16423 -344
rect 16475 -396 16487 -344
rect 16539 -396 16551 -344
rect 16603 -396 16610 -344
rect 2570 -406 16610 -396
rect 1298 -496 17882 -474
rect 1298 -552 1338 -496
rect 1394 -552 1418 -496
rect 1474 -552 1498 -496
rect 1554 -512 8908 -496
rect 1554 -552 1607 -512
rect 1298 -564 1607 -552
rect 1659 -564 1671 -512
rect 1723 -564 1735 -512
rect 1787 -564 2125 -512
rect 2177 -564 2189 -512
rect 2241 -564 2253 -512
rect 2305 -564 3802 -512
rect 3854 -564 3866 -512
rect 3918 -564 3930 -512
rect 3982 -564 4319 -512
rect 4371 -564 4383 -512
rect 4435 -564 4447 -512
rect 4499 -564 5964 -512
rect 6016 -564 6028 -512
rect 6080 -564 6092 -512
rect 6144 -564 6481 -512
rect 6533 -564 6545 -512
rect 6597 -564 6609 -512
rect 6661 -564 8158 -512
rect 8210 -564 8222 -512
rect 8274 -564 8286 -512
rect 8338 -564 8675 -512
rect 8727 -564 8739 -512
rect 8791 -564 8803 -512
rect 8855 -552 8908 -512
rect 8964 -552 8988 -496
rect 9044 -552 9068 -496
rect 9124 -552 10056 -496
rect 10112 -552 10136 -496
rect 10192 -552 10216 -496
rect 10272 -512 17626 -496
rect 10272 -552 10325 -512
rect 8855 -564 10325 -552
rect 10377 -564 10389 -512
rect 10441 -564 10453 -512
rect 10505 -564 10842 -512
rect 10894 -564 10906 -512
rect 10958 -564 10970 -512
rect 11022 -564 12519 -512
rect 12571 -564 12583 -512
rect 12635 -564 12647 -512
rect 12699 -564 13036 -512
rect 13088 -564 13100 -512
rect 13152 -564 13164 -512
rect 13216 -564 14681 -512
rect 14733 -564 14745 -512
rect 14797 -564 14809 -512
rect 14861 -564 15198 -512
rect 15250 -564 15262 -512
rect 15314 -564 15326 -512
rect 15378 -564 16875 -512
rect 16927 -564 16939 -512
rect 16991 -564 17003 -512
rect 17055 -564 17393 -512
rect 17445 -564 17457 -512
rect 17509 -564 17521 -512
rect 17573 -552 17626 -512
rect 17682 -552 17706 -496
rect 17762 -552 17786 -496
rect 17842 -552 17882 -496
rect 17573 -564 17882 -552
rect 1298 -574 17882 -564
rect 2425 -917 2725 -906
rect 7738 -917 8038 -906
rect 11142 -917 11442 -906
rect 16455 -917 16755 -906
rect 1473 -928 17707 -917
rect 1473 -936 2465 -928
rect 1473 -988 1523 -936
rect 1575 -988 1587 -936
rect 1639 -988 1651 -936
rect 1703 -988 1719 -936
rect 1771 -988 1783 -936
rect 1835 -988 1847 -936
rect 1899 -988 2009 -936
rect 2061 -988 2073 -936
rect 2125 -988 2137 -936
rect 2189 -988 2205 -936
rect 2257 -988 2269 -936
rect 2321 -988 2333 -936
rect 2385 -984 2465 -936
rect 2521 -984 2545 -928
rect 2601 -984 2625 -928
rect 2681 -936 7782 -928
rect 2681 -984 3721 -936
rect 2385 -988 3721 -984
rect 3773 -988 3785 -936
rect 3837 -988 3849 -936
rect 3901 -988 3917 -936
rect 3969 -988 3981 -936
rect 4033 -988 4045 -936
rect 4097 -988 4207 -936
rect 4259 -988 4271 -936
rect 4323 -988 4335 -936
rect 4387 -988 4403 -936
rect 4455 -988 4467 -936
rect 4519 -988 4531 -936
rect 4583 -988 5880 -936
rect 5932 -988 5944 -936
rect 5996 -988 6008 -936
rect 6060 -988 6076 -936
rect 6128 -988 6140 -936
rect 6192 -988 6204 -936
rect 6256 -988 6366 -936
rect 6418 -988 6430 -936
rect 6482 -988 6494 -936
rect 6546 -988 6562 -936
rect 6614 -988 6626 -936
rect 6678 -988 6690 -936
rect 6742 -984 7782 -936
rect 7838 -984 7862 -928
rect 7918 -984 7942 -928
rect 7998 -936 11182 -928
rect 7998 -984 8078 -936
rect 6742 -988 8078 -984
rect 8130 -988 8142 -936
rect 8194 -988 8206 -936
rect 8258 -988 8274 -936
rect 8326 -988 8338 -936
rect 8390 -988 8402 -936
rect 8454 -988 8564 -936
rect 8616 -988 8628 -936
rect 8680 -988 8692 -936
rect 8744 -988 8760 -936
rect 8812 -988 8824 -936
rect 8876 -988 8888 -936
rect 8940 -988 10240 -936
rect 10292 -988 10304 -936
rect 10356 -988 10368 -936
rect 10420 -988 10436 -936
rect 10488 -988 10500 -936
rect 10552 -988 10564 -936
rect 10616 -988 10726 -936
rect 10778 -988 10790 -936
rect 10842 -988 10854 -936
rect 10906 -988 10922 -936
rect 10974 -988 10986 -936
rect 11038 -988 11050 -936
rect 11102 -984 11182 -936
rect 11238 -984 11262 -928
rect 11318 -984 11342 -928
rect 11398 -936 16499 -928
rect 11398 -984 12438 -936
rect 11102 -988 12438 -984
rect 12490 -988 12502 -936
rect 12554 -988 12566 -936
rect 12618 -988 12634 -936
rect 12686 -988 12698 -936
rect 12750 -988 12762 -936
rect 12814 -988 12924 -936
rect 12976 -988 12988 -936
rect 13040 -988 13052 -936
rect 13104 -988 13120 -936
rect 13172 -988 13184 -936
rect 13236 -988 13248 -936
rect 13300 -988 14597 -936
rect 14649 -988 14661 -936
rect 14713 -988 14725 -936
rect 14777 -988 14793 -936
rect 14845 -988 14857 -936
rect 14909 -988 14921 -936
rect 14973 -988 15083 -936
rect 15135 -988 15147 -936
rect 15199 -988 15211 -936
rect 15263 -988 15279 -936
rect 15331 -988 15343 -936
rect 15395 -988 15407 -936
rect 15459 -984 16499 -936
rect 16555 -984 16579 -928
rect 16635 -984 16659 -928
rect 16715 -936 17707 -928
rect 16715 -984 16795 -936
rect 15459 -988 16795 -984
rect 16847 -988 16859 -936
rect 16911 -988 16923 -936
rect 16975 -988 16991 -936
rect 17043 -988 17055 -936
rect 17107 -988 17119 -936
rect 17171 -988 17281 -936
rect 17333 -988 17345 -936
rect 17397 -988 17409 -936
rect 17461 -988 17477 -936
rect 17529 -988 17541 -936
rect 17593 -988 17605 -936
rect 17657 -988 17707 -936
rect 1473 -1006 17707 -988
rect 1473 -1074 17707 -1056
rect 1473 -1126 1523 -1074
rect 1575 -1126 1587 -1074
rect 1639 -1126 1651 -1074
rect 1703 -1126 1719 -1074
rect 1771 -1126 1783 -1074
rect 1835 -1126 1847 -1074
rect 1899 -1126 2009 -1074
rect 2061 -1126 2073 -1074
rect 2125 -1126 2137 -1074
rect 2189 -1126 2205 -1074
rect 2257 -1126 2269 -1074
rect 2321 -1126 2333 -1074
rect 2385 -1126 2733 -1074
rect 2785 -1126 2797 -1074
rect 2849 -1126 2861 -1074
rect 2913 -1126 2929 -1074
rect 2981 -1126 2993 -1074
rect 3045 -1126 3057 -1074
rect 3109 -1126 3121 -1074
rect 3173 -1126 3189 -1074
rect 3241 -1126 3253 -1074
rect 3305 -1126 3317 -1074
rect 3369 -1126 3721 -1074
rect 3773 -1126 3785 -1074
rect 3837 -1126 3849 -1074
rect 3901 -1126 3917 -1074
rect 3969 -1126 3981 -1074
rect 4033 -1126 4045 -1074
rect 4097 -1126 4207 -1074
rect 4259 -1126 4271 -1074
rect 4323 -1126 4335 -1074
rect 4387 -1126 4403 -1074
rect 4455 -1126 4467 -1074
rect 4519 -1126 4531 -1074
rect 4583 -1126 5880 -1074
rect 5932 -1126 5944 -1074
rect 5996 -1126 6008 -1074
rect 6060 -1126 6076 -1074
rect 6128 -1126 6140 -1074
rect 6192 -1126 6204 -1074
rect 6256 -1126 6366 -1074
rect 6418 -1126 6430 -1074
rect 6482 -1126 6494 -1074
rect 6546 -1126 6562 -1074
rect 6614 -1126 6626 -1074
rect 6678 -1126 6690 -1074
rect 6742 -1126 7094 -1074
rect 7146 -1126 7158 -1074
rect 7210 -1126 7222 -1074
rect 7274 -1126 7290 -1074
rect 7342 -1126 7354 -1074
rect 7406 -1126 7418 -1074
rect 7470 -1126 7482 -1074
rect 7534 -1126 7550 -1074
rect 7602 -1126 7614 -1074
rect 7666 -1126 7678 -1074
rect 7730 -1126 8078 -1074
rect 8130 -1126 8142 -1074
rect 8194 -1126 8206 -1074
rect 8258 -1126 8274 -1074
rect 8326 -1126 8338 -1074
rect 8390 -1126 8402 -1074
rect 8454 -1126 8564 -1074
rect 8616 -1126 8628 -1074
rect 8680 -1126 8692 -1074
rect 8744 -1126 8760 -1074
rect 8812 -1126 8824 -1074
rect 8876 -1126 8888 -1074
rect 8940 -1126 10240 -1074
rect 10292 -1126 10304 -1074
rect 10356 -1126 10368 -1074
rect 10420 -1126 10436 -1074
rect 10488 -1126 10500 -1074
rect 10552 -1126 10564 -1074
rect 10616 -1126 10726 -1074
rect 10778 -1126 10790 -1074
rect 10842 -1126 10854 -1074
rect 10906 -1126 10922 -1074
rect 10974 -1126 10986 -1074
rect 11038 -1126 11050 -1074
rect 11102 -1126 11450 -1074
rect 11502 -1126 11514 -1074
rect 11566 -1126 11578 -1074
rect 11630 -1126 11646 -1074
rect 11698 -1126 11710 -1074
rect 11762 -1126 11774 -1074
rect 11826 -1126 11838 -1074
rect 11890 -1126 11906 -1074
rect 11958 -1126 11970 -1074
rect 12022 -1126 12034 -1074
rect 12086 -1126 12438 -1074
rect 12490 -1126 12502 -1074
rect 12554 -1126 12566 -1074
rect 12618 -1126 12634 -1074
rect 12686 -1126 12698 -1074
rect 12750 -1126 12762 -1074
rect 12814 -1126 12924 -1074
rect 12976 -1126 12988 -1074
rect 13040 -1126 13052 -1074
rect 13104 -1126 13120 -1074
rect 13172 -1126 13184 -1074
rect 13236 -1126 13248 -1074
rect 13300 -1126 14597 -1074
rect 14649 -1126 14661 -1074
rect 14713 -1126 14725 -1074
rect 14777 -1126 14793 -1074
rect 14845 -1126 14857 -1074
rect 14909 -1126 14921 -1074
rect 14973 -1126 15083 -1074
rect 15135 -1126 15147 -1074
rect 15199 -1126 15211 -1074
rect 15263 -1126 15279 -1074
rect 15331 -1126 15343 -1074
rect 15395 -1126 15407 -1074
rect 15459 -1126 15811 -1074
rect 15863 -1126 15875 -1074
rect 15927 -1126 15939 -1074
rect 15991 -1126 16007 -1074
rect 16059 -1126 16071 -1074
rect 16123 -1126 16135 -1074
rect 16187 -1126 16199 -1074
rect 16251 -1126 16267 -1074
rect 16319 -1126 16331 -1074
rect 16383 -1126 16395 -1074
rect 16447 -1126 16795 -1074
rect 16847 -1126 16859 -1074
rect 16911 -1126 16923 -1074
rect 16975 -1126 16991 -1074
rect 17043 -1126 17055 -1074
rect 17107 -1126 17119 -1074
rect 17171 -1126 17281 -1074
rect 17333 -1126 17345 -1074
rect 17397 -1126 17409 -1074
rect 17461 -1126 17477 -1074
rect 17529 -1126 17541 -1074
rect 17593 -1126 17605 -1074
rect 17657 -1126 17707 -1074
rect 1473 -1144 17707 -1126
rect 3393 -1238 3693 -1226
rect 6770 -1238 7070 -1226
rect 12110 -1238 12410 -1226
rect 15487 -1238 15787 -1226
rect 1473 -1248 17707 -1238
rect 1473 -1252 3433 -1248
rect 1473 -1304 1523 -1252
rect 1575 -1304 1587 -1252
rect 1639 -1304 1651 -1252
rect 1703 -1304 1719 -1252
rect 1771 -1304 1783 -1252
rect 1835 -1304 1847 -1252
rect 1899 -1304 2009 -1252
rect 2061 -1304 2073 -1252
rect 2125 -1304 2137 -1252
rect 2189 -1304 2205 -1252
rect 2257 -1304 2269 -1252
rect 2321 -1304 2333 -1252
rect 2385 -1304 3433 -1252
rect 3489 -1304 3513 -1248
rect 3569 -1304 3593 -1248
rect 3649 -1252 6814 -1248
rect 3649 -1304 3721 -1252
rect 3773 -1304 3785 -1252
rect 3837 -1304 3849 -1252
rect 3901 -1304 3917 -1252
rect 3969 -1304 3981 -1252
rect 4033 -1304 4045 -1252
rect 4097 -1304 4207 -1252
rect 4259 -1304 4271 -1252
rect 4323 -1304 4335 -1252
rect 4387 -1304 4403 -1252
rect 4455 -1304 4467 -1252
rect 4519 -1304 4531 -1252
rect 4583 -1304 5880 -1252
rect 5932 -1304 5944 -1252
rect 5996 -1304 6008 -1252
rect 6060 -1304 6076 -1252
rect 6128 -1304 6140 -1252
rect 6192 -1304 6204 -1252
rect 6256 -1304 6366 -1252
rect 6418 -1304 6430 -1252
rect 6482 -1304 6494 -1252
rect 6546 -1304 6562 -1252
rect 6614 -1304 6626 -1252
rect 6678 -1304 6690 -1252
rect 6742 -1304 6814 -1252
rect 6870 -1304 6894 -1248
rect 6950 -1304 6974 -1248
rect 7030 -1252 12150 -1248
rect 7030 -1304 8078 -1252
rect 8130 -1304 8142 -1252
rect 8194 -1304 8206 -1252
rect 8258 -1304 8274 -1252
rect 8326 -1304 8338 -1252
rect 8390 -1304 8402 -1252
rect 8454 -1304 8564 -1252
rect 8616 -1304 8628 -1252
rect 8680 -1304 8692 -1252
rect 8744 -1304 8760 -1252
rect 8812 -1304 8824 -1252
rect 8876 -1304 8888 -1252
rect 8940 -1304 10240 -1252
rect 10292 -1304 10304 -1252
rect 10356 -1304 10368 -1252
rect 10420 -1304 10436 -1252
rect 10488 -1304 10500 -1252
rect 10552 -1304 10564 -1252
rect 10616 -1304 10726 -1252
rect 10778 -1304 10790 -1252
rect 10842 -1304 10854 -1252
rect 10906 -1304 10922 -1252
rect 10974 -1304 10986 -1252
rect 11038 -1304 11050 -1252
rect 11102 -1304 12150 -1252
rect 12206 -1304 12230 -1248
rect 12286 -1304 12310 -1248
rect 12366 -1252 15531 -1248
rect 12366 -1304 12438 -1252
rect 12490 -1304 12502 -1252
rect 12554 -1304 12566 -1252
rect 12618 -1304 12634 -1252
rect 12686 -1304 12698 -1252
rect 12750 -1304 12762 -1252
rect 12814 -1304 12924 -1252
rect 12976 -1304 12988 -1252
rect 13040 -1304 13052 -1252
rect 13104 -1304 13120 -1252
rect 13172 -1304 13184 -1252
rect 13236 -1304 13248 -1252
rect 13300 -1304 14597 -1252
rect 14649 -1304 14661 -1252
rect 14713 -1304 14725 -1252
rect 14777 -1304 14793 -1252
rect 14845 -1304 14857 -1252
rect 14909 -1304 14921 -1252
rect 14973 -1304 15083 -1252
rect 15135 -1304 15147 -1252
rect 15199 -1304 15211 -1252
rect 15263 -1304 15279 -1252
rect 15331 -1304 15343 -1252
rect 15395 -1304 15407 -1252
rect 15459 -1304 15531 -1252
rect 15587 -1304 15611 -1248
rect 15667 -1304 15691 -1248
rect 15747 -1252 17707 -1248
rect 15747 -1304 16795 -1252
rect 16847 -1304 16859 -1252
rect 16911 -1304 16923 -1252
rect 16975 -1304 16991 -1252
rect 17043 -1304 17055 -1252
rect 17107 -1304 17119 -1252
rect 17171 -1304 17281 -1252
rect 17333 -1304 17345 -1252
rect 17397 -1304 17409 -1252
rect 17461 -1304 17477 -1252
rect 17529 -1304 17541 -1252
rect 17593 -1304 17605 -1252
rect 17657 -1304 17707 -1252
rect 1473 -1326 17707 -1304
rect 1343 -1686 17837 -1664
rect 1343 -1702 4985 -1686
rect 1343 -1754 1350 -1702
rect 1402 -1754 1414 -1702
rect 1466 -1754 1478 -1702
rect 1530 -1754 1865 -1702
rect 1917 -1754 1929 -1702
rect 1981 -1754 1993 -1702
rect 2045 -1754 2383 -1702
rect 2435 -1754 2447 -1702
rect 2499 -1754 2511 -1702
rect 2563 -1754 3543 -1702
rect 3595 -1754 3607 -1702
rect 3659 -1754 3671 -1702
rect 3723 -1754 4060 -1702
rect 4112 -1754 4124 -1702
rect 4176 -1754 4188 -1702
rect 4240 -1754 4577 -1702
rect 4629 -1754 4641 -1702
rect 4693 -1754 4705 -1702
rect 4757 -1742 4985 -1702
rect 5041 -1742 5065 -1686
rect 5121 -1742 5145 -1686
rect 5201 -1742 5262 -1686
rect 5318 -1742 5342 -1686
rect 5398 -1742 5422 -1686
rect 5478 -1702 13702 -1686
rect 5478 -1742 5706 -1702
rect 4757 -1754 5706 -1742
rect 5758 -1754 5770 -1702
rect 5822 -1754 5834 -1702
rect 5886 -1754 6223 -1702
rect 6275 -1754 6287 -1702
rect 6339 -1754 6351 -1702
rect 6403 -1754 6740 -1702
rect 6792 -1754 6804 -1702
rect 6856 -1754 6868 -1702
rect 6920 -1754 7900 -1702
rect 7952 -1754 7964 -1702
rect 8016 -1754 8028 -1702
rect 8080 -1754 8417 -1702
rect 8469 -1754 8481 -1702
rect 8533 -1754 8545 -1702
rect 8597 -1754 8932 -1702
rect 8984 -1754 8996 -1702
rect 9048 -1754 9060 -1702
rect 9112 -1754 10068 -1702
rect 10120 -1754 10132 -1702
rect 10184 -1754 10196 -1702
rect 10248 -1754 10583 -1702
rect 10635 -1754 10647 -1702
rect 10699 -1754 10711 -1702
rect 10763 -1754 11100 -1702
rect 11152 -1754 11164 -1702
rect 11216 -1754 11228 -1702
rect 11280 -1754 12260 -1702
rect 12312 -1754 12324 -1702
rect 12376 -1754 12388 -1702
rect 12440 -1754 12777 -1702
rect 12829 -1754 12841 -1702
rect 12893 -1754 12905 -1702
rect 12957 -1754 13294 -1702
rect 13346 -1754 13358 -1702
rect 13410 -1754 13422 -1702
rect 13474 -1742 13702 -1702
rect 13758 -1742 13782 -1686
rect 13838 -1742 13862 -1686
rect 13918 -1742 13979 -1686
rect 14035 -1742 14059 -1686
rect 14115 -1742 14139 -1686
rect 14195 -1702 17837 -1686
rect 14195 -1742 14423 -1702
rect 13474 -1754 14423 -1742
rect 14475 -1754 14487 -1702
rect 14539 -1754 14551 -1702
rect 14603 -1754 14940 -1702
rect 14992 -1754 15004 -1702
rect 15056 -1754 15068 -1702
rect 15120 -1754 15457 -1702
rect 15509 -1754 15521 -1702
rect 15573 -1754 15585 -1702
rect 15637 -1754 16617 -1702
rect 16669 -1754 16681 -1702
rect 16733 -1754 16745 -1702
rect 16797 -1754 17135 -1702
rect 17187 -1754 17199 -1702
rect 17251 -1754 17263 -1702
rect 17315 -1754 17650 -1702
rect 17702 -1754 17714 -1702
rect 17766 -1754 17778 -1702
rect 17830 -1754 17837 -1702
rect 1343 -1764 17837 -1754
rect 1298 -1826 17882 -1804
rect 1298 -1882 1338 -1826
rect 1394 -1882 1418 -1826
rect 1474 -1882 1498 -1826
rect 1554 -1842 8908 -1826
rect 1554 -1882 2833 -1842
rect 1298 -1894 2833 -1882
rect 2885 -1894 2897 -1842
rect 2949 -1894 2961 -1842
rect 3013 -1894 3350 -1842
rect 3402 -1894 3414 -1842
rect 3466 -1894 3478 -1842
rect 3530 -1894 6933 -1842
rect 6985 -1894 6997 -1842
rect 7049 -1894 7061 -1842
rect 7113 -1894 7450 -1842
rect 7502 -1894 7514 -1842
rect 7566 -1894 7578 -1842
rect 7630 -1882 8908 -1842
rect 8964 -1882 8988 -1826
rect 9044 -1882 9068 -1826
rect 9124 -1882 10056 -1826
rect 10112 -1882 10136 -1826
rect 10192 -1882 10216 -1826
rect 10272 -1842 17626 -1826
rect 10272 -1882 11550 -1842
rect 7630 -1894 11550 -1882
rect 11602 -1894 11614 -1842
rect 11666 -1894 11678 -1842
rect 11730 -1894 12067 -1842
rect 12119 -1894 12131 -1842
rect 12183 -1894 12195 -1842
rect 12247 -1894 15650 -1842
rect 15702 -1894 15714 -1842
rect 15766 -1894 15778 -1842
rect 15830 -1894 16167 -1842
rect 16219 -1894 16231 -1842
rect 16283 -1894 16295 -1842
rect 16347 -1882 17626 -1842
rect 17682 -1882 17706 -1826
rect 17762 -1882 17786 -1826
rect 17842 -1882 17882 -1826
rect 16347 -1894 17882 -1882
rect 1298 -1904 17882 -1894
rect 1601 -1987 17579 -1965
rect 1601 -2003 4550 -1987
rect 1601 -2055 1608 -2003
rect 1660 -2055 1672 -2003
rect 1724 -2055 1736 -2003
rect 1788 -2055 2126 -2003
rect 2178 -2055 2190 -2003
rect 2242 -2055 2254 -2003
rect 2306 -2055 3803 -2003
rect 3855 -2055 3867 -2003
rect 3919 -2055 3931 -2003
rect 3983 -2055 4320 -2003
rect 4372 -2055 4384 -2003
rect 4436 -2055 4448 -2003
rect 4500 -2043 4550 -2003
rect 4606 -2043 4630 -1987
rect 4686 -2043 4710 -1987
rect 4766 -2043 5697 -1987
rect 5753 -2043 5777 -1987
rect 5833 -2043 5857 -1987
rect 5913 -2003 13267 -1987
rect 5913 -2043 5963 -2003
rect 4500 -2055 5963 -2043
rect 6015 -2055 6027 -2003
rect 6079 -2055 6091 -2003
rect 6143 -2055 6480 -2003
rect 6532 -2055 6544 -2003
rect 6596 -2055 6608 -2003
rect 6660 -2055 8157 -2003
rect 8209 -2055 8221 -2003
rect 8273 -2055 8285 -2003
rect 8337 -2055 8674 -2003
rect 8726 -2055 8738 -2003
rect 8790 -2055 8802 -2003
rect 8854 -2055 10326 -2003
rect 10378 -2055 10390 -2003
rect 10442 -2055 10454 -2003
rect 10506 -2055 10843 -2003
rect 10895 -2055 10907 -2003
rect 10959 -2055 10971 -2003
rect 11023 -2055 12520 -2003
rect 12572 -2055 12584 -2003
rect 12636 -2055 12648 -2003
rect 12700 -2055 13037 -2003
rect 13089 -2055 13101 -2003
rect 13153 -2055 13165 -2003
rect 13217 -2043 13267 -2003
rect 13323 -2043 13347 -1987
rect 13403 -2043 13427 -1987
rect 13483 -2043 14414 -1987
rect 14470 -2043 14494 -1987
rect 14550 -2043 14574 -1987
rect 14630 -2003 17579 -1987
rect 14630 -2043 14680 -2003
rect 13217 -2055 14680 -2043
rect 14732 -2055 14744 -2003
rect 14796 -2055 14808 -2003
rect 14860 -2055 15197 -2003
rect 15249 -2055 15261 -2003
rect 15313 -2055 15325 -2003
rect 15377 -2055 16874 -2003
rect 16926 -2055 16938 -2003
rect 16990 -2055 17002 -2003
rect 17054 -2055 17392 -2003
rect 17444 -2055 17456 -2003
rect 17508 -2055 17520 -2003
rect 17572 -2055 17579 -2003
rect 1601 -2065 17579 -2055
rect 865 -2131 18315 -2109
rect 865 -2187 916 -2131
rect 972 -2187 996 -2131
rect 1052 -2187 1076 -2131
rect 1132 -2147 9331 -2131
rect 1132 -2187 2575 -2147
rect 865 -2199 2575 -2187
rect 2627 -2199 2639 -2147
rect 2691 -2199 2703 -2147
rect 2755 -2199 3092 -2147
rect 3144 -2199 3156 -2147
rect 3208 -2199 3220 -2147
rect 3272 -2199 7191 -2147
rect 7243 -2199 7255 -2147
rect 7307 -2199 7319 -2147
rect 7371 -2199 7708 -2147
rect 7760 -2199 7772 -2147
rect 7824 -2199 7836 -2147
rect 7888 -2187 9331 -2147
rect 9387 -2187 9411 -2131
rect 9467 -2187 9491 -2131
rect 9547 -2187 9633 -2131
rect 9689 -2187 9713 -2131
rect 9769 -2187 9793 -2131
rect 9849 -2147 18048 -2131
rect 9849 -2187 11292 -2147
rect 7888 -2199 11292 -2187
rect 11344 -2199 11356 -2147
rect 11408 -2199 11420 -2147
rect 11472 -2199 11809 -2147
rect 11861 -2199 11873 -2147
rect 11925 -2199 11937 -2147
rect 11989 -2199 15908 -2147
rect 15960 -2199 15972 -2147
rect 16024 -2199 16036 -2147
rect 16088 -2199 16425 -2147
rect 16477 -2199 16489 -2147
rect 16541 -2199 16553 -2147
rect 16605 -2187 18048 -2147
rect 18104 -2187 18128 -2131
rect 18184 -2187 18208 -2131
rect 18264 -2187 18315 -2131
rect 16605 -2199 18315 -2187
rect 865 -2209 18315 -2199
rect 3393 -2564 3693 -2553
rect 15487 -2564 15787 -2553
rect 1473 -2575 17707 -2564
rect 1473 -2583 3433 -2575
rect 1473 -2635 1523 -2583
rect 1575 -2635 1587 -2583
rect 1639 -2635 1651 -2583
rect 1703 -2635 1719 -2583
rect 1771 -2635 1783 -2583
rect 1835 -2635 1847 -2583
rect 1899 -2635 2009 -2583
rect 2061 -2635 2073 -2583
rect 2125 -2635 2137 -2583
rect 2189 -2635 2205 -2583
rect 2257 -2635 2269 -2583
rect 2321 -2635 2333 -2583
rect 2385 -2631 3433 -2583
rect 3489 -2631 3513 -2575
rect 3569 -2631 3593 -2575
rect 3649 -2583 15531 -2575
rect 3649 -2631 3721 -2583
rect 2385 -2635 3721 -2631
rect 3773 -2635 3785 -2583
rect 3837 -2635 3849 -2583
rect 3901 -2635 3917 -2583
rect 3969 -2635 3981 -2583
rect 4033 -2635 4045 -2583
rect 4097 -2635 4207 -2583
rect 4259 -2635 4271 -2583
rect 4323 -2635 4335 -2583
rect 4387 -2635 4403 -2583
rect 4455 -2635 4467 -2583
rect 4519 -2635 4531 -2583
rect 4583 -2635 5880 -2583
rect 5932 -2635 5944 -2583
rect 5996 -2635 6008 -2583
rect 6060 -2635 6076 -2583
rect 6128 -2635 6140 -2583
rect 6192 -2635 6204 -2583
rect 6256 -2635 6366 -2583
rect 6418 -2635 6430 -2583
rect 6482 -2635 6494 -2583
rect 6546 -2635 6562 -2583
rect 6614 -2635 6626 -2583
rect 6678 -2635 6690 -2583
rect 6742 -2586 8078 -2583
rect 6742 -2635 6814 -2586
rect 1473 -2642 6814 -2635
rect 6870 -2642 6894 -2586
rect 6950 -2642 6974 -2586
rect 7030 -2635 8078 -2586
rect 8130 -2635 8142 -2583
rect 8194 -2635 8206 -2583
rect 8258 -2635 8274 -2583
rect 8326 -2635 8338 -2583
rect 8390 -2635 8402 -2583
rect 8454 -2635 8564 -2583
rect 8616 -2635 8628 -2583
rect 8680 -2635 8692 -2583
rect 8744 -2635 8760 -2583
rect 8812 -2635 8824 -2583
rect 8876 -2635 8888 -2583
rect 8940 -2635 10240 -2583
rect 10292 -2635 10304 -2583
rect 10356 -2635 10368 -2583
rect 10420 -2635 10436 -2583
rect 10488 -2635 10500 -2583
rect 10552 -2635 10564 -2583
rect 10616 -2635 10726 -2583
rect 10778 -2635 10790 -2583
rect 10842 -2635 10854 -2583
rect 10906 -2635 10922 -2583
rect 10974 -2635 10986 -2583
rect 11038 -2635 11050 -2583
rect 11102 -2586 12438 -2583
rect 11102 -2635 12150 -2586
rect 7030 -2642 12150 -2635
rect 12206 -2642 12230 -2586
rect 12286 -2642 12310 -2586
rect 12366 -2635 12438 -2586
rect 12490 -2635 12502 -2583
rect 12554 -2635 12566 -2583
rect 12618 -2635 12634 -2583
rect 12686 -2635 12698 -2583
rect 12750 -2635 12762 -2583
rect 12814 -2635 12924 -2583
rect 12976 -2635 12988 -2583
rect 13040 -2635 13052 -2583
rect 13104 -2635 13120 -2583
rect 13172 -2635 13184 -2583
rect 13236 -2635 13248 -2583
rect 13300 -2635 14597 -2583
rect 14649 -2635 14661 -2583
rect 14713 -2635 14725 -2583
rect 14777 -2635 14793 -2583
rect 14845 -2635 14857 -2583
rect 14909 -2635 14921 -2583
rect 14973 -2635 15083 -2583
rect 15135 -2635 15147 -2583
rect 15199 -2635 15211 -2583
rect 15263 -2635 15279 -2583
rect 15331 -2635 15343 -2583
rect 15395 -2635 15407 -2583
rect 15459 -2631 15531 -2583
rect 15587 -2631 15611 -2575
rect 15667 -2631 15691 -2575
rect 15747 -2583 17707 -2575
rect 15747 -2631 16795 -2583
rect 15459 -2635 16795 -2631
rect 16847 -2635 16859 -2583
rect 16911 -2635 16923 -2583
rect 16975 -2635 16991 -2583
rect 17043 -2635 17055 -2583
rect 17107 -2635 17119 -2583
rect 17171 -2635 17281 -2583
rect 17333 -2635 17345 -2583
rect 17397 -2635 17409 -2583
rect 17461 -2635 17477 -2583
rect 17529 -2635 17541 -2583
rect 17593 -2635 17605 -2583
rect 17657 -2635 17707 -2583
rect 12366 -2642 17707 -2635
rect 1473 -2653 17707 -2642
rect 6770 -2664 7070 -2653
rect 12110 -2664 12410 -2653
rect 1473 -2721 17707 -2703
rect 1473 -2773 1523 -2721
rect 1575 -2773 1587 -2721
rect 1639 -2773 1651 -2721
rect 1703 -2773 1719 -2721
rect 1771 -2773 1783 -2721
rect 1835 -2773 1847 -2721
rect 1899 -2773 2009 -2721
rect 2061 -2773 2073 -2721
rect 2125 -2773 2137 -2721
rect 2189 -2773 2205 -2721
rect 2257 -2773 2269 -2721
rect 2321 -2773 2333 -2721
rect 2385 -2773 2733 -2721
rect 2785 -2773 2797 -2721
rect 2849 -2773 2861 -2721
rect 2913 -2773 2929 -2721
rect 2981 -2773 2993 -2721
rect 3045 -2773 3057 -2721
rect 3109 -2773 3121 -2721
rect 3173 -2773 3189 -2721
rect 3241 -2773 3253 -2721
rect 3305 -2773 3317 -2721
rect 3369 -2773 3721 -2721
rect 3773 -2773 3785 -2721
rect 3837 -2773 3849 -2721
rect 3901 -2773 3917 -2721
rect 3969 -2773 3981 -2721
rect 4033 -2773 4045 -2721
rect 4097 -2773 4207 -2721
rect 4259 -2773 4271 -2721
rect 4323 -2773 4335 -2721
rect 4387 -2773 4403 -2721
rect 4455 -2773 4467 -2721
rect 4519 -2773 4531 -2721
rect 4583 -2773 5880 -2721
rect 5932 -2773 5944 -2721
rect 5996 -2773 6008 -2721
rect 6060 -2773 6076 -2721
rect 6128 -2773 6140 -2721
rect 6192 -2773 6204 -2721
rect 6256 -2773 6366 -2721
rect 6418 -2773 6430 -2721
rect 6482 -2773 6494 -2721
rect 6546 -2773 6562 -2721
rect 6614 -2773 6626 -2721
rect 6678 -2773 6690 -2721
rect 6742 -2773 7094 -2721
rect 7146 -2773 7158 -2721
rect 7210 -2773 7222 -2721
rect 7274 -2773 7290 -2721
rect 7342 -2773 7354 -2721
rect 7406 -2773 7418 -2721
rect 7470 -2773 7482 -2721
rect 7534 -2773 7550 -2721
rect 7602 -2773 7614 -2721
rect 7666 -2773 7678 -2721
rect 7730 -2773 8078 -2721
rect 8130 -2773 8142 -2721
rect 8194 -2773 8206 -2721
rect 8258 -2773 8274 -2721
rect 8326 -2773 8338 -2721
rect 8390 -2773 8402 -2721
rect 8454 -2773 8564 -2721
rect 8616 -2773 8628 -2721
rect 8680 -2773 8692 -2721
rect 8744 -2773 8760 -2721
rect 8812 -2773 8824 -2721
rect 8876 -2773 8888 -2721
rect 8940 -2773 10240 -2721
rect 10292 -2773 10304 -2721
rect 10356 -2773 10368 -2721
rect 10420 -2773 10436 -2721
rect 10488 -2773 10500 -2721
rect 10552 -2773 10564 -2721
rect 10616 -2773 10726 -2721
rect 10778 -2773 10790 -2721
rect 10842 -2773 10854 -2721
rect 10906 -2773 10922 -2721
rect 10974 -2773 10986 -2721
rect 11038 -2773 11050 -2721
rect 11102 -2773 11450 -2721
rect 11502 -2773 11514 -2721
rect 11566 -2773 11578 -2721
rect 11630 -2773 11646 -2721
rect 11698 -2773 11710 -2721
rect 11762 -2773 11774 -2721
rect 11826 -2773 11838 -2721
rect 11890 -2773 11906 -2721
rect 11958 -2773 11970 -2721
rect 12022 -2773 12034 -2721
rect 12086 -2773 12438 -2721
rect 12490 -2773 12502 -2721
rect 12554 -2773 12566 -2721
rect 12618 -2773 12634 -2721
rect 12686 -2773 12698 -2721
rect 12750 -2773 12762 -2721
rect 12814 -2773 12924 -2721
rect 12976 -2773 12988 -2721
rect 13040 -2773 13052 -2721
rect 13104 -2773 13120 -2721
rect 13172 -2773 13184 -2721
rect 13236 -2773 13248 -2721
rect 13300 -2773 14597 -2721
rect 14649 -2773 14661 -2721
rect 14713 -2773 14725 -2721
rect 14777 -2773 14793 -2721
rect 14845 -2773 14857 -2721
rect 14909 -2773 14921 -2721
rect 14973 -2773 15083 -2721
rect 15135 -2773 15147 -2721
rect 15199 -2773 15211 -2721
rect 15263 -2773 15279 -2721
rect 15331 -2773 15343 -2721
rect 15395 -2773 15407 -2721
rect 15459 -2773 15811 -2721
rect 15863 -2773 15875 -2721
rect 15927 -2773 15939 -2721
rect 15991 -2773 16007 -2721
rect 16059 -2773 16071 -2721
rect 16123 -2773 16135 -2721
rect 16187 -2773 16199 -2721
rect 16251 -2773 16267 -2721
rect 16319 -2773 16331 -2721
rect 16383 -2773 16395 -2721
rect 16447 -2773 16795 -2721
rect 16847 -2773 16859 -2721
rect 16911 -2773 16923 -2721
rect 16975 -2773 16991 -2721
rect 17043 -2773 17055 -2721
rect 17107 -2773 17119 -2721
rect 17171 -2773 17281 -2721
rect 17333 -2773 17345 -2721
rect 17397 -2773 17409 -2721
rect 17461 -2773 17477 -2721
rect 17529 -2773 17541 -2721
rect 17593 -2773 17605 -2721
rect 17657 -2773 17707 -2721
rect 1473 -2791 17707 -2773
rect 1473 -2899 17707 -2885
rect 1473 -2951 1523 -2899
rect 1575 -2951 1587 -2899
rect 1639 -2951 1651 -2899
rect 1703 -2951 1719 -2899
rect 1771 -2951 1783 -2899
rect 1835 -2951 1847 -2899
rect 1899 -2951 2009 -2899
rect 2061 -2951 2073 -2899
rect 2125 -2951 2137 -2899
rect 2189 -2951 2205 -2899
rect 2257 -2951 2269 -2899
rect 2321 -2951 2333 -2899
rect 2385 -2907 3721 -2899
rect 2385 -2951 2465 -2907
rect 1473 -2963 2465 -2951
rect 2521 -2963 2545 -2907
rect 2601 -2963 2625 -2907
rect 2681 -2951 3721 -2907
rect 3773 -2951 3785 -2899
rect 3837 -2951 3849 -2899
rect 3901 -2951 3917 -2899
rect 3969 -2951 3981 -2899
rect 4033 -2951 4045 -2899
rect 4097 -2951 4207 -2899
rect 4259 -2951 4271 -2899
rect 4323 -2951 4335 -2899
rect 4387 -2951 4403 -2899
rect 4455 -2951 4467 -2899
rect 4519 -2951 4531 -2899
rect 4583 -2951 5880 -2899
rect 5932 -2951 5944 -2899
rect 5996 -2951 6008 -2899
rect 6060 -2951 6076 -2899
rect 6128 -2951 6140 -2899
rect 6192 -2951 6204 -2899
rect 6256 -2951 6366 -2899
rect 6418 -2951 6430 -2899
rect 6482 -2951 6494 -2899
rect 6546 -2951 6562 -2899
rect 6614 -2951 6626 -2899
rect 6678 -2951 6690 -2899
rect 6742 -2907 8078 -2899
rect 6742 -2951 7782 -2907
rect 2681 -2963 7782 -2951
rect 7838 -2963 7862 -2907
rect 7918 -2963 7942 -2907
rect 7998 -2951 8078 -2907
rect 8130 -2951 8142 -2899
rect 8194 -2951 8206 -2899
rect 8258 -2951 8274 -2899
rect 8326 -2951 8338 -2899
rect 8390 -2951 8402 -2899
rect 8454 -2951 8564 -2899
rect 8616 -2951 8628 -2899
rect 8680 -2951 8692 -2899
rect 8744 -2951 8760 -2899
rect 8812 -2951 8824 -2899
rect 8876 -2951 8888 -2899
rect 8940 -2951 10240 -2899
rect 10292 -2951 10304 -2899
rect 10356 -2951 10368 -2899
rect 10420 -2951 10436 -2899
rect 10488 -2951 10500 -2899
rect 10552 -2951 10564 -2899
rect 10616 -2951 10726 -2899
rect 10778 -2951 10790 -2899
rect 10842 -2951 10854 -2899
rect 10906 -2951 10922 -2899
rect 10974 -2951 10986 -2899
rect 11038 -2951 11050 -2899
rect 11102 -2907 12438 -2899
rect 11102 -2951 11182 -2907
rect 7998 -2963 11182 -2951
rect 11238 -2963 11262 -2907
rect 11318 -2963 11342 -2907
rect 11398 -2951 12438 -2907
rect 12490 -2951 12502 -2899
rect 12554 -2951 12566 -2899
rect 12618 -2951 12634 -2899
rect 12686 -2951 12698 -2899
rect 12750 -2951 12762 -2899
rect 12814 -2951 12924 -2899
rect 12976 -2951 12988 -2899
rect 13040 -2951 13052 -2899
rect 13104 -2951 13120 -2899
rect 13172 -2951 13184 -2899
rect 13236 -2951 13248 -2899
rect 13300 -2951 14597 -2899
rect 14649 -2951 14661 -2899
rect 14713 -2951 14725 -2899
rect 14777 -2951 14793 -2899
rect 14845 -2951 14857 -2899
rect 14909 -2951 14921 -2899
rect 14973 -2951 15083 -2899
rect 15135 -2951 15147 -2899
rect 15199 -2951 15211 -2899
rect 15263 -2951 15279 -2899
rect 15331 -2951 15343 -2899
rect 15395 -2951 15407 -2899
rect 15459 -2907 16795 -2899
rect 15459 -2951 16499 -2907
rect 11398 -2963 16499 -2951
rect 16555 -2963 16579 -2907
rect 16635 -2963 16659 -2907
rect 16715 -2951 16795 -2907
rect 16847 -2951 16859 -2899
rect 16911 -2951 16923 -2899
rect 16975 -2951 16991 -2899
rect 17043 -2951 17055 -2899
rect 17107 -2951 17119 -2899
rect 17171 -2951 17281 -2899
rect 17333 -2951 17345 -2899
rect 17397 -2951 17409 -2899
rect 17461 -2951 17477 -2899
rect 17529 -2951 17541 -2899
rect 17593 -2951 17605 -2899
rect 17657 -2951 17707 -2899
rect 16715 -2963 17707 -2951
rect 1473 -2973 17707 -2963
rect 2425 -2985 2725 -2973
rect 7738 -2985 8038 -2973
rect 11142 -2985 11442 -2973
rect 16455 -2985 16755 -2973
rect 1298 -3326 17882 -3316
rect 1298 -3338 1607 -3326
rect 1298 -3394 1338 -3338
rect 1394 -3394 1418 -3338
rect 1474 -3394 1498 -3338
rect 1554 -3378 1607 -3338
rect 1659 -3378 1671 -3326
rect 1723 -3378 1735 -3326
rect 1787 -3378 2125 -3326
rect 2177 -3378 2189 -3326
rect 2241 -3378 2253 -3326
rect 2305 -3378 3802 -3326
rect 3854 -3378 3866 -3326
rect 3918 -3378 3930 -3326
rect 3982 -3378 4319 -3326
rect 4371 -3378 4383 -3326
rect 4435 -3378 4447 -3326
rect 4499 -3378 5964 -3326
rect 6016 -3378 6028 -3326
rect 6080 -3378 6092 -3326
rect 6144 -3378 6481 -3326
rect 6533 -3378 6545 -3326
rect 6597 -3378 6609 -3326
rect 6661 -3378 8158 -3326
rect 8210 -3378 8222 -3326
rect 8274 -3378 8286 -3326
rect 8338 -3378 8675 -3326
rect 8727 -3378 8739 -3326
rect 8791 -3378 8803 -3326
rect 8855 -3338 10325 -3326
rect 8855 -3378 8908 -3338
rect 1554 -3394 8908 -3378
rect 8964 -3394 8988 -3338
rect 9044 -3394 9068 -3338
rect 9124 -3394 10056 -3338
rect 10112 -3394 10136 -3338
rect 10192 -3394 10216 -3338
rect 10272 -3378 10325 -3338
rect 10377 -3378 10389 -3326
rect 10441 -3378 10453 -3326
rect 10505 -3378 10842 -3326
rect 10894 -3378 10906 -3326
rect 10958 -3378 10970 -3326
rect 11022 -3378 12519 -3326
rect 12571 -3378 12583 -3326
rect 12635 -3378 12647 -3326
rect 12699 -3378 13036 -3326
rect 13088 -3378 13100 -3326
rect 13152 -3378 13164 -3326
rect 13216 -3378 14681 -3326
rect 14733 -3378 14745 -3326
rect 14797 -3378 14809 -3326
rect 14861 -3378 15198 -3326
rect 15250 -3378 15262 -3326
rect 15314 -3378 15326 -3326
rect 15378 -3378 16875 -3326
rect 16927 -3378 16939 -3326
rect 16991 -3378 17003 -3326
rect 17055 -3378 17393 -3326
rect 17445 -3378 17457 -3326
rect 17509 -3378 17521 -3326
rect 17573 -3338 17882 -3326
rect 17573 -3378 17626 -3338
rect 10272 -3394 17626 -3378
rect 17682 -3394 17706 -3338
rect 17762 -3394 17786 -3338
rect 17842 -3394 17882 -3338
rect 1298 -3416 17882 -3394
rect 2570 -3495 16610 -3485
rect 2570 -3547 2577 -3495
rect 2629 -3547 2641 -3495
rect 2693 -3547 2705 -3495
rect 2757 -3547 3094 -3495
rect 3146 -3547 3158 -3495
rect 3210 -3547 3222 -3495
rect 3274 -3507 7189 -3495
rect 3274 -3547 4550 -3507
rect 2570 -3563 4550 -3547
rect 4606 -3563 4630 -3507
rect 4686 -3563 4710 -3507
rect 4766 -3563 5697 -3507
rect 5753 -3563 5777 -3507
rect 5833 -3563 5857 -3507
rect 5913 -3547 7189 -3507
rect 7241 -3547 7253 -3495
rect 7305 -3547 7317 -3495
rect 7369 -3547 7706 -3495
rect 7758 -3547 7770 -3495
rect 7822 -3547 7834 -3495
rect 7886 -3547 11294 -3495
rect 11346 -3547 11358 -3495
rect 11410 -3547 11422 -3495
rect 11474 -3547 11811 -3495
rect 11863 -3547 11875 -3495
rect 11927 -3547 11939 -3495
rect 11991 -3507 15906 -3495
rect 11991 -3547 13267 -3507
rect 5913 -3563 13267 -3547
rect 13323 -3563 13347 -3507
rect 13403 -3563 13427 -3507
rect 13483 -3563 14414 -3507
rect 14470 -3563 14494 -3507
rect 14550 -3563 14574 -3507
rect 14630 -3547 15906 -3507
rect 15958 -3547 15970 -3495
rect 16022 -3547 16034 -3495
rect 16086 -3547 16423 -3495
rect 16475 -3547 16487 -3495
rect 16539 -3547 16551 -3495
rect 16603 -3547 16610 -3495
rect 14630 -3563 16610 -3547
rect 2570 -3585 16610 -3563
rect 876 -3657 18304 -3647
rect 876 -3669 1348 -3657
rect 876 -3725 916 -3669
rect 972 -3725 996 -3669
rect 1052 -3725 1076 -3669
rect 1132 -3709 1348 -3669
rect 1400 -3709 1412 -3657
rect 1464 -3709 1476 -3657
rect 1528 -3709 1865 -3657
rect 1917 -3709 1929 -3657
rect 1981 -3709 1993 -3657
rect 2045 -3709 2382 -3657
rect 2434 -3709 2446 -3657
rect 2498 -3709 2510 -3657
rect 2562 -3709 3543 -3657
rect 3595 -3709 3607 -3657
rect 3659 -3709 3671 -3657
rect 3723 -3709 4060 -3657
rect 4112 -3709 4124 -3657
rect 4176 -3709 4188 -3657
rect 4240 -3709 4575 -3657
rect 4627 -3709 4639 -3657
rect 4691 -3709 4703 -3657
rect 4755 -3709 5708 -3657
rect 5760 -3709 5772 -3657
rect 5824 -3709 5836 -3657
rect 5888 -3709 6223 -3657
rect 6275 -3709 6287 -3657
rect 6339 -3709 6351 -3657
rect 6403 -3709 6740 -3657
rect 6792 -3709 6804 -3657
rect 6856 -3709 6868 -3657
rect 6920 -3709 7901 -3657
rect 7953 -3709 7965 -3657
rect 8017 -3709 8029 -3657
rect 8081 -3709 8417 -3657
rect 8469 -3709 8481 -3657
rect 8533 -3709 8545 -3657
rect 8597 -3709 8935 -3657
rect 8987 -3709 8999 -3657
rect 9051 -3709 9063 -3657
rect 9115 -3669 10065 -3657
rect 9115 -3709 9331 -3669
rect 1132 -3725 9331 -3709
rect 9387 -3725 9411 -3669
rect 9467 -3725 9491 -3669
rect 9547 -3725 9633 -3669
rect 9689 -3725 9713 -3669
rect 9769 -3725 9793 -3669
rect 9849 -3709 10065 -3669
rect 10117 -3709 10129 -3657
rect 10181 -3709 10193 -3657
rect 10245 -3709 10583 -3657
rect 10635 -3709 10647 -3657
rect 10699 -3709 10711 -3657
rect 10763 -3709 11099 -3657
rect 11151 -3709 11163 -3657
rect 11215 -3709 11227 -3657
rect 11279 -3709 12260 -3657
rect 12312 -3709 12324 -3657
rect 12376 -3709 12388 -3657
rect 12440 -3709 12777 -3657
rect 12829 -3709 12841 -3657
rect 12893 -3709 12905 -3657
rect 12957 -3709 13292 -3657
rect 13344 -3709 13356 -3657
rect 13408 -3709 13420 -3657
rect 13472 -3709 14425 -3657
rect 14477 -3709 14489 -3657
rect 14541 -3709 14553 -3657
rect 14605 -3709 14940 -3657
rect 14992 -3709 15004 -3657
rect 15056 -3709 15068 -3657
rect 15120 -3709 15457 -3657
rect 15509 -3709 15521 -3657
rect 15573 -3709 15585 -3657
rect 15637 -3709 16618 -3657
rect 16670 -3709 16682 -3657
rect 16734 -3709 16746 -3657
rect 16798 -3709 17135 -3657
rect 17187 -3709 17199 -3657
rect 17251 -3709 17263 -3657
rect 17315 -3709 17652 -3657
rect 17704 -3709 17716 -3657
rect 17768 -3709 17780 -3657
rect 17832 -3669 18304 -3657
rect 17832 -3709 18048 -3669
rect 9849 -3725 18048 -3709
rect 18104 -3725 18128 -3669
rect 18184 -3725 18208 -3669
rect 18264 -3725 18304 -3669
rect 876 -3747 18304 -3725
rect 2827 -3826 16353 -3816
rect 2827 -3878 2834 -3826
rect 2886 -3878 2898 -3826
rect 2950 -3878 2962 -3826
rect 3014 -3878 3351 -3826
rect 3403 -3878 3415 -3826
rect 3467 -3878 3479 -3826
rect 3531 -3838 6931 -3826
rect 3531 -3878 4985 -3838
rect 2827 -3894 4985 -3878
rect 5041 -3894 5065 -3838
rect 5121 -3894 5145 -3838
rect 5201 -3894 5262 -3838
rect 5318 -3894 5342 -3838
rect 5398 -3894 5422 -3838
rect 5478 -3878 6931 -3838
rect 6983 -3878 6995 -3826
rect 7047 -3878 7059 -3826
rect 7111 -3878 7449 -3826
rect 7501 -3878 7513 -3826
rect 7565 -3878 7577 -3826
rect 7629 -3878 11551 -3826
rect 11603 -3878 11615 -3826
rect 11667 -3878 11679 -3826
rect 11731 -3878 12069 -3826
rect 12121 -3878 12133 -3826
rect 12185 -3878 12197 -3826
rect 12249 -3838 15649 -3826
rect 12249 -3878 13702 -3838
rect 5478 -3894 13702 -3878
rect 13758 -3894 13782 -3838
rect 13838 -3894 13862 -3838
rect 13918 -3894 13979 -3838
rect 14035 -3894 14059 -3838
rect 14115 -3894 14139 -3838
rect 14195 -3878 15649 -3838
rect 15701 -3878 15713 -3826
rect 15765 -3878 15777 -3826
rect 15829 -3878 16166 -3826
rect 16218 -3878 16230 -3826
rect 16282 -3878 16294 -3826
rect 16346 -3878 16353 -3826
rect 14195 -3894 16353 -3878
rect 2827 -3916 16353 -3894
rect 2827 -4869 16353 -4847
rect 2827 -4885 4985 -4869
rect 2827 -4937 2834 -4885
rect 2886 -4937 2898 -4885
rect 2950 -4937 2962 -4885
rect 3014 -4937 3351 -4885
rect 3403 -4937 3415 -4885
rect 3467 -4937 3479 -4885
rect 3531 -4925 4985 -4885
rect 5041 -4925 5065 -4869
rect 5121 -4925 5145 -4869
rect 5201 -4925 5262 -4869
rect 5318 -4925 5342 -4869
rect 5398 -4925 5422 -4869
rect 5478 -4885 13702 -4869
rect 5478 -4925 6931 -4885
rect 3531 -4937 6931 -4925
rect 6983 -4937 6995 -4885
rect 7047 -4937 7059 -4885
rect 7111 -4937 7449 -4885
rect 7501 -4937 7513 -4885
rect 7565 -4937 7577 -4885
rect 7629 -4937 11551 -4885
rect 11603 -4937 11615 -4885
rect 11667 -4937 11679 -4885
rect 11731 -4937 12069 -4885
rect 12121 -4937 12133 -4885
rect 12185 -4937 12197 -4885
rect 12249 -4925 13702 -4885
rect 13758 -4925 13782 -4869
rect 13838 -4925 13862 -4869
rect 13918 -4925 13979 -4869
rect 14035 -4925 14059 -4869
rect 14115 -4925 14139 -4869
rect 14195 -4885 16353 -4869
rect 14195 -4925 15649 -4885
rect 12249 -4937 15649 -4925
rect 15701 -4937 15713 -4885
rect 15765 -4937 15777 -4885
rect 15829 -4937 16166 -4885
rect 16218 -4937 16230 -4885
rect 16282 -4937 16294 -4885
rect 16346 -4937 16353 -4885
rect 2827 -4947 16353 -4937
rect 876 -5038 18304 -5016
rect 876 -5094 916 -5038
rect 972 -5094 996 -5038
rect 1052 -5094 1076 -5038
rect 1132 -5054 9331 -5038
rect 1132 -5094 1348 -5054
rect 876 -5106 1348 -5094
rect 1400 -5106 1412 -5054
rect 1464 -5106 1476 -5054
rect 1528 -5106 1865 -5054
rect 1917 -5106 1929 -5054
rect 1981 -5106 1993 -5054
rect 2045 -5106 2382 -5054
rect 2434 -5106 2446 -5054
rect 2498 -5106 2510 -5054
rect 2562 -5106 3543 -5054
rect 3595 -5106 3607 -5054
rect 3659 -5106 3671 -5054
rect 3723 -5106 4060 -5054
rect 4112 -5106 4124 -5054
rect 4176 -5106 4188 -5054
rect 4240 -5106 4575 -5054
rect 4627 -5106 4639 -5054
rect 4691 -5106 4703 -5054
rect 4755 -5106 5708 -5054
rect 5760 -5106 5772 -5054
rect 5824 -5106 5836 -5054
rect 5888 -5106 6223 -5054
rect 6275 -5106 6287 -5054
rect 6339 -5106 6351 -5054
rect 6403 -5106 6740 -5054
rect 6792 -5106 6804 -5054
rect 6856 -5106 6868 -5054
rect 6920 -5106 7901 -5054
rect 7953 -5106 7965 -5054
rect 8017 -5106 8029 -5054
rect 8081 -5106 8417 -5054
rect 8469 -5106 8481 -5054
rect 8533 -5106 8545 -5054
rect 8597 -5106 8935 -5054
rect 8987 -5106 8999 -5054
rect 9051 -5106 9063 -5054
rect 9115 -5094 9331 -5054
rect 9387 -5094 9411 -5038
rect 9467 -5094 9491 -5038
rect 9547 -5094 9633 -5038
rect 9689 -5094 9713 -5038
rect 9769 -5094 9793 -5038
rect 9849 -5054 18048 -5038
rect 9849 -5094 10065 -5054
rect 9115 -5106 10065 -5094
rect 10117 -5106 10129 -5054
rect 10181 -5106 10193 -5054
rect 10245 -5106 10583 -5054
rect 10635 -5106 10647 -5054
rect 10699 -5106 10711 -5054
rect 10763 -5106 11099 -5054
rect 11151 -5106 11163 -5054
rect 11215 -5106 11227 -5054
rect 11279 -5106 12260 -5054
rect 12312 -5106 12324 -5054
rect 12376 -5106 12388 -5054
rect 12440 -5106 12777 -5054
rect 12829 -5106 12841 -5054
rect 12893 -5106 12905 -5054
rect 12957 -5106 13292 -5054
rect 13344 -5106 13356 -5054
rect 13408 -5106 13420 -5054
rect 13472 -5106 14425 -5054
rect 14477 -5106 14489 -5054
rect 14541 -5106 14553 -5054
rect 14605 -5106 14940 -5054
rect 14992 -5106 15004 -5054
rect 15056 -5106 15068 -5054
rect 15120 -5106 15457 -5054
rect 15509 -5106 15521 -5054
rect 15573 -5106 15585 -5054
rect 15637 -5106 16618 -5054
rect 16670 -5106 16682 -5054
rect 16734 -5106 16746 -5054
rect 16798 -5106 17135 -5054
rect 17187 -5106 17199 -5054
rect 17251 -5106 17263 -5054
rect 17315 -5106 17652 -5054
rect 17704 -5106 17716 -5054
rect 17768 -5106 17780 -5054
rect 17832 -5094 18048 -5054
rect 18104 -5094 18128 -5038
rect 18184 -5094 18208 -5038
rect 18264 -5094 18304 -5038
rect 17832 -5106 18304 -5094
rect 876 -5116 18304 -5106
rect 2570 -5201 16610 -5179
rect 2570 -5217 4550 -5201
rect 2570 -5269 2577 -5217
rect 2629 -5269 2641 -5217
rect 2693 -5269 2705 -5217
rect 2757 -5269 3094 -5217
rect 3146 -5269 3158 -5217
rect 3210 -5269 3222 -5217
rect 3274 -5257 4550 -5217
rect 4606 -5257 4630 -5201
rect 4686 -5257 4710 -5201
rect 4766 -5257 5697 -5201
rect 5753 -5257 5777 -5201
rect 5833 -5257 5857 -5201
rect 5913 -5217 13267 -5201
rect 5913 -5257 7189 -5217
rect 3274 -5269 7189 -5257
rect 7241 -5269 7253 -5217
rect 7305 -5269 7317 -5217
rect 7369 -5269 7706 -5217
rect 7758 -5269 7770 -5217
rect 7822 -5269 7834 -5217
rect 7886 -5269 11294 -5217
rect 11346 -5269 11358 -5217
rect 11410 -5269 11422 -5217
rect 11474 -5269 11811 -5217
rect 11863 -5269 11875 -5217
rect 11927 -5269 11939 -5217
rect 11991 -5257 13267 -5217
rect 13323 -5257 13347 -5201
rect 13403 -5257 13427 -5201
rect 13483 -5257 14414 -5201
rect 14470 -5257 14494 -5201
rect 14550 -5257 14574 -5201
rect 14630 -5217 16610 -5201
rect 14630 -5257 15906 -5217
rect 11991 -5269 15906 -5257
rect 15958 -5269 15970 -5217
rect 16022 -5269 16034 -5217
rect 16086 -5269 16423 -5217
rect 16475 -5269 16487 -5217
rect 16539 -5269 16551 -5217
rect 16603 -5269 16610 -5217
rect 2570 -5279 16610 -5269
rect 1298 -5370 17882 -5348
rect 1298 -5426 1338 -5370
rect 1394 -5426 1418 -5370
rect 1474 -5426 1498 -5370
rect 1554 -5386 8908 -5370
rect 1554 -5426 1607 -5386
rect 1298 -5438 1607 -5426
rect 1659 -5438 1671 -5386
rect 1723 -5438 1735 -5386
rect 1787 -5438 2125 -5386
rect 2177 -5438 2189 -5386
rect 2241 -5438 2253 -5386
rect 2305 -5438 3802 -5386
rect 3854 -5438 3866 -5386
rect 3918 -5438 3930 -5386
rect 3982 -5438 4319 -5386
rect 4371 -5438 4383 -5386
rect 4435 -5438 4447 -5386
rect 4499 -5438 5964 -5386
rect 6016 -5438 6028 -5386
rect 6080 -5438 6092 -5386
rect 6144 -5438 6481 -5386
rect 6533 -5438 6545 -5386
rect 6597 -5438 6609 -5386
rect 6661 -5438 8158 -5386
rect 8210 -5438 8222 -5386
rect 8274 -5438 8286 -5386
rect 8338 -5438 8675 -5386
rect 8727 -5438 8739 -5386
rect 8791 -5438 8803 -5386
rect 8855 -5426 8908 -5386
rect 8964 -5426 8988 -5370
rect 9044 -5426 9068 -5370
rect 9124 -5426 10056 -5370
rect 10112 -5426 10136 -5370
rect 10192 -5426 10216 -5370
rect 10272 -5386 17626 -5370
rect 10272 -5426 10325 -5386
rect 8855 -5438 10325 -5426
rect 10377 -5438 10389 -5386
rect 10441 -5438 10453 -5386
rect 10505 -5438 10842 -5386
rect 10894 -5438 10906 -5386
rect 10958 -5438 10970 -5386
rect 11022 -5438 12519 -5386
rect 12571 -5438 12583 -5386
rect 12635 -5438 12647 -5386
rect 12699 -5438 13036 -5386
rect 13088 -5438 13100 -5386
rect 13152 -5438 13164 -5386
rect 13216 -5438 14681 -5386
rect 14733 -5438 14745 -5386
rect 14797 -5438 14809 -5386
rect 14861 -5438 15198 -5386
rect 15250 -5438 15262 -5386
rect 15314 -5438 15326 -5386
rect 15378 -5438 16875 -5386
rect 16927 -5438 16939 -5386
rect 16991 -5438 17003 -5386
rect 17055 -5438 17393 -5386
rect 17445 -5438 17457 -5386
rect 17509 -5438 17521 -5386
rect 17573 -5426 17626 -5386
rect 17682 -5426 17706 -5370
rect 17762 -5426 17786 -5370
rect 17842 -5426 17882 -5370
rect 17573 -5438 17882 -5426
rect 1298 -5448 17882 -5438
rect 2425 -5791 2725 -5779
rect 7738 -5791 8038 -5779
rect 11142 -5791 11442 -5779
rect 16455 -5791 16755 -5779
rect 1473 -5801 17707 -5791
rect 1473 -5812 2465 -5801
rect 1473 -5864 1523 -5812
rect 1575 -5864 1587 -5812
rect 1639 -5864 1651 -5812
rect 1703 -5864 1719 -5812
rect 1771 -5864 1783 -5812
rect 1835 -5864 1847 -5812
rect 1899 -5864 2009 -5812
rect 2061 -5864 2073 -5812
rect 2125 -5864 2137 -5812
rect 2189 -5864 2205 -5812
rect 2257 -5864 2269 -5812
rect 2321 -5864 2333 -5812
rect 2385 -5857 2465 -5812
rect 2521 -5857 2545 -5801
rect 2601 -5857 2625 -5801
rect 2681 -5812 7782 -5801
rect 2681 -5857 3721 -5812
rect 2385 -5864 3721 -5857
rect 3773 -5864 3785 -5812
rect 3837 -5864 3849 -5812
rect 3901 -5864 3917 -5812
rect 3969 -5864 3981 -5812
rect 4033 -5864 4045 -5812
rect 4097 -5864 4207 -5812
rect 4259 -5864 4271 -5812
rect 4323 -5864 4335 -5812
rect 4387 -5864 4403 -5812
rect 4455 -5864 4467 -5812
rect 4519 -5864 4531 -5812
rect 4583 -5864 5880 -5812
rect 5932 -5864 5944 -5812
rect 5996 -5864 6008 -5812
rect 6060 -5864 6076 -5812
rect 6128 -5864 6140 -5812
rect 6192 -5864 6204 -5812
rect 6256 -5864 6366 -5812
rect 6418 -5864 6430 -5812
rect 6482 -5864 6494 -5812
rect 6546 -5864 6562 -5812
rect 6614 -5864 6626 -5812
rect 6678 -5864 6690 -5812
rect 6742 -5857 7782 -5812
rect 7838 -5857 7862 -5801
rect 7918 -5857 7942 -5801
rect 7998 -5812 11182 -5801
rect 7998 -5857 8078 -5812
rect 6742 -5864 8078 -5857
rect 8130 -5864 8142 -5812
rect 8194 -5864 8206 -5812
rect 8258 -5864 8274 -5812
rect 8326 -5864 8338 -5812
rect 8390 -5864 8402 -5812
rect 8454 -5864 8564 -5812
rect 8616 -5864 8628 -5812
rect 8680 -5864 8692 -5812
rect 8744 -5864 8760 -5812
rect 8812 -5864 8824 -5812
rect 8876 -5864 8888 -5812
rect 8940 -5864 10240 -5812
rect 10292 -5864 10304 -5812
rect 10356 -5864 10368 -5812
rect 10420 -5864 10436 -5812
rect 10488 -5864 10500 -5812
rect 10552 -5864 10564 -5812
rect 10616 -5864 10726 -5812
rect 10778 -5864 10790 -5812
rect 10842 -5864 10854 -5812
rect 10906 -5864 10922 -5812
rect 10974 -5864 10986 -5812
rect 11038 -5864 11050 -5812
rect 11102 -5857 11182 -5812
rect 11238 -5857 11262 -5801
rect 11318 -5857 11342 -5801
rect 11398 -5812 16499 -5801
rect 11398 -5857 12438 -5812
rect 11102 -5864 12438 -5857
rect 12490 -5864 12502 -5812
rect 12554 -5864 12566 -5812
rect 12618 -5864 12634 -5812
rect 12686 -5864 12698 -5812
rect 12750 -5864 12762 -5812
rect 12814 -5864 12924 -5812
rect 12976 -5864 12988 -5812
rect 13040 -5864 13052 -5812
rect 13104 -5864 13120 -5812
rect 13172 -5864 13184 -5812
rect 13236 -5864 13248 -5812
rect 13300 -5864 14597 -5812
rect 14649 -5864 14661 -5812
rect 14713 -5864 14725 -5812
rect 14777 -5864 14793 -5812
rect 14845 -5864 14857 -5812
rect 14909 -5864 14921 -5812
rect 14973 -5864 15083 -5812
rect 15135 -5864 15147 -5812
rect 15199 -5864 15211 -5812
rect 15263 -5864 15279 -5812
rect 15331 -5864 15343 -5812
rect 15395 -5864 15407 -5812
rect 15459 -5857 16499 -5812
rect 16555 -5857 16579 -5801
rect 16635 -5857 16659 -5801
rect 16715 -5812 17707 -5801
rect 16715 -5857 16795 -5812
rect 15459 -5864 16795 -5857
rect 16847 -5864 16859 -5812
rect 16911 -5864 16923 -5812
rect 16975 -5864 16991 -5812
rect 17043 -5864 17055 -5812
rect 17107 -5864 17119 -5812
rect 17171 -5864 17281 -5812
rect 17333 -5864 17345 -5812
rect 17397 -5864 17409 -5812
rect 17461 -5864 17477 -5812
rect 17529 -5864 17541 -5812
rect 17593 -5864 17605 -5812
rect 17657 -5864 17707 -5812
rect 1473 -5879 17707 -5864
rect 1473 -5990 17707 -5973
rect 1473 -6042 1523 -5990
rect 1575 -6042 1587 -5990
rect 1639 -6042 1651 -5990
rect 1703 -6042 1719 -5990
rect 1771 -6042 1783 -5990
rect 1835 -6042 1847 -5990
rect 1899 -6042 2009 -5990
rect 2061 -6042 2073 -5990
rect 2125 -6042 2137 -5990
rect 2189 -6042 2205 -5990
rect 2257 -6042 2269 -5990
rect 2321 -6042 2333 -5990
rect 2385 -6042 2733 -5990
rect 2785 -6042 2797 -5990
rect 2849 -6042 2861 -5990
rect 2913 -6042 2929 -5990
rect 2981 -6042 2993 -5990
rect 3045 -6042 3057 -5990
rect 3109 -6042 3121 -5990
rect 3173 -6042 3189 -5990
rect 3241 -6042 3253 -5990
rect 3305 -6042 3317 -5990
rect 3369 -6042 3721 -5990
rect 3773 -6042 3785 -5990
rect 3837 -6042 3849 -5990
rect 3901 -6042 3917 -5990
rect 3969 -6042 3981 -5990
rect 4033 -6042 4045 -5990
rect 4097 -6042 4207 -5990
rect 4259 -6042 4271 -5990
rect 4323 -6042 4335 -5990
rect 4387 -6042 4403 -5990
rect 4455 -6042 4467 -5990
rect 4519 -6042 4531 -5990
rect 4583 -6042 5880 -5990
rect 5932 -6042 5944 -5990
rect 5996 -6042 6008 -5990
rect 6060 -6042 6076 -5990
rect 6128 -6042 6140 -5990
rect 6192 -6042 6204 -5990
rect 6256 -6042 6366 -5990
rect 6418 -6042 6430 -5990
rect 6482 -6042 6494 -5990
rect 6546 -6042 6562 -5990
rect 6614 -6042 6626 -5990
rect 6678 -6042 6690 -5990
rect 6742 -6042 7094 -5990
rect 7146 -6042 7158 -5990
rect 7210 -6042 7222 -5990
rect 7274 -6042 7290 -5990
rect 7342 -6042 7354 -5990
rect 7406 -6042 7418 -5990
rect 7470 -6042 7482 -5990
rect 7534 -6042 7550 -5990
rect 7602 -6042 7614 -5990
rect 7666 -6042 7678 -5990
rect 7730 -6042 8078 -5990
rect 8130 -6042 8142 -5990
rect 8194 -6042 8206 -5990
rect 8258 -6042 8274 -5990
rect 8326 -6042 8338 -5990
rect 8390 -6042 8402 -5990
rect 8454 -6042 8564 -5990
rect 8616 -6042 8628 -5990
rect 8680 -6042 8692 -5990
rect 8744 -6042 8760 -5990
rect 8812 -6042 8824 -5990
rect 8876 -6042 8888 -5990
rect 8940 -6042 10240 -5990
rect 10292 -6042 10304 -5990
rect 10356 -6042 10368 -5990
rect 10420 -6042 10436 -5990
rect 10488 -6042 10500 -5990
rect 10552 -6042 10564 -5990
rect 10616 -6042 10726 -5990
rect 10778 -6042 10790 -5990
rect 10842 -6042 10854 -5990
rect 10906 -6042 10922 -5990
rect 10974 -6042 10986 -5990
rect 11038 -6042 11050 -5990
rect 11102 -6042 11450 -5990
rect 11502 -6042 11514 -5990
rect 11566 -6042 11578 -5990
rect 11630 -6042 11646 -5990
rect 11698 -6042 11710 -5990
rect 11762 -6042 11774 -5990
rect 11826 -6042 11838 -5990
rect 11890 -6042 11906 -5990
rect 11958 -6042 11970 -5990
rect 12022 -6042 12034 -5990
rect 12086 -6042 12438 -5990
rect 12490 -6042 12502 -5990
rect 12554 -6042 12566 -5990
rect 12618 -6042 12634 -5990
rect 12686 -6042 12698 -5990
rect 12750 -6042 12762 -5990
rect 12814 -6042 12924 -5990
rect 12976 -6042 12988 -5990
rect 13040 -6042 13052 -5990
rect 13104 -6042 13120 -5990
rect 13172 -6042 13184 -5990
rect 13236 -6042 13248 -5990
rect 13300 -6042 14597 -5990
rect 14649 -6042 14661 -5990
rect 14713 -6042 14725 -5990
rect 14777 -6042 14793 -5990
rect 14845 -6042 14857 -5990
rect 14909 -6042 14921 -5990
rect 14973 -6042 15083 -5990
rect 15135 -6042 15147 -5990
rect 15199 -6042 15211 -5990
rect 15263 -6042 15279 -5990
rect 15331 -6042 15343 -5990
rect 15395 -6042 15407 -5990
rect 15459 -6042 15811 -5990
rect 15863 -6042 15875 -5990
rect 15927 -6042 15939 -5990
rect 15991 -6042 16007 -5990
rect 16059 -6042 16071 -5990
rect 16123 -6042 16135 -5990
rect 16187 -6042 16199 -5990
rect 16251 -6042 16267 -5990
rect 16319 -6042 16331 -5990
rect 16383 -6042 16395 -5990
rect 16447 -6042 16795 -5990
rect 16847 -6042 16859 -5990
rect 16911 -6042 16923 -5990
rect 16975 -6042 16991 -5990
rect 17043 -6042 17055 -5990
rect 17107 -6042 17119 -5990
rect 17171 -6042 17281 -5990
rect 17333 -6042 17345 -5990
rect 17397 -6042 17409 -5990
rect 17461 -6042 17477 -5990
rect 17529 -6042 17541 -5990
rect 17593 -6042 17605 -5990
rect 17657 -6042 17707 -5990
rect 1473 -6061 17707 -6042
rect 1473 -6129 17707 -6111
rect 1473 -6181 1523 -6129
rect 1575 -6181 1587 -6129
rect 1639 -6181 1651 -6129
rect 1703 -6181 1719 -6129
rect 1771 -6181 1783 -6129
rect 1835 -6181 1847 -6129
rect 1899 -6181 2009 -6129
rect 2061 -6181 2073 -6129
rect 2125 -6181 2137 -6129
rect 2189 -6181 2205 -6129
rect 2257 -6181 2269 -6129
rect 2321 -6181 2333 -6129
rect 2385 -6133 3721 -6129
rect 2385 -6181 3433 -6133
rect 1473 -6189 3433 -6181
rect 3489 -6189 3513 -6133
rect 3569 -6189 3593 -6133
rect 3649 -6181 3721 -6133
rect 3773 -6181 3785 -6129
rect 3837 -6181 3849 -6129
rect 3901 -6181 3917 -6129
rect 3969 -6181 3981 -6129
rect 4033 -6181 4045 -6129
rect 4097 -6181 4207 -6129
rect 4259 -6181 4271 -6129
rect 4323 -6181 4335 -6129
rect 4387 -6181 4403 -6129
rect 4455 -6181 4467 -6129
rect 4519 -6181 4531 -6129
rect 4583 -6181 5880 -6129
rect 5932 -6181 5944 -6129
rect 5996 -6181 6008 -6129
rect 6060 -6181 6076 -6129
rect 6128 -6181 6140 -6129
rect 6192 -6181 6204 -6129
rect 6256 -6181 6366 -6129
rect 6418 -6181 6430 -6129
rect 6482 -6181 6494 -6129
rect 6546 -6181 6562 -6129
rect 6614 -6181 6626 -6129
rect 6678 -6181 6690 -6129
rect 6742 -6133 8078 -6129
rect 6742 -6181 6814 -6133
rect 3649 -6189 6814 -6181
rect 6870 -6189 6894 -6133
rect 6950 -6189 6974 -6133
rect 7030 -6181 8078 -6133
rect 8130 -6181 8142 -6129
rect 8194 -6181 8206 -6129
rect 8258 -6181 8274 -6129
rect 8326 -6181 8338 -6129
rect 8390 -6181 8402 -6129
rect 8454 -6181 8564 -6129
rect 8616 -6181 8628 -6129
rect 8680 -6181 8692 -6129
rect 8744 -6181 8760 -6129
rect 8812 -6181 8824 -6129
rect 8876 -6181 8888 -6129
rect 8940 -6181 10240 -6129
rect 10292 -6181 10304 -6129
rect 10356 -6181 10368 -6129
rect 10420 -6181 10436 -6129
rect 10488 -6181 10500 -6129
rect 10552 -6181 10564 -6129
rect 10616 -6181 10726 -6129
rect 10778 -6181 10790 -6129
rect 10842 -6181 10854 -6129
rect 10906 -6181 10922 -6129
rect 10974 -6181 10986 -6129
rect 11038 -6181 11050 -6129
rect 11102 -6133 12438 -6129
rect 11102 -6181 12150 -6133
rect 7030 -6189 12150 -6181
rect 12206 -6189 12230 -6133
rect 12286 -6189 12310 -6133
rect 12366 -6181 12438 -6133
rect 12490 -6181 12502 -6129
rect 12554 -6181 12566 -6129
rect 12618 -6181 12634 -6129
rect 12686 -6181 12698 -6129
rect 12750 -6181 12762 -6129
rect 12814 -6181 12924 -6129
rect 12976 -6181 12988 -6129
rect 13040 -6181 13052 -6129
rect 13104 -6181 13120 -6129
rect 13172 -6181 13184 -6129
rect 13236 -6181 13248 -6129
rect 13300 -6181 14597 -6129
rect 14649 -6181 14661 -6129
rect 14713 -6181 14725 -6129
rect 14777 -6181 14793 -6129
rect 14845 -6181 14857 -6129
rect 14909 -6181 14921 -6129
rect 14973 -6181 15083 -6129
rect 15135 -6181 15147 -6129
rect 15199 -6181 15211 -6129
rect 15263 -6181 15279 -6129
rect 15331 -6181 15343 -6129
rect 15395 -6181 15407 -6129
rect 15459 -6133 16795 -6129
rect 15459 -6181 15531 -6133
rect 12366 -6189 15531 -6181
rect 15587 -6189 15611 -6133
rect 15667 -6189 15691 -6133
rect 15747 -6181 16795 -6133
rect 16847 -6181 16859 -6129
rect 16911 -6181 16923 -6129
rect 16975 -6181 16991 -6129
rect 17043 -6181 17055 -6129
rect 17107 -6181 17119 -6129
rect 17171 -6181 17281 -6129
rect 17333 -6181 17345 -6129
rect 17397 -6181 17409 -6129
rect 17461 -6181 17477 -6129
rect 17529 -6181 17541 -6129
rect 17593 -6181 17605 -6129
rect 17657 -6181 17707 -6129
rect 15747 -6189 17707 -6181
rect 1473 -6199 17707 -6189
rect 3393 -6211 3693 -6199
rect 6770 -6211 7070 -6199
rect 12110 -6211 12410 -6199
rect 15487 -6211 15787 -6199
rect 865 -6564 18315 -6554
rect 865 -6576 2575 -6564
rect 865 -6632 916 -6576
rect 972 -6632 996 -6576
rect 1052 -6632 1076 -6576
rect 1132 -6616 2575 -6576
rect 2627 -6616 2639 -6564
rect 2691 -6616 2703 -6564
rect 2755 -6616 3092 -6564
rect 3144 -6616 3156 -6564
rect 3208 -6616 3220 -6564
rect 3272 -6616 7191 -6564
rect 7243 -6616 7255 -6564
rect 7307 -6616 7319 -6564
rect 7371 -6616 7708 -6564
rect 7760 -6616 7772 -6564
rect 7824 -6616 7836 -6564
rect 7888 -6576 11292 -6564
rect 7888 -6616 9331 -6576
rect 1132 -6632 9331 -6616
rect 9387 -6632 9411 -6576
rect 9467 -6632 9491 -6576
rect 9547 -6632 9633 -6576
rect 9689 -6632 9713 -6576
rect 9769 -6632 9793 -6576
rect 9849 -6616 11292 -6576
rect 11344 -6616 11356 -6564
rect 11408 -6616 11420 -6564
rect 11472 -6616 11809 -6564
rect 11861 -6616 11873 -6564
rect 11925 -6616 11937 -6564
rect 11989 -6616 15908 -6564
rect 15960 -6616 15972 -6564
rect 16024 -6616 16036 -6564
rect 16088 -6616 16425 -6564
rect 16477 -6616 16489 -6564
rect 16541 -6616 16553 -6564
rect 16605 -6576 18315 -6564
rect 16605 -6616 18048 -6576
rect 9849 -6632 18048 -6616
rect 18104 -6632 18128 -6576
rect 18184 -6632 18208 -6576
rect 18264 -6632 18315 -6576
rect 865 -6654 18315 -6632
rect 1601 -6709 17579 -6699
rect 1601 -6761 1608 -6709
rect 1660 -6761 1672 -6709
rect 1724 -6761 1736 -6709
rect 1788 -6761 2126 -6709
rect 2178 -6761 2190 -6709
rect 2242 -6761 2254 -6709
rect 2306 -6761 3803 -6709
rect 3855 -6761 3867 -6709
rect 3919 -6761 3931 -6709
rect 3983 -6761 4320 -6709
rect 4372 -6761 4384 -6709
rect 4436 -6761 4448 -6709
rect 4500 -6721 5963 -6709
rect 4500 -6761 4550 -6721
rect 1601 -6777 4550 -6761
rect 4606 -6777 4630 -6721
rect 4686 -6777 4710 -6721
rect 4766 -6777 5697 -6721
rect 5753 -6777 5777 -6721
rect 5833 -6777 5857 -6721
rect 5913 -6761 5963 -6721
rect 6015 -6761 6027 -6709
rect 6079 -6761 6091 -6709
rect 6143 -6761 6480 -6709
rect 6532 -6761 6544 -6709
rect 6596 -6761 6608 -6709
rect 6660 -6761 8157 -6709
rect 8209 -6761 8221 -6709
rect 8273 -6761 8285 -6709
rect 8337 -6761 8674 -6709
rect 8726 -6761 8738 -6709
rect 8790 -6761 8802 -6709
rect 8854 -6761 10326 -6709
rect 10378 -6761 10390 -6709
rect 10442 -6761 10454 -6709
rect 10506 -6761 10843 -6709
rect 10895 -6761 10907 -6709
rect 10959 -6761 10971 -6709
rect 11023 -6761 12520 -6709
rect 12572 -6761 12584 -6709
rect 12636 -6761 12648 -6709
rect 12700 -6761 13037 -6709
rect 13089 -6761 13101 -6709
rect 13153 -6761 13165 -6709
rect 13217 -6721 14680 -6709
rect 13217 -6761 13267 -6721
rect 5913 -6777 13267 -6761
rect 13323 -6777 13347 -6721
rect 13403 -6777 13427 -6721
rect 13483 -6777 14414 -6721
rect 14470 -6777 14494 -6721
rect 14550 -6777 14574 -6721
rect 14630 -6761 14680 -6721
rect 14732 -6761 14744 -6709
rect 14796 -6761 14808 -6709
rect 14860 -6761 15197 -6709
rect 15249 -6761 15261 -6709
rect 15313 -6761 15325 -6709
rect 15377 -6761 16874 -6709
rect 16926 -6761 16938 -6709
rect 16990 -6761 17002 -6709
rect 17054 -6761 17392 -6709
rect 17444 -6761 17456 -6709
rect 17508 -6761 17520 -6709
rect 17572 -6761 17579 -6709
rect 14630 -6777 17579 -6761
rect 1601 -6799 17579 -6777
rect 1298 -6870 17882 -6860
rect 1298 -6882 2833 -6870
rect 1298 -6938 1338 -6882
rect 1394 -6938 1418 -6882
rect 1474 -6938 1498 -6882
rect 1554 -6922 2833 -6882
rect 2885 -6922 2897 -6870
rect 2949 -6922 2961 -6870
rect 3013 -6922 3350 -6870
rect 3402 -6922 3414 -6870
rect 3466 -6922 3478 -6870
rect 3530 -6922 6933 -6870
rect 6985 -6922 6997 -6870
rect 7049 -6922 7061 -6870
rect 7113 -6922 7450 -6870
rect 7502 -6922 7514 -6870
rect 7566 -6922 7578 -6870
rect 7630 -6882 11550 -6870
rect 7630 -6922 8908 -6882
rect 1554 -6938 8908 -6922
rect 8964 -6938 8988 -6882
rect 9044 -6938 9068 -6882
rect 9124 -6938 10056 -6882
rect 10112 -6938 10136 -6882
rect 10192 -6938 10216 -6882
rect 10272 -6922 11550 -6882
rect 11602 -6922 11614 -6870
rect 11666 -6922 11678 -6870
rect 11730 -6922 12067 -6870
rect 12119 -6922 12131 -6870
rect 12183 -6922 12195 -6870
rect 12247 -6922 15650 -6870
rect 15702 -6922 15714 -6870
rect 15766 -6922 15778 -6870
rect 15830 -6922 16167 -6870
rect 16219 -6922 16231 -6870
rect 16283 -6922 16295 -6870
rect 16347 -6882 17882 -6870
rect 16347 -6922 17626 -6882
rect 10272 -6938 17626 -6922
rect 17682 -6938 17706 -6882
rect 17762 -6938 17786 -6882
rect 17842 -6938 17882 -6882
rect 1298 -6960 17882 -6938
rect 1343 -7010 17837 -7000
rect 1343 -7062 1350 -7010
rect 1402 -7062 1414 -7010
rect 1466 -7062 1478 -7010
rect 1530 -7062 1865 -7010
rect 1917 -7062 1929 -7010
rect 1981 -7062 1993 -7010
rect 2045 -7062 2383 -7010
rect 2435 -7062 2447 -7010
rect 2499 -7062 2511 -7010
rect 2563 -7062 3543 -7010
rect 3595 -7062 3607 -7010
rect 3659 -7062 3671 -7010
rect 3723 -7062 4060 -7010
rect 4112 -7062 4124 -7010
rect 4176 -7062 4188 -7010
rect 4240 -7062 4577 -7010
rect 4629 -7062 4641 -7010
rect 4693 -7062 4705 -7010
rect 4757 -7022 5706 -7010
rect 4757 -7062 4985 -7022
rect 1343 -7078 4985 -7062
rect 5041 -7078 5065 -7022
rect 5121 -7078 5145 -7022
rect 5201 -7078 5262 -7022
rect 5318 -7078 5342 -7022
rect 5398 -7078 5422 -7022
rect 5478 -7062 5706 -7022
rect 5758 -7062 5770 -7010
rect 5822 -7062 5834 -7010
rect 5886 -7062 6223 -7010
rect 6275 -7062 6287 -7010
rect 6339 -7062 6351 -7010
rect 6403 -7062 6740 -7010
rect 6792 -7062 6804 -7010
rect 6856 -7062 6868 -7010
rect 6920 -7062 7900 -7010
rect 7952 -7062 7964 -7010
rect 8016 -7062 8028 -7010
rect 8080 -7062 8417 -7010
rect 8469 -7062 8481 -7010
rect 8533 -7062 8545 -7010
rect 8597 -7062 8932 -7010
rect 8984 -7062 8996 -7010
rect 9048 -7062 9060 -7010
rect 9112 -7062 10068 -7010
rect 10120 -7062 10132 -7010
rect 10184 -7062 10196 -7010
rect 10248 -7062 10583 -7010
rect 10635 -7062 10647 -7010
rect 10699 -7062 10711 -7010
rect 10763 -7062 11100 -7010
rect 11152 -7062 11164 -7010
rect 11216 -7062 11228 -7010
rect 11280 -7062 12260 -7010
rect 12312 -7062 12324 -7010
rect 12376 -7062 12388 -7010
rect 12440 -7062 12777 -7010
rect 12829 -7062 12841 -7010
rect 12893 -7062 12905 -7010
rect 12957 -7062 13294 -7010
rect 13346 -7062 13358 -7010
rect 13410 -7062 13422 -7010
rect 13474 -7022 14423 -7010
rect 13474 -7062 13702 -7022
rect 5478 -7078 13702 -7062
rect 13758 -7078 13782 -7022
rect 13838 -7078 13862 -7022
rect 13918 -7078 13979 -7022
rect 14035 -7078 14059 -7022
rect 14115 -7078 14139 -7022
rect 14195 -7062 14423 -7022
rect 14475 -7062 14487 -7010
rect 14539 -7062 14551 -7010
rect 14603 -7062 14940 -7010
rect 14992 -7062 15004 -7010
rect 15056 -7062 15068 -7010
rect 15120 -7062 15457 -7010
rect 15509 -7062 15521 -7010
rect 15573 -7062 15585 -7010
rect 15637 -7062 16617 -7010
rect 16669 -7062 16681 -7010
rect 16733 -7062 16745 -7010
rect 16797 -7062 17135 -7010
rect 17187 -7062 17199 -7010
rect 17251 -7062 17263 -7010
rect 17315 -7062 17650 -7010
rect 17702 -7062 17714 -7010
rect 17766 -7062 17778 -7010
rect 17830 -7062 17837 -7010
rect 14195 -7078 17837 -7062
rect 1343 -7100 17837 -7078
rect 1473 -7459 17707 -7438
rect 1473 -7511 1523 -7459
rect 1575 -7511 1587 -7459
rect 1639 -7511 1651 -7459
rect 1703 -7511 1719 -7459
rect 1771 -7511 1783 -7459
rect 1835 -7511 1847 -7459
rect 1899 -7511 2009 -7459
rect 2061 -7511 2073 -7459
rect 2125 -7511 2137 -7459
rect 2189 -7511 2205 -7459
rect 2257 -7511 2269 -7459
rect 2321 -7511 2333 -7459
rect 2385 -7460 3721 -7459
rect 2385 -7511 3433 -7460
rect 1473 -7516 3433 -7511
rect 3489 -7516 3513 -7460
rect 3569 -7516 3593 -7460
rect 3649 -7511 3721 -7460
rect 3773 -7511 3785 -7459
rect 3837 -7511 3849 -7459
rect 3901 -7511 3917 -7459
rect 3969 -7511 3981 -7459
rect 4033 -7511 4045 -7459
rect 4097 -7511 4207 -7459
rect 4259 -7511 4271 -7459
rect 4323 -7511 4335 -7459
rect 4387 -7511 4403 -7459
rect 4455 -7511 4467 -7459
rect 4519 -7511 4531 -7459
rect 4583 -7511 5880 -7459
rect 5932 -7511 5944 -7459
rect 5996 -7511 6008 -7459
rect 6060 -7511 6076 -7459
rect 6128 -7511 6140 -7459
rect 6192 -7511 6204 -7459
rect 6256 -7511 6366 -7459
rect 6418 -7511 6430 -7459
rect 6482 -7511 6494 -7459
rect 6546 -7511 6562 -7459
rect 6614 -7511 6626 -7459
rect 6678 -7511 6690 -7459
rect 6742 -7460 8078 -7459
rect 6742 -7511 6814 -7460
rect 3649 -7516 6814 -7511
rect 6870 -7516 6894 -7460
rect 6950 -7516 6974 -7460
rect 7030 -7511 8078 -7460
rect 8130 -7511 8142 -7459
rect 8194 -7511 8206 -7459
rect 8258 -7511 8274 -7459
rect 8326 -7511 8338 -7459
rect 8390 -7511 8402 -7459
rect 8454 -7511 8564 -7459
rect 8616 -7511 8628 -7459
rect 8680 -7511 8692 -7459
rect 8744 -7511 8760 -7459
rect 8812 -7511 8824 -7459
rect 8876 -7511 8888 -7459
rect 8940 -7511 10240 -7459
rect 10292 -7511 10304 -7459
rect 10356 -7511 10368 -7459
rect 10420 -7511 10436 -7459
rect 10488 -7511 10500 -7459
rect 10552 -7511 10564 -7459
rect 10616 -7511 10726 -7459
rect 10778 -7511 10790 -7459
rect 10842 -7511 10854 -7459
rect 10906 -7511 10922 -7459
rect 10974 -7511 10986 -7459
rect 11038 -7511 11050 -7459
rect 11102 -7460 12438 -7459
rect 11102 -7511 12150 -7460
rect 7030 -7516 12150 -7511
rect 12206 -7516 12230 -7460
rect 12286 -7516 12310 -7460
rect 12366 -7511 12438 -7460
rect 12490 -7511 12502 -7459
rect 12554 -7511 12566 -7459
rect 12618 -7511 12634 -7459
rect 12686 -7511 12698 -7459
rect 12750 -7511 12762 -7459
rect 12814 -7511 12924 -7459
rect 12976 -7511 12988 -7459
rect 13040 -7511 13052 -7459
rect 13104 -7511 13120 -7459
rect 13172 -7511 13184 -7459
rect 13236 -7511 13248 -7459
rect 13300 -7511 14597 -7459
rect 14649 -7511 14661 -7459
rect 14713 -7511 14725 -7459
rect 14777 -7511 14793 -7459
rect 14845 -7511 14857 -7459
rect 14909 -7511 14921 -7459
rect 14973 -7511 15083 -7459
rect 15135 -7511 15147 -7459
rect 15199 -7511 15211 -7459
rect 15263 -7511 15279 -7459
rect 15331 -7511 15343 -7459
rect 15395 -7511 15407 -7459
rect 15459 -7460 16795 -7459
rect 15459 -7511 15531 -7460
rect 12366 -7516 15531 -7511
rect 15587 -7516 15611 -7460
rect 15667 -7516 15691 -7460
rect 15747 -7511 16795 -7460
rect 16847 -7511 16859 -7459
rect 16911 -7511 16923 -7459
rect 16975 -7511 16991 -7459
rect 17043 -7511 17055 -7459
rect 17107 -7511 17119 -7459
rect 17171 -7511 17281 -7459
rect 17333 -7511 17345 -7459
rect 17397 -7511 17409 -7459
rect 17461 -7511 17477 -7459
rect 17529 -7511 17541 -7459
rect 17593 -7511 17605 -7459
rect 17657 -7511 17707 -7459
rect 15747 -7516 17707 -7511
rect 1473 -7526 17707 -7516
rect 3393 -7538 3693 -7526
rect 6770 -7538 7070 -7526
rect 12110 -7538 12410 -7526
rect 15487 -7538 15787 -7526
rect 1473 -7637 17707 -7620
rect 1473 -7689 1523 -7637
rect 1575 -7689 1587 -7637
rect 1639 -7689 1651 -7637
rect 1703 -7689 1719 -7637
rect 1771 -7689 1783 -7637
rect 1835 -7689 1847 -7637
rect 1899 -7689 2009 -7637
rect 2061 -7689 2073 -7637
rect 2125 -7689 2137 -7637
rect 2189 -7689 2205 -7637
rect 2257 -7689 2269 -7637
rect 2321 -7689 2333 -7637
rect 2385 -7689 2733 -7637
rect 2785 -7689 2797 -7637
rect 2849 -7689 2861 -7637
rect 2913 -7689 2929 -7637
rect 2981 -7689 2993 -7637
rect 3045 -7689 3057 -7637
rect 3109 -7689 3121 -7637
rect 3173 -7689 3189 -7637
rect 3241 -7689 3253 -7637
rect 3305 -7689 3317 -7637
rect 3369 -7689 3721 -7637
rect 3773 -7689 3785 -7637
rect 3837 -7689 3849 -7637
rect 3901 -7689 3917 -7637
rect 3969 -7689 3981 -7637
rect 4033 -7689 4045 -7637
rect 4097 -7689 4207 -7637
rect 4259 -7689 4271 -7637
rect 4323 -7689 4335 -7637
rect 4387 -7689 4403 -7637
rect 4455 -7689 4467 -7637
rect 4519 -7689 4531 -7637
rect 4583 -7689 5880 -7637
rect 5932 -7689 5944 -7637
rect 5996 -7689 6008 -7637
rect 6060 -7689 6076 -7637
rect 6128 -7689 6140 -7637
rect 6192 -7689 6204 -7637
rect 6256 -7689 6366 -7637
rect 6418 -7689 6430 -7637
rect 6482 -7689 6494 -7637
rect 6546 -7689 6562 -7637
rect 6614 -7689 6626 -7637
rect 6678 -7689 6690 -7637
rect 6742 -7689 7094 -7637
rect 7146 -7689 7158 -7637
rect 7210 -7689 7222 -7637
rect 7274 -7689 7290 -7637
rect 7342 -7689 7354 -7637
rect 7406 -7689 7418 -7637
rect 7470 -7689 7482 -7637
rect 7534 -7689 7550 -7637
rect 7602 -7689 7614 -7637
rect 7666 -7689 7678 -7637
rect 7730 -7689 8078 -7637
rect 8130 -7689 8142 -7637
rect 8194 -7689 8206 -7637
rect 8258 -7689 8274 -7637
rect 8326 -7689 8338 -7637
rect 8390 -7689 8402 -7637
rect 8454 -7689 8564 -7637
rect 8616 -7689 8628 -7637
rect 8680 -7689 8692 -7637
rect 8744 -7689 8760 -7637
rect 8812 -7689 8824 -7637
rect 8876 -7689 8888 -7637
rect 8940 -7689 10240 -7637
rect 10292 -7689 10304 -7637
rect 10356 -7689 10368 -7637
rect 10420 -7689 10436 -7637
rect 10488 -7689 10500 -7637
rect 10552 -7689 10564 -7637
rect 10616 -7689 10726 -7637
rect 10778 -7689 10790 -7637
rect 10842 -7689 10854 -7637
rect 10906 -7689 10922 -7637
rect 10974 -7689 10986 -7637
rect 11038 -7689 11050 -7637
rect 11102 -7689 11450 -7637
rect 11502 -7689 11514 -7637
rect 11566 -7689 11578 -7637
rect 11630 -7689 11646 -7637
rect 11698 -7689 11710 -7637
rect 11762 -7689 11774 -7637
rect 11826 -7689 11838 -7637
rect 11890 -7689 11906 -7637
rect 11958 -7689 11970 -7637
rect 12022 -7689 12034 -7637
rect 12086 -7689 12438 -7637
rect 12490 -7689 12502 -7637
rect 12554 -7689 12566 -7637
rect 12618 -7689 12634 -7637
rect 12686 -7689 12698 -7637
rect 12750 -7689 12762 -7637
rect 12814 -7689 12924 -7637
rect 12976 -7689 12988 -7637
rect 13040 -7689 13052 -7637
rect 13104 -7689 13120 -7637
rect 13172 -7689 13184 -7637
rect 13236 -7689 13248 -7637
rect 13300 -7689 14597 -7637
rect 14649 -7689 14661 -7637
rect 14713 -7689 14725 -7637
rect 14777 -7689 14793 -7637
rect 14845 -7689 14857 -7637
rect 14909 -7689 14921 -7637
rect 14973 -7689 15083 -7637
rect 15135 -7689 15147 -7637
rect 15199 -7689 15211 -7637
rect 15263 -7689 15279 -7637
rect 15331 -7689 15343 -7637
rect 15395 -7689 15407 -7637
rect 15459 -7689 15811 -7637
rect 15863 -7689 15875 -7637
rect 15927 -7689 15939 -7637
rect 15991 -7689 16007 -7637
rect 16059 -7689 16071 -7637
rect 16123 -7689 16135 -7637
rect 16187 -7689 16199 -7637
rect 16251 -7689 16267 -7637
rect 16319 -7689 16331 -7637
rect 16383 -7689 16395 -7637
rect 16447 -7689 16795 -7637
rect 16847 -7689 16859 -7637
rect 16911 -7689 16923 -7637
rect 16975 -7689 16991 -7637
rect 17043 -7689 17055 -7637
rect 17107 -7689 17119 -7637
rect 17171 -7689 17281 -7637
rect 17333 -7689 17345 -7637
rect 17397 -7689 17409 -7637
rect 17461 -7689 17477 -7637
rect 17529 -7689 17541 -7637
rect 17593 -7689 17605 -7637
rect 17657 -7689 17707 -7637
rect 1473 -7708 17707 -7689
rect 1473 -7776 17707 -7758
rect 1473 -7828 1523 -7776
rect 1575 -7828 1587 -7776
rect 1639 -7828 1651 -7776
rect 1703 -7828 1719 -7776
rect 1771 -7828 1783 -7776
rect 1835 -7828 1847 -7776
rect 1899 -7828 2009 -7776
rect 2061 -7828 2073 -7776
rect 2125 -7828 2137 -7776
rect 2189 -7828 2205 -7776
rect 2257 -7828 2269 -7776
rect 2321 -7828 2333 -7776
rect 2385 -7780 3721 -7776
rect 2385 -7828 2465 -7780
rect 1473 -7836 2465 -7828
rect 2521 -7836 2545 -7780
rect 2601 -7836 2625 -7780
rect 2681 -7828 3721 -7780
rect 3773 -7828 3785 -7776
rect 3837 -7828 3849 -7776
rect 3901 -7828 3917 -7776
rect 3969 -7828 3981 -7776
rect 4033 -7828 4045 -7776
rect 4097 -7828 4207 -7776
rect 4259 -7828 4271 -7776
rect 4323 -7828 4335 -7776
rect 4387 -7828 4403 -7776
rect 4455 -7828 4467 -7776
rect 4519 -7828 4531 -7776
rect 4583 -7828 5880 -7776
rect 5932 -7828 5944 -7776
rect 5996 -7828 6008 -7776
rect 6060 -7828 6076 -7776
rect 6128 -7828 6140 -7776
rect 6192 -7828 6204 -7776
rect 6256 -7828 6366 -7776
rect 6418 -7828 6430 -7776
rect 6482 -7828 6494 -7776
rect 6546 -7828 6562 -7776
rect 6614 -7828 6626 -7776
rect 6678 -7828 6690 -7776
rect 6742 -7780 8078 -7776
rect 6742 -7828 7782 -7780
rect 2681 -7836 7782 -7828
rect 7838 -7836 7862 -7780
rect 7918 -7836 7942 -7780
rect 7998 -7828 8078 -7780
rect 8130 -7828 8142 -7776
rect 8194 -7828 8206 -7776
rect 8258 -7828 8274 -7776
rect 8326 -7828 8338 -7776
rect 8390 -7828 8402 -7776
rect 8454 -7828 8564 -7776
rect 8616 -7828 8628 -7776
rect 8680 -7828 8692 -7776
rect 8744 -7828 8760 -7776
rect 8812 -7828 8824 -7776
rect 8876 -7828 8888 -7776
rect 8940 -7828 10240 -7776
rect 10292 -7828 10304 -7776
rect 10356 -7828 10368 -7776
rect 10420 -7828 10436 -7776
rect 10488 -7828 10500 -7776
rect 10552 -7828 10564 -7776
rect 10616 -7828 10726 -7776
rect 10778 -7828 10790 -7776
rect 10842 -7828 10854 -7776
rect 10906 -7828 10922 -7776
rect 10974 -7828 10986 -7776
rect 11038 -7828 11050 -7776
rect 11102 -7780 12438 -7776
rect 11102 -7828 11182 -7780
rect 7998 -7836 11182 -7828
rect 11238 -7836 11262 -7780
rect 11318 -7836 11342 -7780
rect 11398 -7828 12438 -7780
rect 12490 -7828 12502 -7776
rect 12554 -7828 12566 -7776
rect 12618 -7828 12634 -7776
rect 12686 -7828 12698 -7776
rect 12750 -7828 12762 -7776
rect 12814 -7828 12924 -7776
rect 12976 -7828 12988 -7776
rect 13040 -7828 13052 -7776
rect 13104 -7828 13120 -7776
rect 13172 -7828 13184 -7776
rect 13236 -7828 13248 -7776
rect 13300 -7828 14597 -7776
rect 14649 -7828 14661 -7776
rect 14713 -7828 14725 -7776
rect 14777 -7828 14793 -7776
rect 14845 -7828 14857 -7776
rect 14909 -7828 14921 -7776
rect 14973 -7828 15083 -7776
rect 15135 -7828 15147 -7776
rect 15199 -7828 15211 -7776
rect 15263 -7828 15279 -7776
rect 15331 -7828 15343 -7776
rect 15395 -7828 15407 -7776
rect 15459 -7780 16795 -7776
rect 15459 -7828 16499 -7780
rect 11398 -7836 16499 -7828
rect 16555 -7836 16579 -7780
rect 16635 -7836 16659 -7780
rect 16715 -7828 16795 -7780
rect 16847 -7828 16859 -7776
rect 16911 -7828 16923 -7776
rect 16975 -7828 16991 -7776
rect 17043 -7828 17055 -7776
rect 17107 -7828 17119 -7776
rect 17171 -7828 17281 -7776
rect 17333 -7828 17345 -7776
rect 17397 -7828 17409 -7776
rect 17461 -7828 17477 -7776
rect 17529 -7828 17541 -7776
rect 17593 -7828 17605 -7776
rect 17657 -7828 17707 -7776
rect 16715 -7836 17707 -7828
rect 1473 -7846 17707 -7836
rect 2425 -7858 2725 -7846
rect 7738 -7858 8038 -7846
rect 11142 -7858 11442 -7846
rect 16455 -7858 16755 -7846
rect 1298 -8199 17882 -8189
rect 1298 -8211 1607 -8199
rect 1298 -8267 1338 -8211
rect 1394 -8267 1418 -8211
rect 1474 -8267 1498 -8211
rect 1554 -8251 1607 -8211
rect 1659 -8251 1671 -8199
rect 1723 -8251 1735 -8199
rect 1787 -8251 2125 -8199
rect 2177 -8251 2189 -8199
rect 2241 -8251 2253 -8199
rect 2305 -8251 3802 -8199
rect 3854 -8251 3866 -8199
rect 3918 -8251 3930 -8199
rect 3982 -8251 4319 -8199
rect 4371 -8251 4383 -8199
rect 4435 -8251 4447 -8199
rect 4499 -8251 5964 -8199
rect 6016 -8251 6028 -8199
rect 6080 -8251 6092 -8199
rect 6144 -8251 6481 -8199
rect 6533 -8251 6545 -8199
rect 6597 -8251 6609 -8199
rect 6661 -8251 8158 -8199
rect 8210 -8251 8222 -8199
rect 8274 -8251 8286 -8199
rect 8338 -8251 8675 -8199
rect 8727 -8251 8739 -8199
rect 8791 -8251 8803 -8199
rect 8855 -8211 10325 -8199
rect 8855 -8251 8908 -8211
rect 1554 -8267 8908 -8251
rect 8964 -8267 8988 -8211
rect 9044 -8267 9068 -8211
rect 9124 -8267 10056 -8211
rect 10112 -8267 10136 -8211
rect 10192 -8267 10216 -8211
rect 10272 -8251 10325 -8211
rect 10377 -8251 10389 -8199
rect 10441 -8251 10453 -8199
rect 10505 -8251 10842 -8199
rect 10894 -8251 10906 -8199
rect 10958 -8251 10970 -8199
rect 11022 -8251 12519 -8199
rect 12571 -8251 12583 -8199
rect 12635 -8251 12647 -8199
rect 12699 -8251 13036 -8199
rect 13088 -8251 13100 -8199
rect 13152 -8251 13164 -8199
rect 13216 -8251 14681 -8199
rect 14733 -8251 14745 -8199
rect 14797 -8251 14809 -8199
rect 14861 -8251 15198 -8199
rect 15250 -8251 15262 -8199
rect 15314 -8251 15326 -8199
rect 15378 -8251 16875 -8199
rect 16927 -8251 16939 -8199
rect 16991 -8251 17003 -8199
rect 17055 -8251 17393 -8199
rect 17445 -8251 17457 -8199
rect 17509 -8251 17521 -8199
rect 17573 -8211 17882 -8199
rect 17573 -8251 17626 -8211
rect 10272 -8267 17626 -8251
rect 17682 -8267 17706 -8211
rect 17762 -8267 17786 -8211
rect 17842 -8267 17882 -8211
rect 1298 -8289 17882 -8267
rect 2570 -8368 16610 -8358
rect 2570 -8420 2577 -8368
rect 2629 -8420 2641 -8368
rect 2693 -8420 2705 -8368
rect 2757 -8420 3094 -8368
rect 3146 -8420 3158 -8368
rect 3210 -8420 3222 -8368
rect 3274 -8380 7189 -8368
rect 3274 -8420 4550 -8380
rect 2570 -8436 4550 -8420
rect 4606 -8436 4630 -8380
rect 4686 -8436 4710 -8380
rect 4766 -8436 5697 -8380
rect 5753 -8436 5777 -8380
rect 5833 -8436 5857 -8380
rect 5913 -8420 7189 -8380
rect 7241 -8420 7253 -8368
rect 7305 -8420 7317 -8368
rect 7369 -8420 7706 -8368
rect 7758 -8420 7770 -8368
rect 7822 -8420 7834 -8368
rect 7886 -8420 11294 -8368
rect 11346 -8420 11358 -8368
rect 11410 -8420 11422 -8368
rect 11474 -8420 11811 -8368
rect 11863 -8420 11875 -8368
rect 11927 -8420 11939 -8368
rect 11991 -8380 15906 -8368
rect 11991 -8420 13267 -8380
rect 5913 -8436 13267 -8420
rect 13323 -8436 13347 -8380
rect 13403 -8436 13427 -8380
rect 13483 -8436 14414 -8380
rect 14470 -8436 14494 -8380
rect 14550 -8436 14574 -8380
rect 14630 -8420 15906 -8380
rect 15958 -8420 15970 -8368
rect 16022 -8420 16034 -8368
rect 16086 -8420 16423 -8368
rect 16475 -8420 16487 -8368
rect 16539 -8420 16551 -8368
rect 16603 -8420 16610 -8368
rect 14630 -8436 16610 -8420
rect 2570 -8458 16610 -8436
rect 876 -8531 18304 -8521
rect 876 -8543 1348 -8531
rect 876 -8599 916 -8543
rect 972 -8599 996 -8543
rect 1052 -8599 1076 -8543
rect 1132 -8583 1348 -8543
rect 1400 -8583 1412 -8531
rect 1464 -8583 1476 -8531
rect 1528 -8583 1865 -8531
rect 1917 -8583 1929 -8531
rect 1981 -8583 1993 -8531
rect 2045 -8583 2382 -8531
rect 2434 -8583 2446 -8531
rect 2498 -8583 2510 -8531
rect 2562 -8583 3543 -8531
rect 3595 -8583 3607 -8531
rect 3659 -8583 3671 -8531
rect 3723 -8583 4060 -8531
rect 4112 -8583 4124 -8531
rect 4176 -8583 4188 -8531
rect 4240 -8583 4575 -8531
rect 4627 -8583 4639 -8531
rect 4691 -8583 4703 -8531
rect 4755 -8583 5708 -8531
rect 5760 -8583 5772 -8531
rect 5824 -8583 5836 -8531
rect 5888 -8583 6223 -8531
rect 6275 -8583 6287 -8531
rect 6339 -8583 6351 -8531
rect 6403 -8583 6740 -8531
rect 6792 -8583 6804 -8531
rect 6856 -8583 6868 -8531
rect 6920 -8583 7901 -8531
rect 7953 -8583 7965 -8531
rect 8017 -8583 8029 -8531
rect 8081 -8583 8417 -8531
rect 8469 -8583 8481 -8531
rect 8533 -8583 8545 -8531
rect 8597 -8583 8935 -8531
rect 8987 -8583 8999 -8531
rect 9051 -8583 9063 -8531
rect 9115 -8543 10065 -8531
rect 9115 -8583 9331 -8543
rect 1132 -8599 9331 -8583
rect 9387 -8599 9411 -8543
rect 9467 -8599 9491 -8543
rect 9547 -8599 9633 -8543
rect 9689 -8599 9713 -8543
rect 9769 -8599 9793 -8543
rect 9849 -8583 10065 -8543
rect 10117 -8583 10129 -8531
rect 10181 -8583 10193 -8531
rect 10245 -8583 10583 -8531
rect 10635 -8583 10647 -8531
rect 10699 -8583 10711 -8531
rect 10763 -8583 11099 -8531
rect 11151 -8583 11163 -8531
rect 11215 -8583 11227 -8531
rect 11279 -8583 12260 -8531
rect 12312 -8583 12324 -8531
rect 12376 -8583 12388 -8531
rect 12440 -8583 12777 -8531
rect 12829 -8583 12841 -8531
rect 12893 -8583 12905 -8531
rect 12957 -8583 13292 -8531
rect 13344 -8583 13356 -8531
rect 13408 -8583 13420 -8531
rect 13472 -8583 14425 -8531
rect 14477 -8583 14489 -8531
rect 14541 -8583 14553 -8531
rect 14605 -8583 14940 -8531
rect 14992 -8583 15004 -8531
rect 15056 -8583 15068 -8531
rect 15120 -8583 15457 -8531
rect 15509 -8583 15521 -8531
rect 15573 -8583 15585 -8531
rect 15637 -8583 16618 -8531
rect 16670 -8583 16682 -8531
rect 16734 -8583 16746 -8531
rect 16798 -8583 17135 -8531
rect 17187 -8583 17199 -8531
rect 17251 -8583 17263 -8531
rect 17315 -8583 17652 -8531
rect 17704 -8583 17716 -8531
rect 17768 -8583 17780 -8531
rect 17832 -8543 18304 -8531
rect 17832 -8583 18048 -8543
rect 9849 -8599 18048 -8583
rect 18104 -8599 18128 -8543
rect 18184 -8599 18208 -8543
rect 18264 -8599 18304 -8543
rect 876 -8621 18304 -8599
rect 2827 -8699 16353 -8689
rect 2827 -8751 2834 -8699
rect 2886 -8751 2898 -8699
rect 2950 -8751 2962 -8699
rect 3014 -8751 3351 -8699
rect 3403 -8751 3415 -8699
rect 3467 -8751 3479 -8699
rect 3531 -8711 6931 -8699
rect 3531 -8751 4985 -8711
rect 2827 -8767 4985 -8751
rect 5041 -8767 5065 -8711
rect 5121 -8767 5145 -8711
rect 5201 -8767 5262 -8711
rect 5318 -8767 5342 -8711
rect 5398 -8767 5422 -8711
rect 5478 -8751 6931 -8711
rect 6983 -8751 6995 -8699
rect 7047 -8751 7059 -8699
rect 7111 -8751 7449 -8699
rect 7501 -8751 7513 -8699
rect 7565 -8751 7577 -8699
rect 7629 -8751 11551 -8699
rect 11603 -8751 11615 -8699
rect 11667 -8751 11679 -8699
rect 11731 -8751 12069 -8699
rect 12121 -8751 12133 -8699
rect 12185 -8751 12197 -8699
rect 12249 -8711 15649 -8699
rect 12249 -8751 13702 -8711
rect 5478 -8767 13702 -8751
rect 13758 -8767 13782 -8711
rect 13838 -8767 13862 -8711
rect 13918 -8767 13979 -8711
rect 14035 -8767 14059 -8711
rect 14115 -8767 14139 -8711
rect 14195 -8751 15649 -8711
rect 15701 -8751 15713 -8699
rect 15765 -8751 15777 -8699
rect 15829 -8751 16166 -8699
rect 16218 -8751 16230 -8699
rect 16282 -8751 16294 -8699
rect 16346 -8751 16353 -8699
rect 14195 -8767 16353 -8751
rect 2827 -8789 16353 -8767
<< via2 >>
rect 4985 -52 5041 4
rect 5065 -52 5121 4
rect 5145 -52 5201 4
rect 5262 -52 5318 4
rect 5342 -52 5398 4
rect 5422 -52 5478 4
rect 13702 -52 13758 4
rect 13782 -52 13838 4
rect 13862 -52 13918 4
rect 13979 -52 14035 4
rect 14059 -52 14115 4
rect 14139 -52 14195 4
rect 916 -221 972 -165
rect 996 -221 1052 -165
rect 1076 -221 1132 -165
rect 9331 -221 9387 -165
rect 9411 -221 9467 -165
rect 9491 -221 9547 -165
rect 9633 -221 9689 -165
rect 9713 -221 9769 -165
rect 9793 -221 9849 -165
rect 18048 -221 18104 -165
rect 18128 -221 18184 -165
rect 18208 -221 18264 -165
rect 4550 -384 4606 -328
rect 4630 -384 4686 -328
rect 4710 -384 4766 -328
rect 5697 -384 5753 -328
rect 5777 -384 5833 -328
rect 5857 -384 5913 -328
rect 13267 -384 13323 -328
rect 13347 -384 13403 -328
rect 13427 -384 13483 -328
rect 14414 -384 14470 -328
rect 14494 -384 14550 -328
rect 14574 -384 14630 -328
rect 1338 -552 1394 -496
rect 1418 -552 1474 -496
rect 1498 -552 1554 -496
rect 8908 -552 8964 -496
rect 8988 -552 9044 -496
rect 9068 -552 9124 -496
rect 10056 -552 10112 -496
rect 10136 -552 10192 -496
rect 10216 -552 10272 -496
rect 17626 -552 17682 -496
rect 17706 -552 17762 -496
rect 17786 -552 17842 -496
rect 2465 -984 2521 -928
rect 2545 -984 2601 -928
rect 2625 -984 2681 -928
rect 7782 -984 7838 -928
rect 7862 -984 7918 -928
rect 7942 -984 7998 -928
rect 11182 -984 11238 -928
rect 11262 -984 11318 -928
rect 11342 -984 11398 -928
rect 16499 -984 16555 -928
rect 16579 -984 16635 -928
rect 16659 -984 16715 -928
rect 3433 -1304 3489 -1248
rect 3513 -1304 3569 -1248
rect 3593 -1304 3649 -1248
rect 6814 -1304 6870 -1248
rect 6894 -1304 6950 -1248
rect 6974 -1304 7030 -1248
rect 12150 -1304 12206 -1248
rect 12230 -1304 12286 -1248
rect 12310 -1304 12366 -1248
rect 15531 -1304 15587 -1248
rect 15611 -1304 15667 -1248
rect 15691 -1304 15747 -1248
rect 4985 -1742 5041 -1686
rect 5065 -1742 5121 -1686
rect 5145 -1742 5201 -1686
rect 5262 -1742 5318 -1686
rect 5342 -1742 5398 -1686
rect 5422 -1742 5478 -1686
rect 13702 -1742 13758 -1686
rect 13782 -1742 13838 -1686
rect 13862 -1742 13918 -1686
rect 13979 -1742 14035 -1686
rect 14059 -1742 14115 -1686
rect 14139 -1742 14195 -1686
rect 1338 -1882 1394 -1826
rect 1418 -1882 1474 -1826
rect 1498 -1882 1554 -1826
rect 8908 -1882 8964 -1826
rect 8988 -1882 9044 -1826
rect 9068 -1882 9124 -1826
rect 10056 -1882 10112 -1826
rect 10136 -1882 10192 -1826
rect 10216 -1882 10272 -1826
rect 17626 -1882 17682 -1826
rect 17706 -1882 17762 -1826
rect 17786 -1882 17842 -1826
rect 4550 -2043 4606 -1987
rect 4630 -2043 4686 -1987
rect 4710 -2043 4766 -1987
rect 5697 -2043 5753 -1987
rect 5777 -2043 5833 -1987
rect 5857 -2043 5913 -1987
rect 13267 -2043 13323 -1987
rect 13347 -2043 13403 -1987
rect 13427 -2043 13483 -1987
rect 14414 -2043 14470 -1987
rect 14494 -2043 14550 -1987
rect 14574 -2043 14630 -1987
rect 916 -2187 972 -2131
rect 996 -2187 1052 -2131
rect 1076 -2187 1132 -2131
rect 9331 -2187 9387 -2131
rect 9411 -2187 9467 -2131
rect 9491 -2187 9547 -2131
rect 9633 -2187 9689 -2131
rect 9713 -2187 9769 -2131
rect 9793 -2187 9849 -2131
rect 18048 -2187 18104 -2131
rect 18128 -2187 18184 -2131
rect 18208 -2187 18264 -2131
rect 3433 -2631 3489 -2575
rect 3513 -2631 3569 -2575
rect 3593 -2631 3649 -2575
rect 6814 -2642 6870 -2586
rect 6894 -2642 6950 -2586
rect 6974 -2642 7030 -2586
rect 12150 -2642 12206 -2586
rect 12230 -2642 12286 -2586
rect 12310 -2642 12366 -2586
rect 15531 -2631 15587 -2575
rect 15611 -2631 15667 -2575
rect 15691 -2631 15747 -2575
rect 2465 -2963 2521 -2907
rect 2545 -2963 2601 -2907
rect 2625 -2963 2681 -2907
rect 7782 -2963 7838 -2907
rect 7862 -2963 7918 -2907
rect 7942 -2963 7998 -2907
rect 11182 -2963 11238 -2907
rect 11262 -2963 11318 -2907
rect 11342 -2963 11398 -2907
rect 16499 -2963 16555 -2907
rect 16579 -2963 16635 -2907
rect 16659 -2963 16715 -2907
rect 1338 -3394 1394 -3338
rect 1418 -3394 1474 -3338
rect 1498 -3394 1554 -3338
rect 8908 -3394 8964 -3338
rect 8988 -3394 9044 -3338
rect 9068 -3394 9124 -3338
rect 10056 -3394 10112 -3338
rect 10136 -3394 10192 -3338
rect 10216 -3394 10272 -3338
rect 17626 -3394 17682 -3338
rect 17706 -3394 17762 -3338
rect 17786 -3394 17842 -3338
rect 4550 -3563 4606 -3507
rect 4630 -3563 4686 -3507
rect 4710 -3563 4766 -3507
rect 5697 -3563 5753 -3507
rect 5777 -3563 5833 -3507
rect 5857 -3563 5913 -3507
rect 13267 -3563 13323 -3507
rect 13347 -3563 13403 -3507
rect 13427 -3563 13483 -3507
rect 14414 -3563 14470 -3507
rect 14494 -3563 14550 -3507
rect 14574 -3563 14630 -3507
rect 916 -3725 972 -3669
rect 996 -3725 1052 -3669
rect 1076 -3725 1132 -3669
rect 9331 -3725 9387 -3669
rect 9411 -3725 9467 -3669
rect 9491 -3725 9547 -3669
rect 9633 -3725 9689 -3669
rect 9713 -3725 9769 -3669
rect 9793 -3725 9849 -3669
rect 18048 -3725 18104 -3669
rect 18128 -3725 18184 -3669
rect 18208 -3725 18264 -3669
rect 4985 -3894 5041 -3838
rect 5065 -3894 5121 -3838
rect 5145 -3894 5201 -3838
rect 5262 -3894 5318 -3838
rect 5342 -3894 5398 -3838
rect 5422 -3894 5478 -3838
rect 13702 -3894 13758 -3838
rect 13782 -3894 13838 -3838
rect 13862 -3894 13918 -3838
rect 13979 -3894 14035 -3838
rect 14059 -3894 14115 -3838
rect 14139 -3894 14195 -3838
rect 4985 -4925 5041 -4869
rect 5065 -4925 5121 -4869
rect 5145 -4925 5201 -4869
rect 5262 -4925 5318 -4869
rect 5342 -4925 5398 -4869
rect 5422 -4925 5478 -4869
rect 13702 -4925 13758 -4869
rect 13782 -4925 13838 -4869
rect 13862 -4925 13918 -4869
rect 13979 -4925 14035 -4869
rect 14059 -4925 14115 -4869
rect 14139 -4925 14195 -4869
rect 916 -5094 972 -5038
rect 996 -5094 1052 -5038
rect 1076 -5094 1132 -5038
rect 9331 -5094 9387 -5038
rect 9411 -5094 9467 -5038
rect 9491 -5094 9547 -5038
rect 9633 -5094 9689 -5038
rect 9713 -5094 9769 -5038
rect 9793 -5094 9849 -5038
rect 18048 -5094 18104 -5038
rect 18128 -5094 18184 -5038
rect 18208 -5094 18264 -5038
rect 4550 -5257 4606 -5201
rect 4630 -5257 4686 -5201
rect 4710 -5257 4766 -5201
rect 5697 -5257 5753 -5201
rect 5777 -5257 5833 -5201
rect 5857 -5257 5913 -5201
rect 13267 -5257 13323 -5201
rect 13347 -5257 13403 -5201
rect 13427 -5257 13483 -5201
rect 14414 -5257 14470 -5201
rect 14494 -5257 14550 -5201
rect 14574 -5257 14630 -5201
rect 1338 -5426 1394 -5370
rect 1418 -5426 1474 -5370
rect 1498 -5426 1554 -5370
rect 8908 -5426 8964 -5370
rect 8988 -5426 9044 -5370
rect 9068 -5426 9124 -5370
rect 10056 -5426 10112 -5370
rect 10136 -5426 10192 -5370
rect 10216 -5426 10272 -5370
rect 17626 -5426 17682 -5370
rect 17706 -5426 17762 -5370
rect 17786 -5426 17842 -5370
rect 2465 -5857 2521 -5801
rect 2545 -5857 2601 -5801
rect 2625 -5857 2681 -5801
rect 7782 -5857 7838 -5801
rect 7862 -5857 7918 -5801
rect 7942 -5857 7998 -5801
rect 11182 -5857 11238 -5801
rect 11262 -5857 11318 -5801
rect 11342 -5857 11398 -5801
rect 16499 -5857 16555 -5801
rect 16579 -5857 16635 -5801
rect 16659 -5857 16715 -5801
rect 3433 -6189 3489 -6133
rect 3513 -6189 3569 -6133
rect 3593 -6189 3649 -6133
rect 6814 -6189 6870 -6133
rect 6894 -6189 6950 -6133
rect 6974 -6189 7030 -6133
rect 12150 -6189 12206 -6133
rect 12230 -6189 12286 -6133
rect 12310 -6189 12366 -6133
rect 15531 -6189 15587 -6133
rect 15611 -6189 15667 -6133
rect 15691 -6189 15747 -6133
rect 916 -6632 972 -6576
rect 996 -6632 1052 -6576
rect 1076 -6632 1132 -6576
rect 9331 -6632 9387 -6576
rect 9411 -6632 9467 -6576
rect 9491 -6632 9547 -6576
rect 9633 -6632 9689 -6576
rect 9713 -6632 9769 -6576
rect 9793 -6632 9849 -6576
rect 18048 -6632 18104 -6576
rect 18128 -6632 18184 -6576
rect 18208 -6632 18264 -6576
rect 4550 -6777 4606 -6721
rect 4630 -6777 4686 -6721
rect 4710 -6777 4766 -6721
rect 5697 -6777 5753 -6721
rect 5777 -6777 5833 -6721
rect 5857 -6777 5913 -6721
rect 13267 -6777 13323 -6721
rect 13347 -6777 13403 -6721
rect 13427 -6777 13483 -6721
rect 14414 -6777 14470 -6721
rect 14494 -6777 14550 -6721
rect 14574 -6777 14630 -6721
rect 1338 -6938 1394 -6882
rect 1418 -6938 1474 -6882
rect 1498 -6938 1554 -6882
rect 8908 -6938 8964 -6882
rect 8988 -6938 9044 -6882
rect 9068 -6938 9124 -6882
rect 10056 -6938 10112 -6882
rect 10136 -6938 10192 -6882
rect 10216 -6938 10272 -6882
rect 17626 -6938 17682 -6882
rect 17706 -6938 17762 -6882
rect 17786 -6938 17842 -6882
rect 4985 -7078 5041 -7022
rect 5065 -7078 5121 -7022
rect 5145 -7078 5201 -7022
rect 5262 -7078 5318 -7022
rect 5342 -7078 5398 -7022
rect 5422 -7078 5478 -7022
rect 13702 -7078 13758 -7022
rect 13782 -7078 13838 -7022
rect 13862 -7078 13918 -7022
rect 13979 -7078 14035 -7022
rect 14059 -7078 14115 -7022
rect 14139 -7078 14195 -7022
rect 3433 -7516 3489 -7460
rect 3513 -7516 3569 -7460
rect 3593 -7516 3649 -7460
rect 6814 -7516 6870 -7460
rect 6894 -7516 6950 -7460
rect 6974 -7516 7030 -7460
rect 12150 -7516 12206 -7460
rect 12230 -7516 12286 -7460
rect 12310 -7516 12366 -7460
rect 15531 -7516 15587 -7460
rect 15611 -7516 15667 -7460
rect 15691 -7516 15747 -7460
rect 2465 -7836 2521 -7780
rect 2545 -7836 2601 -7780
rect 2625 -7836 2681 -7780
rect 7782 -7836 7838 -7780
rect 7862 -7836 7918 -7780
rect 7942 -7836 7998 -7780
rect 11182 -7836 11238 -7780
rect 11262 -7836 11318 -7780
rect 11342 -7836 11398 -7780
rect 16499 -7836 16555 -7780
rect 16579 -7836 16635 -7780
rect 16659 -7836 16715 -7780
rect 1338 -8267 1394 -8211
rect 1418 -8267 1474 -8211
rect 1498 -8267 1554 -8211
rect 8908 -8267 8964 -8211
rect 8988 -8267 9044 -8211
rect 9068 -8267 9124 -8211
rect 10056 -8267 10112 -8211
rect 10136 -8267 10192 -8211
rect 10216 -8267 10272 -8211
rect 17626 -8267 17682 -8211
rect 17706 -8267 17762 -8211
rect 17786 -8267 17842 -8211
rect 4550 -8436 4606 -8380
rect 4630 -8436 4686 -8380
rect 4710 -8436 4766 -8380
rect 5697 -8436 5753 -8380
rect 5777 -8436 5833 -8380
rect 5857 -8436 5913 -8380
rect 13267 -8436 13323 -8380
rect 13347 -8436 13403 -8380
rect 13427 -8436 13483 -8380
rect 14414 -8436 14470 -8380
rect 14494 -8436 14550 -8380
rect 14574 -8436 14630 -8380
rect 916 -8599 972 -8543
rect 996 -8599 1052 -8543
rect 1076 -8599 1132 -8543
rect 9331 -8599 9387 -8543
rect 9411 -8599 9467 -8543
rect 9491 -8599 9547 -8543
rect 9633 -8599 9689 -8543
rect 9713 -8599 9769 -8543
rect 9793 -8599 9849 -8543
rect 18048 -8599 18104 -8543
rect 18128 -8599 18184 -8543
rect 18208 -8599 18264 -8543
rect 4985 -8767 5041 -8711
rect 5065 -8767 5121 -8711
rect 5145 -8767 5201 -8711
rect 5262 -8767 5318 -8711
rect 5342 -8767 5398 -8711
rect 5422 -8767 5478 -8711
rect 13702 -8767 13758 -8711
rect 13782 -8767 13838 -8711
rect 13862 -8767 13918 -8711
rect 13979 -8767 14035 -8711
rect 14059 -8767 14115 -8711
rect 14139 -8767 14195 -8711
<< metal3 >>
rect 4941 4 5522 26
rect 4941 -52 4985 4
rect 5041 -52 5065 4
rect 5121 -52 5145 4
rect 5201 -52 5262 4
rect 5318 -52 5342 4
rect 5398 -52 5422 4
rect 5478 -52 5522 4
rect 876 -165 1176 -143
rect 876 -221 916 -165
rect 972 -221 996 -165
rect 1052 -221 1076 -165
rect 1132 -221 1176 -165
rect 876 -2131 1176 -221
rect 4506 -328 4806 -306
rect 4506 -384 4550 -328
rect 4606 -384 4630 -328
rect 4686 -384 4710 -328
rect 4766 -384 4806 -328
rect 876 -2187 916 -2131
rect 972 -2187 996 -2131
rect 1052 -2187 1076 -2131
rect 1132 -2187 1176 -2131
rect 876 -3669 1176 -2187
rect 876 -3725 916 -3669
rect 972 -3725 996 -3669
rect 1052 -3725 1076 -3669
rect 1132 -3725 1176 -3669
rect 876 -5038 1176 -3725
rect 876 -5094 916 -5038
rect 972 -5094 996 -5038
rect 1052 -5094 1076 -5038
rect 1132 -5094 1176 -5038
rect 876 -6576 1176 -5094
rect 876 -6632 916 -6576
rect 972 -6632 996 -6576
rect 1052 -6632 1076 -6576
rect 1132 -6632 1176 -6576
rect 876 -8543 1176 -6632
rect 1298 -496 1598 -474
rect 1298 -552 1338 -496
rect 1394 -552 1418 -496
rect 1474 -552 1498 -496
rect 1554 -552 1598 -496
rect 1298 -1826 1598 -552
rect 1298 -1882 1338 -1826
rect 1394 -1882 1418 -1826
rect 1474 -1882 1498 -1826
rect 1554 -1882 1598 -1826
rect 1298 -3338 1598 -1882
rect 1298 -3394 1338 -3338
rect 1394 -3394 1418 -3338
rect 1474 -3394 1498 -3338
rect 1554 -3394 1598 -3338
rect 1298 -5370 1598 -3394
rect 1298 -5426 1338 -5370
rect 1394 -5426 1418 -5370
rect 1474 -5426 1498 -5370
rect 1554 -5426 1598 -5370
rect 1298 -6882 1598 -5426
rect 1298 -6938 1338 -6882
rect 1394 -6938 1418 -6882
rect 1474 -6938 1498 -6882
rect 1554 -6938 1598 -6882
rect 1298 -8211 1598 -6938
rect 2425 -928 2725 -906
rect 2425 -984 2465 -928
rect 2521 -984 2545 -928
rect 2601 -984 2625 -928
rect 2681 -984 2725 -928
rect 2425 -2907 2725 -984
rect 2425 -2963 2465 -2907
rect 2521 -2963 2545 -2907
rect 2601 -2963 2625 -2907
rect 2681 -2963 2725 -2907
rect 2425 -5801 2725 -2963
rect 2425 -5857 2465 -5801
rect 2521 -5857 2545 -5801
rect 2601 -5857 2625 -5801
rect 2681 -5857 2725 -5801
rect 2425 -7780 2725 -5857
rect 3393 -1248 3693 -1226
rect 3393 -1304 3433 -1248
rect 3489 -1304 3513 -1248
rect 3569 -1304 3593 -1248
rect 3649 -1304 3693 -1248
rect 3393 -2575 3693 -1304
rect 3393 -2631 3433 -2575
rect 3489 -2631 3513 -2575
rect 3569 -2631 3593 -2575
rect 3649 -2631 3693 -2575
rect 3393 -6133 3693 -2631
rect 3393 -6189 3433 -6133
rect 3489 -6189 3513 -6133
rect 3569 -6189 3593 -6133
rect 3649 -6189 3693 -6133
rect 3393 -7460 3693 -6189
rect 3393 -7516 3433 -7460
rect 3489 -7516 3513 -7460
rect 3569 -7516 3593 -7460
rect 3649 -7516 3693 -7460
rect 3393 -7538 3693 -7516
rect 4506 -1987 4806 -384
rect 4506 -2043 4550 -1987
rect 4606 -2043 4630 -1987
rect 4686 -2043 4710 -1987
rect 4766 -2043 4806 -1987
rect 4506 -3507 4806 -2043
rect 4506 -3563 4550 -3507
rect 4606 -3563 4630 -3507
rect 4686 -3563 4710 -3507
rect 4766 -3563 4806 -3507
rect 4506 -5201 4806 -3563
rect 4506 -5257 4550 -5201
rect 4606 -5257 4630 -5201
rect 4686 -5257 4710 -5201
rect 4766 -5257 4806 -5201
rect 4506 -6721 4806 -5257
rect 4506 -6777 4550 -6721
rect 4606 -6777 4630 -6721
rect 4686 -6777 4710 -6721
rect 4766 -6777 4806 -6721
rect 2425 -7836 2465 -7780
rect 2521 -7836 2545 -7780
rect 2601 -7836 2625 -7780
rect 2681 -7836 2725 -7780
rect 2425 -7858 2725 -7836
rect 1298 -8267 1338 -8211
rect 1394 -8267 1418 -8211
rect 1474 -8267 1498 -8211
rect 1554 -8267 1598 -8211
rect 1298 -8289 1598 -8267
rect 4506 -8380 4806 -6777
rect 4506 -8436 4550 -8380
rect 4606 -8436 4630 -8380
rect 4686 -8436 4710 -8380
rect 4766 -8436 4806 -8380
rect 4506 -8458 4806 -8436
rect 4941 -1686 5522 -52
rect 13658 4 14239 26
rect 13658 -52 13702 4
rect 13758 -52 13782 4
rect 13838 -52 13862 4
rect 13918 -52 13979 4
rect 14035 -52 14059 4
rect 14115 -52 14139 4
rect 14195 -52 14239 4
rect 9287 -165 9893 -143
rect 9287 -221 9331 -165
rect 9387 -221 9411 -165
rect 9467 -221 9491 -165
rect 9547 -221 9633 -165
rect 9689 -221 9713 -165
rect 9769 -221 9793 -165
rect 9849 -221 9893 -165
rect 4941 -1742 4985 -1686
rect 5041 -1742 5065 -1686
rect 5121 -1742 5145 -1686
rect 5201 -1742 5262 -1686
rect 5318 -1742 5342 -1686
rect 5398 -1742 5422 -1686
rect 5478 -1742 5522 -1686
rect 4941 -3838 5522 -1742
rect 4941 -3894 4985 -3838
rect 5041 -3894 5065 -3838
rect 5121 -3894 5145 -3838
rect 5201 -3894 5262 -3838
rect 5318 -3894 5342 -3838
rect 5398 -3894 5422 -3838
rect 5478 -3894 5522 -3838
rect 4941 -4869 5522 -3894
rect 4941 -4925 4985 -4869
rect 5041 -4925 5065 -4869
rect 5121 -4925 5145 -4869
rect 5201 -4925 5262 -4869
rect 5318 -4925 5342 -4869
rect 5398 -4925 5422 -4869
rect 5478 -4925 5522 -4869
rect 4941 -7022 5522 -4925
rect 4941 -7078 4985 -7022
rect 5041 -7078 5065 -7022
rect 5121 -7078 5145 -7022
rect 5201 -7078 5262 -7022
rect 5318 -7078 5342 -7022
rect 5398 -7078 5422 -7022
rect 5478 -7078 5522 -7022
rect 876 -8599 916 -8543
rect 972 -8599 996 -8543
rect 1052 -8599 1076 -8543
rect 1132 -8599 1176 -8543
rect 876 -8621 1176 -8599
rect 4941 -8711 5522 -7078
rect 5657 -328 5957 -306
rect 5657 -384 5697 -328
rect 5753 -384 5777 -328
rect 5833 -384 5857 -328
rect 5913 -384 5957 -328
rect 5657 -1987 5957 -384
rect 8864 -496 9164 -474
rect 8864 -552 8908 -496
rect 8964 -552 8988 -496
rect 9044 -552 9068 -496
rect 9124 -552 9164 -496
rect 7738 -928 8038 -906
rect 7738 -984 7782 -928
rect 7838 -984 7862 -928
rect 7918 -984 7942 -928
rect 7998 -984 8038 -928
rect 5657 -2043 5697 -1987
rect 5753 -2043 5777 -1987
rect 5833 -2043 5857 -1987
rect 5913 -2043 5957 -1987
rect 5657 -3507 5957 -2043
rect 5657 -3563 5697 -3507
rect 5753 -3563 5777 -3507
rect 5833 -3563 5857 -3507
rect 5913 -3563 5957 -3507
rect 5657 -5201 5957 -3563
rect 5657 -5257 5697 -5201
rect 5753 -5257 5777 -5201
rect 5833 -5257 5857 -5201
rect 5913 -5257 5957 -5201
rect 5657 -6721 5957 -5257
rect 5657 -6777 5697 -6721
rect 5753 -6777 5777 -6721
rect 5833 -6777 5857 -6721
rect 5913 -6777 5957 -6721
rect 5657 -8380 5957 -6777
rect 6770 -1248 7070 -1226
rect 6770 -1304 6814 -1248
rect 6870 -1304 6894 -1248
rect 6950 -1304 6974 -1248
rect 7030 -1304 7070 -1248
rect 6770 -2586 7070 -1304
rect 6770 -2642 6814 -2586
rect 6870 -2642 6894 -2586
rect 6950 -2642 6974 -2586
rect 7030 -2642 7070 -2586
rect 6770 -6133 7070 -2642
rect 6770 -6189 6814 -6133
rect 6870 -6189 6894 -6133
rect 6950 -6189 6974 -6133
rect 7030 -6189 7070 -6133
rect 6770 -7460 7070 -6189
rect 6770 -7516 6814 -7460
rect 6870 -7516 6894 -7460
rect 6950 -7516 6974 -7460
rect 7030 -7516 7070 -7460
rect 6770 -7538 7070 -7516
rect 7738 -2907 8038 -984
rect 7738 -2963 7782 -2907
rect 7838 -2963 7862 -2907
rect 7918 -2963 7942 -2907
rect 7998 -2963 8038 -2907
rect 7738 -5801 8038 -2963
rect 7738 -5857 7782 -5801
rect 7838 -5857 7862 -5801
rect 7918 -5857 7942 -5801
rect 7998 -5857 8038 -5801
rect 7738 -7780 8038 -5857
rect 7738 -7836 7782 -7780
rect 7838 -7836 7862 -7780
rect 7918 -7836 7942 -7780
rect 7998 -7836 8038 -7780
rect 7738 -7858 8038 -7836
rect 8864 -1826 9164 -552
rect 8864 -1882 8908 -1826
rect 8964 -1882 8988 -1826
rect 9044 -1882 9068 -1826
rect 9124 -1882 9164 -1826
rect 8864 -3338 9164 -1882
rect 8864 -3394 8908 -3338
rect 8964 -3394 8988 -3338
rect 9044 -3394 9068 -3338
rect 9124 -3394 9164 -3338
rect 8864 -5370 9164 -3394
rect 8864 -5426 8908 -5370
rect 8964 -5426 8988 -5370
rect 9044 -5426 9068 -5370
rect 9124 -5426 9164 -5370
rect 8864 -6882 9164 -5426
rect 8864 -6938 8908 -6882
rect 8964 -6938 8988 -6882
rect 9044 -6938 9068 -6882
rect 9124 -6938 9164 -6882
rect 8864 -8211 9164 -6938
rect 8864 -8267 8908 -8211
rect 8964 -8267 8988 -8211
rect 9044 -8267 9068 -8211
rect 9124 -8267 9164 -8211
rect 8864 -8289 9164 -8267
rect 9287 -2131 9893 -221
rect 13223 -328 13523 -306
rect 13223 -384 13267 -328
rect 13323 -384 13347 -328
rect 13403 -384 13427 -328
rect 13483 -384 13523 -328
rect 9287 -2187 9331 -2131
rect 9387 -2187 9411 -2131
rect 9467 -2187 9491 -2131
rect 9547 -2187 9633 -2131
rect 9689 -2187 9713 -2131
rect 9769 -2187 9793 -2131
rect 9849 -2187 9893 -2131
rect 9287 -3669 9893 -2187
rect 9287 -3725 9331 -3669
rect 9387 -3725 9411 -3669
rect 9467 -3725 9491 -3669
rect 9547 -3725 9633 -3669
rect 9689 -3725 9713 -3669
rect 9769 -3725 9793 -3669
rect 9849 -3725 9893 -3669
rect 9287 -5038 9893 -3725
rect 9287 -5094 9331 -5038
rect 9387 -5094 9411 -5038
rect 9467 -5094 9491 -5038
rect 9547 -5094 9633 -5038
rect 9689 -5094 9713 -5038
rect 9769 -5094 9793 -5038
rect 9849 -5094 9893 -5038
rect 9287 -6576 9893 -5094
rect 9287 -6632 9331 -6576
rect 9387 -6632 9411 -6576
rect 9467 -6632 9491 -6576
rect 9547 -6632 9633 -6576
rect 9689 -6632 9713 -6576
rect 9769 -6632 9793 -6576
rect 9849 -6632 9893 -6576
rect 5657 -8436 5697 -8380
rect 5753 -8436 5777 -8380
rect 5833 -8436 5857 -8380
rect 5913 -8436 5957 -8380
rect 5657 -8458 5957 -8436
rect 9287 -8543 9893 -6632
rect 10016 -496 10316 -474
rect 10016 -552 10056 -496
rect 10112 -552 10136 -496
rect 10192 -552 10216 -496
rect 10272 -552 10316 -496
rect 10016 -1826 10316 -552
rect 10016 -1882 10056 -1826
rect 10112 -1882 10136 -1826
rect 10192 -1882 10216 -1826
rect 10272 -1882 10316 -1826
rect 10016 -3338 10316 -1882
rect 10016 -3394 10056 -3338
rect 10112 -3394 10136 -3338
rect 10192 -3394 10216 -3338
rect 10272 -3394 10316 -3338
rect 10016 -5370 10316 -3394
rect 10016 -5426 10056 -5370
rect 10112 -5426 10136 -5370
rect 10192 -5426 10216 -5370
rect 10272 -5426 10316 -5370
rect 10016 -6882 10316 -5426
rect 10016 -6938 10056 -6882
rect 10112 -6938 10136 -6882
rect 10192 -6938 10216 -6882
rect 10272 -6938 10316 -6882
rect 10016 -8211 10316 -6938
rect 11142 -928 11442 -906
rect 11142 -984 11182 -928
rect 11238 -984 11262 -928
rect 11318 -984 11342 -928
rect 11398 -984 11442 -928
rect 11142 -2907 11442 -984
rect 11142 -2963 11182 -2907
rect 11238 -2963 11262 -2907
rect 11318 -2963 11342 -2907
rect 11398 -2963 11442 -2907
rect 11142 -5801 11442 -2963
rect 11142 -5857 11182 -5801
rect 11238 -5857 11262 -5801
rect 11318 -5857 11342 -5801
rect 11398 -5857 11442 -5801
rect 11142 -7780 11442 -5857
rect 12110 -1248 12410 -1226
rect 12110 -1304 12150 -1248
rect 12206 -1304 12230 -1248
rect 12286 -1304 12310 -1248
rect 12366 -1304 12410 -1248
rect 12110 -2586 12410 -1304
rect 12110 -2642 12150 -2586
rect 12206 -2642 12230 -2586
rect 12286 -2642 12310 -2586
rect 12366 -2642 12410 -2586
rect 12110 -6133 12410 -2642
rect 12110 -6189 12150 -6133
rect 12206 -6189 12230 -6133
rect 12286 -6189 12310 -6133
rect 12366 -6189 12410 -6133
rect 12110 -7460 12410 -6189
rect 12110 -7516 12150 -7460
rect 12206 -7516 12230 -7460
rect 12286 -7516 12310 -7460
rect 12366 -7516 12410 -7460
rect 12110 -7538 12410 -7516
rect 13223 -1987 13523 -384
rect 13223 -2043 13267 -1987
rect 13323 -2043 13347 -1987
rect 13403 -2043 13427 -1987
rect 13483 -2043 13523 -1987
rect 13223 -3507 13523 -2043
rect 13223 -3563 13267 -3507
rect 13323 -3563 13347 -3507
rect 13403 -3563 13427 -3507
rect 13483 -3563 13523 -3507
rect 13223 -5201 13523 -3563
rect 13223 -5257 13267 -5201
rect 13323 -5257 13347 -5201
rect 13403 -5257 13427 -5201
rect 13483 -5257 13523 -5201
rect 13223 -6721 13523 -5257
rect 13223 -6777 13267 -6721
rect 13323 -6777 13347 -6721
rect 13403 -6777 13427 -6721
rect 13483 -6777 13523 -6721
rect 11142 -7836 11182 -7780
rect 11238 -7836 11262 -7780
rect 11318 -7836 11342 -7780
rect 11398 -7836 11442 -7780
rect 11142 -7858 11442 -7836
rect 10016 -8267 10056 -8211
rect 10112 -8267 10136 -8211
rect 10192 -8267 10216 -8211
rect 10272 -8267 10316 -8211
rect 10016 -8289 10316 -8267
rect 13223 -8380 13523 -6777
rect 13223 -8436 13267 -8380
rect 13323 -8436 13347 -8380
rect 13403 -8436 13427 -8380
rect 13483 -8436 13523 -8380
rect 13223 -8458 13523 -8436
rect 13658 -1686 14239 -52
rect 18004 -165 18304 -143
rect 18004 -221 18048 -165
rect 18104 -221 18128 -165
rect 18184 -221 18208 -165
rect 18264 -221 18304 -165
rect 13658 -1742 13702 -1686
rect 13758 -1742 13782 -1686
rect 13838 -1742 13862 -1686
rect 13918 -1742 13979 -1686
rect 14035 -1742 14059 -1686
rect 14115 -1742 14139 -1686
rect 14195 -1742 14239 -1686
rect 13658 -3838 14239 -1742
rect 13658 -3894 13702 -3838
rect 13758 -3894 13782 -3838
rect 13838 -3894 13862 -3838
rect 13918 -3894 13979 -3838
rect 14035 -3894 14059 -3838
rect 14115 -3894 14139 -3838
rect 14195 -3894 14239 -3838
rect 13658 -4869 14239 -3894
rect 13658 -4925 13702 -4869
rect 13758 -4925 13782 -4869
rect 13838 -4925 13862 -4869
rect 13918 -4925 13979 -4869
rect 14035 -4925 14059 -4869
rect 14115 -4925 14139 -4869
rect 14195 -4925 14239 -4869
rect 13658 -7022 14239 -4925
rect 13658 -7078 13702 -7022
rect 13758 -7078 13782 -7022
rect 13838 -7078 13862 -7022
rect 13918 -7078 13979 -7022
rect 14035 -7078 14059 -7022
rect 14115 -7078 14139 -7022
rect 14195 -7078 14239 -7022
rect 9287 -8599 9331 -8543
rect 9387 -8599 9411 -8543
rect 9467 -8599 9491 -8543
rect 9547 -8599 9633 -8543
rect 9689 -8599 9713 -8543
rect 9769 -8599 9793 -8543
rect 9849 -8599 9893 -8543
rect 9287 -8621 9893 -8599
rect 4941 -8767 4985 -8711
rect 5041 -8767 5065 -8711
rect 5121 -8767 5145 -8711
rect 5201 -8767 5262 -8711
rect 5318 -8767 5342 -8711
rect 5398 -8767 5422 -8711
rect 5478 -8767 5522 -8711
rect 4941 -8789 5522 -8767
rect 13658 -8711 14239 -7078
rect 14374 -328 14674 -306
rect 14374 -384 14414 -328
rect 14470 -384 14494 -328
rect 14550 -384 14574 -328
rect 14630 -384 14674 -328
rect 14374 -1987 14674 -384
rect 17582 -496 17882 -474
rect 17582 -552 17626 -496
rect 17682 -552 17706 -496
rect 17762 -552 17786 -496
rect 17842 -552 17882 -496
rect 16455 -928 16755 -906
rect 16455 -984 16499 -928
rect 16555 -984 16579 -928
rect 16635 -984 16659 -928
rect 16715 -984 16755 -928
rect 14374 -2043 14414 -1987
rect 14470 -2043 14494 -1987
rect 14550 -2043 14574 -1987
rect 14630 -2043 14674 -1987
rect 14374 -3507 14674 -2043
rect 14374 -3563 14414 -3507
rect 14470 -3563 14494 -3507
rect 14550 -3563 14574 -3507
rect 14630 -3563 14674 -3507
rect 14374 -5201 14674 -3563
rect 14374 -5257 14414 -5201
rect 14470 -5257 14494 -5201
rect 14550 -5257 14574 -5201
rect 14630 -5257 14674 -5201
rect 14374 -6721 14674 -5257
rect 14374 -6777 14414 -6721
rect 14470 -6777 14494 -6721
rect 14550 -6777 14574 -6721
rect 14630 -6777 14674 -6721
rect 14374 -8380 14674 -6777
rect 15487 -1248 15787 -1226
rect 15487 -1304 15531 -1248
rect 15587 -1304 15611 -1248
rect 15667 -1304 15691 -1248
rect 15747 -1304 15787 -1248
rect 15487 -2575 15787 -1304
rect 15487 -2631 15531 -2575
rect 15587 -2631 15611 -2575
rect 15667 -2631 15691 -2575
rect 15747 -2631 15787 -2575
rect 15487 -6133 15787 -2631
rect 15487 -6189 15531 -6133
rect 15587 -6189 15611 -6133
rect 15667 -6189 15691 -6133
rect 15747 -6189 15787 -6133
rect 15487 -7460 15787 -6189
rect 15487 -7516 15531 -7460
rect 15587 -7516 15611 -7460
rect 15667 -7516 15691 -7460
rect 15747 -7516 15787 -7460
rect 15487 -7538 15787 -7516
rect 16455 -2907 16755 -984
rect 16455 -2963 16499 -2907
rect 16555 -2963 16579 -2907
rect 16635 -2963 16659 -2907
rect 16715 -2963 16755 -2907
rect 16455 -5801 16755 -2963
rect 16455 -5857 16499 -5801
rect 16555 -5857 16579 -5801
rect 16635 -5857 16659 -5801
rect 16715 -5857 16755 -5801
rect 16455 -7780 16755 -5857
rect 16455 -7836 16499 -7780
rect 16555 -7836 16579 -7780
rect 16635 -7836 16659 -7780
rect 16715 -7836 16755 -7780
rect 16455 -7858 16755 -7836
rect 17582 -1826 17882 -552
rect 17582 -1882 17626 -1826
rect 17682 -1882 17706 -1826
rect 17762 -1882 17786 -1826
rect 17842 -1882 17882 -1826
rect 17582 -3338 17882 -1882
rect 17582 -3394 17626 -3338
rect 17682 -3394 17706 -3338
rect 17762 -3394 17786 -3338
rect 17842 -3394 17882 -3338
rect 17582 -5370 17882 -3394
rect 17582 -5426 17626 -5370
rect 17682 -5426 17706 -5370
rect 17762 -5426 17786 -5370
rect 17842 -5426 17882 -5370
rect 17582 -6882 17882 -5426
rect 17582 -6938 17626 -6882
rect 17682 -6938 17706 -6882
rect 17762 -6938 17786 -6882
rect 17842 -6938 17882 -6882
rect 17582 -8211 17882 -6938
rect 17582 -8267 17626 -8211
rect 17682 -8267 17706 -8211
rect 17762 -8267 17786 -8211
rect 17842 -8267 17882 -8211
rect 17582 -8289 17882 -8267
rect 18004 -2131 18304 -221
rect 18004 -2187 18048 -2131
rect 18104 -2187 18128 -2131
rect 18184 -2187 18208 -2131
rect 18264 -2187 18304 -2131
rect 18004 -3669 18304 -2187
rect 18004 -3725 18048 -3669
rect 18104 -3725 18128 -3669
rect 18184 -3725 18208 -3669
rect 18264 -3725 18304 -3669
rect 18004 -5038 18304 -3725
rect 18004 -5094 18048 -5038
rect 18104 -5094 18128 -5038
rect 18184 -5094 18208 -5038
rect 18264 -5094 18304 -5038
rect 18004 -6576 18304 -5094
rect 18004 -6632 18048 -6576
rect 18104 -6632 18128 -6576
rect 18184 -6632 18208 -6576
rect 18264 -6632 18304 -6576
rect 14374 -8436 14414 -8380
rect 14470 -8436 14494 -8380
rect 14550 -8436 14574 -8380
rect 14630 -8436 14674 -8380
rect 14374 -8458 14674 -8436
rect 18004 -8543 18304 -6632
rect 18004 -8599 18048 -8543
rect 18104 -8599 18128 -8543
rect 18184 -8599 18208 -8543
rect 18264 -8599 18304 -8543
rect 18004 -8621 18304 -8599
rect 13658 -8767 13702 -8711
rect 13758 -8767 13782 -8711
rect 13838 -8767 13862 -8711
rect 13918 -8767 13979 -8711
rect 14035 -8767 14059 -8711
rect 14115 -8767 14139 -8711
rect 14195 -8767 14239 -8711
rect 13658 -8789 14239 -8767
<< end >>
