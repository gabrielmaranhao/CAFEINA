* NGSPICE file created from esd_structure.ext - technology: sky130A

.subckt esd_structure VDD VSS PAD GATE
D0 VSS.t5 PAD.t1 sky130_fd_pr__diode_pw2nd_11v0 pj=2.2e+07 area=1e+13
D1 GATE.t1 VDD.t0 sky130_fd_pr__diode_pd2nw_05v5 pj=1.8e+06 area=2.025e+11
D2 VSS.t4 PAD.t2 sky130_fd_pr__diode_pw2nd_11v0 pj=2.2e+07 area=1e+13
D3 PAD.t3 VDD.t5 sky130_fd_pr__diode_pd2nw_11v0 pj=2.2e+07 area=1e+13
D4 PAD.t4 VDD.t4 sky130_fd_pr__diode_pd2nw_11v0 pj=2.2e+07 area=1e+13
D5 VSS.t3 PAD.t5 sky130_fd_pr__diode_pw2nd_11v0 pj=2.2e+07 area=1e+13
D6 VSS.t0 GATE.t2 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
D7 PAD.t6 VDD.t3 sky130_fd_pr__diode_pd2nw_11v0 pj=2.2e+07 area=1e+13
D8 VSS.t2 PAD.t7 sky130_fd_pr__diode_pw2nd_11v0 pj=2.2e+07 area=1e+13
D9 VSS.t1 PAD.t8 sky130_fd_pr__diode_pw2nd_11v0 pj=2.2e+07 area=1e+13
D10 PAD.t9 VDD.t2 sky130_fd_pr__diode_pd2nw_11v0 pj=2.2e+07 area=1e+13
D11 PAD.t10 VDD.t1 sky130_fd_pr__diode_pd2nw_11v0 pj=2.2e+07 area=1e+13
X0 GATE PAD VSS.t6 sky130_fd_pr__res_high_po_0p35 l=10
R0 PAD.n1 PAD.t10 7.88381
R1 PAD.n4 PAD.t9 7.88381
R2 PAD.n0 PAD.t4 7.86996
R3 PAD.n2 PAD.t6 7.86996
R4 PAD.n3 PAD.t3 7.85667
R5 PAD.n3 PAD.t8 3.12876
R6 PAD.n4 PAD.t7 3.08886
R7 PAD.n2 PAD.t1 3.08268
R8 PAD.n1 PAD.t2 3.03726
R9 PAD.n0 PAD.t5 2.98039
R10 PAD PAD.n4 0.496594
R11 PAD.n2 PAD.n1 0.335321
R12 PAD.n3 PAD.n2 0.335321
R13 PAD.n1 PAD.n0 0.330857
R14 PAD.n4 PAD.n3 0.328625
R15 VSS.n60 VSS.n59 41845.4
R16 VSS.n60 VSS.n58 37037.8
R17 VSS.n84 VSS.n29 9710.94
R18 VSS.n94 VSS.n29 9710.94
R19 VSS.n84 VSS.n30 9710.94
R20 VSS.n94 VSS.n30 9710.94
R21 VSS.n53 VSS.n52 9513.78
R22 VSS.n61 VSS.n52 9513.78
R23 VSS.n54 VSS.n53 9513.78
R24 VSS.n61 VSS.n54 9513.78
R25 VSS.n59 VSS.n6 8944.64
R26 VSS.n58 VSS.n55 8226.36
R27 VSS.n125 VSS.n3 4231.64
R28 VSS.n125 VSS.n4 4231.64
R29 VSS.n126 VSS.n4 4231.64
R30 VSS.n126 VSS.n3 4231.64
R31 VSS.n120 VSS.n9 4231.64
R32 VSS.n120 VSS.n10 4231.64
R33 VSS.n117 VSS.n10 4231.64
R34 VSS.n117 VSS.n9 4231.64
R35 VSS.n111 VSS.n13 4231.64
R36 VSS.n112 VSS.n13 4231.64
R37 VSS.n112 VSS.n15 4231.64
R38 VSS.n111 VSS.n15 4231.64
R39 VSS.n107 VSS.n21 4231.64
R40 VSS.n106 VSS.n21 4231.64
R41 VSS.n106 VSS.n20 4231.64
R42 VSS.n107 VSS.n20 4231.64
R43 VSS.n100 VSS.n28 4231.64
R44 VSS.n101 VSS.n28 4231.64
R45 VSS.n101 VSS.n27 4231.64
R46 VSS.n100 VSS.n27 4231.64
R47 VSS.n56 VSS.n40 3657.19
R48 VSS.n79 VSS.n37 3007.15
R49 VSS.n87 VSS.n37 3007.15
R50 VSS.n87 VSS.n38 3007.15
R51 VSS.n79 VSS.n38 3007.15
R52 VSS.n78 VSS.n77 2840.43
R53 VSS.n78 VSS.n39 2715.27
R54 VSS.n76 VSS.n44 1407.97
R55 VSS.n45 VSS.n44 1407.97
R56 VSS.n76 VSS.n47 1407.97
R57 VSS.n47 VSS.n45 1407.97
R58 VSS.n73 VSS.n48 1242.12
R59 VSS.n62 VSS.n51 1092.14
R60 VSS.n49 VSS.n32 1090.26
R61 VSS.n63 VSS.n62 859.838
R62 VSS.n92 VSS.n32 797.26
R63 VSS.n96 VSS.n95 771.23
R64 VSS.n86 VSS.n85 608.38
R65 VSS.n104 VSS.n103 602.678
R66 VSS.n57 VSS.n56 600.646
R67 VSS.n34 VSS.n33 563.201
R68 VSS.n91 VSS.n34 512.63
R69 VSS.n124 VSS.n2 488.283
R70 VSS.n127 VSS.n2 488.283
R71 VSS.n121 VSS.n8 488.283
R72 VSS.n102 VSS.n26 488.283
R73 VSS.n99 VSS.n26 488.283
R74 VSS.n108 VSS.n19 464.377
R75 VSS.n104 VSS.n24 392.178
R76 VSS.n58 VSS.n57 355.413
R77 VSS.t3 VSS.n96 318.017
R78 VSS.t3 VSS.n97 318.017
R79 VSS.t4 VSS.n22 318.017
R80 VSS.t4 VSS.n23 318.017
R81 VSS.t5 VSS.n16 318.017
R82 VSS.t1 VSS.n118 318.017
R83 VSS.n119 VSS.t1 318.017
R84 VSS.t2 VSS.n5 318.017
R85 VSS.t2 VSS.n6 318.017
R86 VSS.n97 VSS.n22 310.336
R87 VSS.n23 VSS.n16 310.336
R88 VSS.n118 VSS.n11 310.336
R89 VSS.n119 VSS.n5 310.336
R90 VSS.n17 VSS.n11 302.654
R91 VSS.n45 VSS.n41 292.5
R92 VSS.n46 VSS.n45 292.5
R93 VSS.n47 VSS.n42 292.5
R94 VSS.n47 VSS.t0 292.5
R95 VSS.n76 VSS.n75 292.5
R96 VSS.n77 VSS.n76 292.5
R97 VSS.n74 VSS.n44 292.5
R98 VSS.t0 VSS.n44 292.5
R99 VSS.n48 VSS.n29 292.5
R100 VSS.n29 VSS.t6 292.5
R101 VSS.n90 VSS.n30 292.5
R102 VSS.n56 VSS.n30 292.5
R103 VSS.n55 VSS.n39 245.845
R104 VSS.t0 VSS.n46 237.739
R105 VSS.n95 VSS.t6 227.375
R106 VSS.n77 VSS.n43 223.109
R107 VSS.n92 VSS.n33 212.978
R108 VSS.n85 VSS.n40 212.012
R109 VSS.n63 VSS.n50 204.089
R110 VSS.n80 VSS.n35 195.388
R111 VSS.n100 VSS.n99 146.25
R112 VSS.t3 VSS.n100 146.25
R113 VSS.n102 VSS.n101 146.25
R114 VSS.n101 VSS.t3 146.25
R115 VSS.n108 VSS.n107 146.25
R116 VSS.n107 VSS.t4 146.25
R117 VSS.n106 VSS.n105 146.25
R118 VSS.t4 VSS.n106 146.25
R119 VSS.n111 VSS.n110 146.25
R120 VSS.t5 VSS.n111 146.25
R121 VSS.n113 VSS.n112 146.25
R122 VSS.n112 VSS.t5 146.25
R123 VSS.n9 VSS.n7 146.25
R124 VSS.t1 VSS.n9 146.25
R125 VSS.n10 VSS.n8 146.25
R126 VSS.t1 VSS.n10 146.25
R127 VSS.n127 VSS.n126 146.25
R128 VSS.n126 VSS.t2 146.25
R129 VSS.n125 VSS.n124 146.25
R130 VSS.t2 VSS.n125 146.25
R131 VSS.n99 VSS.n98 141.423
R132 VSS.n128 VSS.n127 141.169
R133 VSS.n86 VSS.n39 130.588
R134 VSS.n48 VSS.n31 123.504
R135 VSS.n90 VSS.n89 120.712
R136 VSS.n81 VSS.n80 108.171
R137 VSS.n81 VSS.n37 104.344
R138 VSS.n80 VSS.n79 97.5005
R139 VSS.n79 VSS.n78 97.5005
R140 VSS.n43 VSS.n37 97.5005
R141 VSS.n38 VSS.n35 97.5005
R142 VSS.n55 VSS.n38 97.5005
R143 VSS.n88 VSS.n87 97.5005
R144 VSS.n87 VSS.n86 97.5005
R145 VSS.n89 VSS.n35 94.4946
R146 VSS.n75 VSS.n74 91.4829
R147 VSS.n123 VSS.n7 90.8926
R148 VSS.n46 VSS.n39 82.2948
R149 VSS.n124 VSS.n123 74.7894
R150 VSS.n105 VSS.n14 71.5299
R151 VSS.n110 VSS.n109 71.5299
R152 VSS.n110 VSS.n12 71.5299
R153 VSS.n12 VSS.n7 71.5299
R154 VSS.n114 VSS.n8 71.5299
R155 VSS.n113 VSS.n14 71.5299
R156 VSS.n114 VSS.n113 71.5299
R157 VSS.n109 VSS.n108 71.5299
R158 VSS.n103 VSS.n102 71.5299
R159 VSS.n105 VSS.n104 70.777
R160 VSS.n103 VSS.n25 69.0698
R161 VSS.n116 VSS.n12 60.0412
R162 VSS.n109 VSS.n18 60.0412
R163 VSS.n67 VSS.n14 59.6073
R164 VSS.n115 VSS.n114 58.9564
R165 VSS.n123 VSS.n122 56.8726
R166 VSS.n50 VSS.n33 53.6894
R167 VSS.n91 VSS.n90 49.3181
R168 VSS.n93 VSS.n92 47.3101
R169 VSS.n75 VSS.n42 43.3786
R170 VSS.n64 VSS.n63 42.9823
R171 VSS.n74 VSS.n73 42.5417
R172 VSS.n93 VSS.n31 32.1381
R173 VSS.n92 VSS.n91 21.4941
R174 VSS.n27 VSS.n26 19.5005
R175 VSS.n96 VSS.n27 19.5005
R176 VSS.n98 VSS.n28 19.5005
R177 VSS.n97 VSS.n28 19.5005
R178 VSS.n20 VSS.n19 19.5005
R179 VSS.n22 VSS.n20 19.5005
R180 VSS.n21 VSS.n18 19.5005
R181 VSS.n23 VSS.n21 19.5005
R182 VSS.n18 VSS.n15 19.5005
R183 VSS.n16 VSS.n15 19.5005
R184 VSS.n116 VSS.n13 19.5005
R185 VSS.n13 VSS.n11 19.5005
R186 VSS.n117 VSS.n116 19.5005
R187 VSS.n118 VSS.n117 19.5005
R188 VSS.n121 VSS.n120 19.5005
R189 VSS.n120 VSS.n119 19.5005
R190 VSS.n3 VSS.n1 19.5005
R191 VSS.n5 VSS.n3 19.5005
R192 VSS.n4 VSS.n2 19.5005
R193 VSS.n6 VSS.n4 19.5005
R194 VSS.n54 VSS.n51 16.2505
R195 VSS.n59 VSS.n54 16.2505
R196 VSS.n52 VSS.n50 16.2505
R197 VSS.n57 VSS.n52 16.2505
R198 VSS.t5 VSS.n17 15.3636
R199 VSS.n40 VSS.t6 15.236
R200 VSS.t0 VSS.n43 14.6306
R201 VSS.n94 VSS.n93 13.6052
R202 VSS.n95 VSS.n94 13.6052
R203 VSS.n84 VSS.n83 13.6052
R204 VSS.n85 VSS.n84 13.6052
R205 VSS.n62 VSS.n61 13.0005
R206 VSS.n61 VSS.n60 13.0005
R207 VSS.n53 VSS.n32 13.0005
R208 VSS.n53 VSS.n17 13.0005
R209 VSS.n64 VSS.n34 9.67323
R210 VSS.n89 VSS.n88 7.97817
R211 VSS.n82 VSS.n42 7.08973
R212 VSS.n82 VSS.n41 6.26336
R213 VSS.n83 VSS.n36 5.1205
R214 VSS.n65 VSS.n49 4.21093
R215 VSS.n83 VSS.n82 3.97817
R216 VSS.n73 VSS.n72 2.69764
R217 VSS.n122 VSS.n121 2.63579
R218 VSS.n71 VSS.n31 2.3005
R219 VSS.n88 VSS.n36 2.05445
R220 VSS.n51 VSS.n49 1.88285
R221 VSS.n24 VSS.n19 1.42272
R222 VSS.n66 VSS.n36 1.40956
R223 VSS.n72 VSS.n71 1.18164
R224 VSS.n66 VSS.n65 1.1131
R225 VSS.n116 VSS.n115 0.922534
R226 VSS.n25 VSS.n24 0.824262
R227 VSS.n69 VSS.n25 0.461815
R228 VSS.n68 VSS.n67 0.461815
R229 VSS.n115 VSS.n0 0.461815
R230 VSS.n129 VSS.n128 0.461815
R231 VSS.n122 VSS.n1 0.444064
R232 VSS.n72 VSS.n41 0.274786
R233 VSS.n67 VSS.n18 0.271686
R234 VSS.n98 VSS.n24 0.253965
R235 VSS.n82 VSS.n81 0.246654
R236 VSS.n65 VSS.n64 0.133357
R237 VSS.n128 VSS.n1 0.0638663
R238 VSS.n70 VSS.n66 0.0637184
R239 VSS VSS.n129 0.0630545
R240 VSS.n71 VSS.n70 0.0496247
R241 VSS.n70 VSS.n69 0.0416399
R242 VSS.n129 VSS.n0 0.0343928
R243 VSS.n69 VSS.n68 0.0342838
R244 VSS.n68 VSS.n0 0.0336299
R245 GATE.n0 GATE.t1 594.694
R246 GATE.n0 GATE.t2 194.549
R247 GATE GATE.n0 0.230151
R248 VDD.n64 VDD.n9 2509.97
R249 VDD.n63 VDD.n9 2509.97
R250 VDD.n63 VDD.n8 2509.97
R251 VDD.n64 VDD.n8 2509.97
R252 VDD.n59 VDD.n10 2509.97
R253 VDD.n59 VDD.n11 2509.97
R254 VDD.n38 VDD.n11 2509.97
R255 VDD.n38 VDD.n10 2509.97
R256 VDD.n43 VDD.n37 2509.97
R257 VDD.n43 VDD.n42 2509.97
R258 VDD.n41 VDD.n37 2509.97
R259 VDD.n42 VDD.n41 2509.97
R260 VDD.n31 VDD.n30 2509.97
R261 VDD.n46 VDD.n31 2509.97
R262 VDD.n47 VDD.n46 2509.97
R263 VDD.n68 VDD.n5 2509.97
R264 VDD.n70 VDD.n4 2509.97
R265 VDD.n68 VDD.n4 2509.97
R266 VDD.n23 VDD.n22 857.648
R267 VDD.n20 VDD.n18 857.648
R268 VDD.n48 VDD.n28 485.272
R269 VDD.n32 VDD.n28 485.272
R270 VDD.n67 VDD.n3 485.272
R271 VDD.n71 VDD.n3 485.272
R272 VDD.n23 VDD.n17 267.182
R273 VDD.n21 VDD.n20 267.182
R274 VDD.n18 VDD.n15 92.5005
R275 VDD.n20 VDD.n19 92.5005
R276 VDD.n22 VDD.n16 92.5005
R277 VDD.n24 VDD.n23 92.5005
R278 VDD.n30 VDD.n29 82.2983
R279 VDD.n69 VDD.n5 82.2983
R280 VDD.n45 VDD.t4 80.4888
R281 VDD.n44 VDD.t1 80.4888
R282 VDD.n40 VDD.t1 80.4888
R283 VDD.n39 VDD.t3 80.4888
R284 VDD.n60 VDD.t3 80.4888
R285 VDD.t5 VDD.n61 80.4888
R286 VDD.t5 VDD.n62 80.4888
R287 VDD.t2 VDD.n6 80.4888
R288 VDD.n45 VDD.n44 75.3344
R289 VDD.n40 VDD.n39 75.3344
R290 VDD.n61 VDD.n60 75.3344
R291 VDD.n62 VDD.n6 75.3344
R292 VDD.n65 VDD.n7 70.024
R293 VDD.n66 VDD.n65 70.024
R294 VDD.n35 VDD.n34 70.024
R295 VDD.n49 VDD.n12 70.024
R296 VDD.n54 VDD.n12 70.024
R297 VDD.n67 VDD.n66 70.024
R298 VDD.n72 VDD.n71 70.024
R299 VDD.n56 VDD.n2 70.024
R300 VDD.n72 VDD.n2 70.024
R301 VDD.n55 VDD.n54 70.024
R302 VDD.n36 VDD.n33 70.024
R303 VDD.n36 VDD.n35 70.024
R304 VDD.n34 VDD.n7 68.5181
R305 VDD.n49 VDD.n48 68.5181
R306 VDD.n56 VDD.n55 68.5181
R307 VDD.n33 VDD.n32 68.5181
R308 VDD.n66 VDD.n1 63.0291
R309 VDD.n35 VDD.n13 63.0291
R310 VDD.n73 VDD.n72 62.7434
R311 VDD.n58 VDD.n7 61.9233
R312 VDD.n33 VDD.n27 61.9233
R313 VDD.n57 VDD.n56 61.5303
R314 VDD.n50 VDD.n49 61.5303
R315 VDD.n54 VDD.n53 61.3719
R316 VDD.n25 VDD.n15 60.593
R317 VDD.n18 VDD.n17 57.4849
R318 VDD.n22 VDD.n21 57.4849
R319 VDD.n15 VDD.n14 55.4189
R320 VDD.n48 VDD.n47 46.2505
R321 VDD.n42 VDD.n12 46.2505
R322 VDD.n42 VDD.t1 46.2505
R323 VDD.n34 VDD.n10 46.2505
R324 VDD.n10 VDD.t3 46.2505
R325 VDD.n65 VDD.n64 46.2505
R326 VDD.n64 VDD.t5 46.2505
R327 VDD.n68 VDD.n67 46.2505
R328 VDD.t2 VDD.n68 46.2505
R329 VDD.n71 VDD.n70 46.2505
R330 VDD.n63 VDD.n2 46.2505
R331 VDD.t5 VDD.n63 46.2505
R332 VDD.n55 VDD.n11 46.2505
R333 VDD.n11 VDD.t3 46.2505
R334 VDD.n37 VDD.n36 46.2505
R335 VDD.n37 VDD.t1 46.2505
R336 VDD.n32 VDD.n31 46.2505
R337 VDD.t4 VDD.n31 46.2505
R338 VDD.n47 VDD.n29 43.9252
R339 VDD.n70 VDD.n69 43.9252
R340 VDD.n24 VDD.n16 43.0241
R341 VDD.n19 VDD.n16 40.9441
R342 VDD.n21 VDD.t0 28.8172
R343 VDD.t0 VDD.n17 28.8172
R344 VDD.n30 VDD.n28 6.16717
R345 VDD.n5 VDD.n3 6.16717
R346 VDD.n9 VDD.n1 6.16717
R347 VDD.n62 VDD.n9 6.16717
R348 VDD.n4 VDD.n1 6.16717
R349 VDD.n6 VDD.n4 6.16717
R350 VDD.n59 VDD.n58 6.16717
R351 VDD.n60 VDD.n59 6.16717
R352 VDD.n58 VDD.n8 6.16717
R353 VDD.n61 VDD.n8 6.16717
R354 VDD.n41 VDD.n13 6.16717
R355 VDD.n41 VDD.n40 6.16717
R356 VDD.n38 VDD.n13 6.16717
R357 VDD.n39 VDD.n38 6.16717
R358 VDD.n46 VDD.n27 6.16717
R359 VDD.n46 VDD.n45 6.16717
R360 VDD.n43 VDD.n27 6.16717
R361 VDD.n44 VDD.n43 6.16717
R362 VDD.n19 VDD.n14 3.93896
R363 VDD.n25 VDD.n24 3.28255
R364 VDD.n26 VDD.n14 2.77474
R365 VDD.n26 VDD.n25 2.7652
R366 VDD.n53 VDD.n13 1.54336
R367 VDD.n69 VDD.t2 1.51745
R368 VDD.t4 VDD.n29 1.51745
R369 VDD.n51 VDD.n26 1.47074
R370 VDD.n51 VDD.n50 0.461815
R371 VDD.n53 VDD.n52 0.461815
R372 VDD.n57 VDD.n0 0.461815
R373 VDD.n74 VDD.n73 0.461815
R374 VDD.n50 VDD.n27 0.393482
R375 VDD.n73 VDD.n1 0.171929
R376 VDD.n58 VDD.n57 0.168921
R377 VDD VDD.n74 0.0638174
R378 VDD.n52 VDD.n51 0.032976
R379 VDD.n52 VDD.n0 0.032976
R380 VDD.n74 VDD.n0 0.0327581
C0 VDD GATE 0.429f
C1 PAD GATE 0.113f
C2 VDD PAD 21.6f
.ends

