magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< nwell >>
rect 816 -8987 9679 813
<< pmoshvt >>
rect 1033 361 1233 561
rect 1485 361 1685 561
rect 1743 361 1943 561
rect 2001 361 2201 561
rect 2259 361 2459 561
rect 2711 361 2911 561
rect 2969 361 3169 561
rect 3227 361 3427 561
rect 3679 361 3879 561
rect 3937 361 4137 561
rect 4195 361 4395 561
rect 4453 361 4653 561
rect 4905 361 5105 561
rect 5391 361 5591 561
rect 5842 361 6042 561
rect 6100 361 6300 561
rect 6358 361 6558 561
rect 6616 361 6816 561
rect 7068 361 7268 561
rect 7326 361 7526 561
rect 7584 361 7784 561
rect 8036 361 8236 561
rect 8294 361 8494 561
rect 8552 361 8752 561
rect 8810 361 9010 561
rect 9262 361 9462 561
rect 1033 -583 1233 -383
rect 1485 -583 1685 -383
rect 1743 -583 1943 -383
rect 2001 -583 2201 -383
rect 2259 -583 2459 -383
rect 2711 -583 2911 -383
rect 2969 -583 3169 -383
rect 3227 -583 3427 -383
rect 3679 -583 3879 -383
rect 3937 -583 4137 -383
rect 4195 -583 4395 -383
rect 4453 -583 4653 -383
rect 4905 -583 5105 -383
rect 5391 -583 5591 -383
rect 5842 -583 6042 -383
rect 6100 -583 6300 -383
rect 6358 -583 6558 -383
rect 6616 -583 6816 -383
rect 7068 -583 7268 -383
rect 7326 -583 7526 -383
rect 7584 -583 7784 -383
rect 8036 -583 8236 -383
rect 8294 -583 8494 -383
rect 8552 -583 8752 -383
rect 8810 -583 9010 -383
rect 9262 -583 9462 -383
rect 1033 -1274 1233 -1074
rect 1485 -1274 1685 -1074
rect 1743 -1274 1943 -1074
rect 2001 -1274 2201 -1074
rect 2259 -1274 2459 -1074
rect 2711 -1274 2911 -1074
rect 2969 -1274 3169 -1074
rect 3227 -1274 3427 -1074
rect 3679 -1274 3879 -1074
rect 3937 -1274 4137 -1074
rect 4195 -1274 4395 -1074
rect 4453 -1274 4653 -1074
rect 4905 -1274 5105 -1074
rect 5391 -1274 5591 -1074
rect 5842 -1274 6042 -1074
rect 6100 -1274 6300 -1074
rect 6358 -1274 6558 -1074
rect 6616 -1274 6816 -1074
rect 7068 -1274 7268 -1074
rect 7326 -1274 7526 -1074
rect 7584 -1274 7784 -1074
rect 8036 -1274 8236 -1074
rect 8294 -1274 8494 -1074
rect 8552 -1274 8752 -1074
rect 8810 -1274 9010 -1074
rect 9262 -1274 9462 -1074
rect 1033 -2230 1233 -2030
rect 1485 -2230 1685 -2030
rect 1743 -2230 1943 -2030
rect 2001 -2230 2201 -2030
rect 2259 -2230 2459 -2030
rect 2711 -2230 2911 -2030
rect 2969 -2230 3169 -2030
rect 3227 -2230 3427 -2030
rect 3679 -2230 3879 -2030
rect 3937 -2230 4137 -2030
rect 4195 -2230 4395 -2030
rect 4453 -2230 4653 -2030
rect 4905 -2230 5105 -2030
rect 5391 -2230 5591 -2030
rect 5842 -2230 6042 -2030
rect 6100 -2230 6300 -2030
rect 6358 -2230 6558 -2030
rect 6616 -2230 6816 -2030
rect 7068 -2230 7268 -2030
rect 7326 -2230 7526 -2030
rect 7584 -2230 7784 -2030
rect 8036 -2230 8236 -2030
rect 8294 -2230 8494 -2030
rect 8552 -2230 8752 -2030
rect 8810 -2230 9010 -2030
rect 9262 -2230 9462 -2030
rect 1033 -2921 1233 -2721
rect 1485 -2921 1685 -2721
rect 1743 -2921 1943 -2721
rect 2001 -2921 2201 -2721
rect 2259 -2921 2459 -2721
rect 2711 -2921 2911 -2721
rect 2969 -2921 3169 -2721
rect 3227 -2921 3427 -2721
rect 3679 -2921 3879 -2721
rect 3937 -2921 4137 -2721
rect 4195 -2921 4395 -2721
rect 4453 -2921 4653 -2721
rect 4905 -2921 5105 -2721
rect 5391 -2921 5591 -2721
rect 5842 -2921 6042 -2721
rect 6100 -2921 6300 -2721
rect 6358 -2921 6558 -2721
rect 6616 -2921 6816 -2721
rect 7068 -2921 7268 -2721
rect 7326 -2921 7526 -2721
rect 7584 -2921 7784 -2721
rect 8036 -2921 8236 -2721
rect 8294 -2921 8494 -2721
rect 8552 -2921 8752 -2721
rect 8810 -2921 9010 -2721
rect 9262 -2921 9462 -2721
rect 1033 -3911 1233 -3711
rect 1485 -3911 1685 -3711
rect 1743 -3911 1943 -3711
rect 2001 -3911 2201 -3711
rect 2259 -3911 2459 -3711
rect 2711 -3911 2911 -3711
rect 2969 -3911 3169 -3711
rect 3227 -3911 3427 -3711
rect 3679 -3911 3879 -3711
rect 3937 -3911 4137 -3711
rect 4195 -3911 4395 -3711
rect 4453 -3911 4653 -3711
rect 4905 -3911 5105 -3711
rect 5391 -3911 5591 -3711
rect 5842 -3911 6042 -3711
rect 6100 -3911 6300 -3711
rect 6358 -3911 6558 -3711
rect 6616 -3911 6816 -3711
rect 7068 -3911 7268 -3711
rect 7326 -3911 7526 -3711
rect 7584 -3911 7784 -3711
rect 8036 -3911 8236 -3711
rect 8294 -3911 8494 -3711
rect 8552 -3911 8752 -3711
rect 8810 -3911 9010 -3711
rect 9262 -3911 9462 -3711
rect 1033 -4467 1233 -4267
rect 1485 -4467 1685 -4267
rect 1743 -4467 1943 -4267
rect 2001 -4467 2201 -4267
rect 2259 -4467 2459 -4267
rect 2711 -4467 2911 -4267
rect 2969 -4467 3169 -4267
rect 3227 -4467 3427 -4267
rect 3679 -4467 3879 -4267
rect 3937 -4467 4137 -4267
rect 4195 -4467 4395 -4267
rect 4453 -4467 4653 -4267
rect 4905 -4467 5105 -4267
rect 5391 -4467 5591 -4267
rect 5842 -4467 6042 -4267
rect 6100 -4467 6300 -4267
rect 6358 -4467 6558 -4267
rect 6616 -4467 6816 -4267
rect 7068 -4467 7268 -4267
rect 7326 -4467 7526 -4267
rect 7584 -4467 7784 -4267
rect 8036 -4467 8236 -4267
rect 8294 -4467 8494 -4267
rect 8552 -4467 8752 -4267
rect 8810 -4467 9010 -4267
rect 9262 -4467 9462 -4267
rect 1033 -5457 1233 -5257
rect 1485 -5457 1685 -5257
rect 1743 -5457 1943 -5257
rect 2001 -5457 2201 -5257
rect 2259 -5457 2459 -5257
rect 2711 -5457 2911 -5257
rect 2969 -5457 3169 -5257
rect 3227 -5457 3427 -5257
rect 3679 -5457 3879 -5257
rect 3937 -5457 4137 -5257
rect 4195 -5457 4395 -5257
rect 4453 -5457 4653 -5257
rect 4905 -5457 5105 -5257
rect 5391 -5457 5591 -5257
rect 5842 -5457 6042 -5257
rect 6100 -5457 6300 -5257
rect 6358 -5457 6558 -5257
rect 6616 -5457 6816 -5257
rect 7068 -5457 7268 -5257
rect 7326 -5457 7526 -5257
rect 7584 -5457 7784 -5257
rect 8036 -5457 8236 -5257
rect 8294 -5457 8494 -5257
rect 8552 -5457 8752 -5257
rect 8810 -5457 9010 -5257
rect 9262 -5457 9462 -5257
rect 1033 -6147 1233 -5947
rect 1485 -6147 1685 -5947
rect 1743 -6147 1943 -5947
rect 2001 -6147 2201 -5947
rect 2259 -6147 2459 -5947
rect 2711 -6147 2911 -5947
rect 2969 -6147 3169 -5947
rect 3227 -6147 3427 -5947
rect 3679 -6147 3879 -5947
rect 3937 -6147 4137 -5947
rect 4195 -6147 4395 -5947
rect 4453 -6147 4653 -5947
rect 4905 -6147 5105 -5947
rect 5391 -6147 5591 -5947
rect 5842 -6147 6042 -5947
rect 6100 -6147 6300 -5947
rect 6358 -6147 6558 -5947
rect 6616 -6147 6816 -5947
rect 7068 -6147 7268 -5947
rect 7326 -6147 7526 -5947
rect 7584 -6147 7784 -5947
rect 8036 -6147 8236 -5947
rect 8294 -6147 8494 -5947
rect 8552 -6147 8752 -5947
rect 8810 -6147 9010 -5947
rect 9262 -6147 9462 -5947
rect 1033 -7104 1233 -6904
rect 1485 -7104 1685 -6904
rect 1743 -7104 1943 -6904
rect 2001 -7104 2201 -6904
rect 2259 -7104 2459 -6904
rect 2711 -7104 2911 -6904
rect 2969 -7104 3169 -6904
rect 3227 -7104 3427 -6904
rect 3679 -7104 3879 -6904
rect 3937 -7104 4137 -6904
rect 4195 -7104 4395 -6904
rect 4453 -7104 4653 -6904
rect 4905 -7104 5105 -6904
rect 5391 -7104 5591 -6904
rect 5842 -7104 6042 -6904
rect 6100 -7104 6300 -6904
rect 6358 -7104 6558 -6904
rect 6616 -7104 6816 -6904
rect 7068 -7104 7268 -6904
rect 7326 -7104 7526 -6904
rect 7584 -7104 7784 -6904
rect 8036 -7104 8236 -6904
rect 8294 -7104 8494 -6904
rect 8552 -7104 8752 -6904
rect 8810 -7104 9010 -6904
rect 9262 -7104 9462 -6904
rect 1033 -7794 1233 -7594
rect 1485 -7794 1685 -7594
rect 1743 -7794 1943 -7594
rect 2001 -7794 2201 -7594
rect 2259 -7794 2459 -7594
rect 2711 -7794 2911 -7594
rect 2969 -7794 3169 -7594
rect 3227 -7794 3427 -7594
rect 3679 -7794 3879 -7594
rect 3937 -7794 4137 -7594
rect 4195 -7794 4395 -7594
rect 4453 -7794 4653 -7594
rect 4905 -7794 5105 -7594
rect 5391 -7794 5591 -7594
rect 5842 -7794 6042 -7594
rect 6100 -7794 6300 -7594
rect 6358 -7794 6558 -7594
rect 6616 -7794 6816 -7594
rect 7068 -7794 7268 -7594
rect 7326 -7794 7526 -7594
rect 7584 -7794 7784 -7594
rect 8036 -7794 8236 -7594
rect 8294 -7794 8494 -7594
rect 8552 -7794 8752 -7594
rect 8810 -7794 9010 -7594
rect 9262 -7794 9462 -7594
rect 1033 -8738 1233 -8538
rect 1485 -8738 1685 -8538
rect 1743 -8738 1943 -8538
rect 2001 -8738 2201 -8538
rect 2259 -8738 2459 -8538
rect 2711 -8738 2911 -8538
rect 2969 -8738 3169 -8538
rect 3227 -8738 3427 -8538
rect 3679 -8738 3879 -8538
rect 3937 -8738 4137 -8538
rect 4195 -8738 4395 -8538
rect 4453 -8738 4653 -8538
rect 4905 -8738 5105 -8538
rect 5391 -8738 5591 -8538
rect 5842 -8738 6042 -8538
rect 6100 -8738 6300 -8538
rect 6358 -8738 6558 -8538
rect 6616 -8738 6816 -8538
rect 7068 -8738 7268 -8538
rect 7326 -8738 7526 -8538
rect 7584 -8738 7784 -8538
rect 8036 -8738 8236 -8538
rect 8294 -8738 8494 -8538
rect 8552 -8738 8752 -8538
rect 8810 -8738 9010 -8538
rect 9262 -8738 9462 -8538
<< pdiff >>
rect 975 546 1033 561
rect 975 512 987 546
rect 1021 512 1033 546
rect 975 478 1033 512
rect 975 444 987 478
rect 1021 444 1033 478
rect 975 410 1033 444
rect 975 376 987 410
rect 1021 376 1033 410
rect 975 361 1033 376
rect 1233 546 1291 561
rect 1233 512 1245 546
rect 1279 512 1291 546
rect 1233 478 1291 512
rect 1233 444 1245 478
rect 1279 444 1291 478
rect 1233 410 1291 444
rect 1233 376 1245 410
rect 1279 376 1291 410
rect 1233 361 1291 376
rect 1427 546 1485 561
rect 1427 512 1439 546
rect 1473 512 1485 546
rect 1427 478 1485 512
rect 1427 444 1439 478
rect 1473 444 1485 478
rect 1427 410 1485 444
rect 1427 376 1439 410
rect 1473 376 1485 410
rect 1427 361 1485 376
rect 1685 546 1743 561
rect 1685 512 1697 546
rect 1731 512 1743 546
rect 1685 478 1743 512
rect 1685 444 1697 478
rect 1731 444 1743 478
rect 1685 410 1743 444
rect 1685 376 1697 410
rect 1731 376 1743 410
rect 1685 361 1743 376
rect 1943 546 2001 561
rect 1943 512 1955 546
rect 1989 512 2001 546
rect 1943 478 2001 512
rect 1943 444 1955 478
rect 1989 444 2001 478
rect 1943 410 2001 444
rect 1943 376 1955 410
rect 1989 376 2001 410
rect 1943 361 2001 376
rect 2201 546 2259 561
rect 2201 512 2213 546
rect 2247 512 2259 546
rect 2201 478 2259 512
rect 2201 444 2213 478
rect 2247 444 2259 478
rect 2201 410 2259 444
rect 2201 376 2213 410
rect 2247 376 2259 410
rect 2201 361 2259 376
rect 2459 546 2517 561
rect 2459 512 2471 546
rect 2505 512 2517 546
rect 2459 478 2517 512
rect 2459 444 2471 478
rect 2505 444 2517 478
rect 2459 410 2517 444
rect 2459 376 2471 410
rect 2505 376 2517 410
rect 2459 361 2517 376
rect 2653 546 2711 561
rect 2653 512 2665 546
rect 2699 512 2711 546
rect 2653 478 2711 512
rect 2653 444 2665 478
rect 2699 444 2711 478
rect 2653 410 2711 444
rect 2653 376 2665 410
rect 2699 376 2711 410
rect 2653 361 2711 376
rect 2911 546 2969 561
rect 2911 512 2923 546
rect 2957 512 2969 546
rect 2911 478 2969 512
rect 2911 444 2923 478
rect 2957 444 2969 478
rect 2911 410 2969 444
rect 2911 376 2923 410
rect 2957 376 2969 410
rect 2911 361 2969 376
rect 3169 546 3227 561
rect 3169 512 3181 546
rect 3215 512 3227 546
rect 3169 478 3227 512
rect 3169 444 3181 478
rect 3215 444 3227 478
rect 3169 410 3227 444
rect 3169 376 3181 410
rect 3215 376 3227 410
rect 3169 361 3227 376
rect 3427 546 3485 561
rect 3427 512 3439 546
rect 3473 512 3485 546
rect 3427 478 3485 512
rect 3427 444 3439 478
rect 3473 444 3485 478
rect 3427 410 3485 444
rect 3427 376 3439 410
rect 3473 376 3485 410
rect 3427 361 3485 376
rect 3621 546 3679 561
rect 3621 512 3633 546
rect 3667 512 3679 546
rect 3621 478 3679 512
rect 3621 444 3633 478
rect 3667 444 3679 478
rect 3621 410 3679 444
rect 3621 376 3633 410
rect 3667 376 3679 410
rect 3621 361 3679 376
rect 3879 546 3937 561
rect 3879 512 3891 546
rect 3925 512 3937 546
rect 3879 478 3937 512
rect 3879 444 3891 478
rect 3925 444 3937 478
rect 3879 410 3937 444
rect 3879 376 3891 410
rect 3925 376 3937 410
rect 3879 361 3937 376
rect 4137 546 4195 561
rect 4137 512 4149 546
rect 4183 512 4195 546
rect 4137 478 4195 512
rect 4137 444 4149 478
rect 4183 444 4195 478
rect 4137 410 4195 444
rect 4137 376 4149 410
rect 4183 376 4195 410
rect 4137 361 4195 376
rect 4395 546 4453 561
rect 4395 512 4407 546
rect 4441 512 4453 546
rect 4395 478 4453 512
rect 4395 444 4407 478
rect 4441 444 4453 478
rect 4395 410 4453 444
rect 4395 376 4407 410
rect 4441 376 4453 410
rect 4395 361 4453 376
rect 4653 546 4711 561
rect 4653 512 4665 546
rect 4699 512 4711 546
rect 4653 478 4711 512
rect 4653 444 4665 478
rect 4699 444 4711 478
rect 4653 410 4711 444
rect 4653 376 4665 410
rect 4699 376 4711 410
rect 4653 361 4711 376
rect 4847 546 4905 561
rect 4847 512 4859 546
rect 4893 512 4905 546
rect 4847 478 4905 512
rect 4847 444 4859 478
rect 4893 444 4905 478
rect 4847 410 4905 444
rect 4847 376 4859 410
rect 4893 376 4905 410
rect 4847 361 4905 376
rect 5105 546 5163 561
rect 5105 512 5117 546
rect 5151 512 5163 546
rect 5105 478 5163 512
rect 5105 444 5117 478
rect 5151 444 5163 478
rect 5105 410 5163 444
rect 5105 376 5117 410
rect 5151 376 5163 410
rect 5105 361 5163 376
rect 5333 546 5391 561
rect 5333 512 5345 546
rect 5379 512 5391 546
rect 5333 478 5391 512
rect 5333 444 5345 478
rect 5379 444 5391 478
rect 5333 410 5391 444
rect 5333 376 5345 410
rect 5379 376 5391 410
rect 5333 361 5391 376
rect 5591 546 5649 561
rect 5591 512 5603 546
rect 5637 512 5649 546
rect 5591 478 5649 512
rect 5591 444 5603 478
rect 5637 444 5649 478
rect 5591 410 5649 444
rect 5591 376 5603 410
rect 5637 376 5649 410
rect 5591 361 5649 376
rect 5784 546 5842 561
rect 5784 512 5796 546
rect 5830 512 5842 546
rect 5784 478 5842 512
rect 5784 444 5796 478
rect 5830 444 5842 478
rect 5784 410 5842 444
rect 5784 376 5796 410
rect 5830 376 5842 410
rect 5784 361 5842 376
rect 6042 546 6100 561
rect 6042 512 6054 546
rect 6088 512 6100 546
rect 6042 478 6100 512
rect 6042 444 6054 478
rect 6088 444 6100 478
rect 6042 410 6100 444
rect 6042 376 6054 410
rect 6088 376 6100 410
rect 6042 361 6100 376
rect 6300 546 6358 561
rect 6300 512 6312 546
rect 6346 512 6358 546
rect 6300 478 6358 512
rect 6300 444 6312 478
rect 6346 444 6358 478
rect 6300 410 6358 444
rect 6300 376 6312 410
rect 6346 376 6358 410
rect 6300 361 6358 376
rect 6558 546 6616 561
rect 6558 512 6570 546
rect 6604 512 6616 546
rect 6558 478 6616 512
rect 6558 444 6570 478
rect 6604 444 6616 478
rect 6558 410 6616 444
rect 6558 376 6570 410
rect 6604 376 6616 410
rect 6558 361 6616 376
rect 6816 546 6874 561
rect 6816 512 6828 546
rect 6862 512 6874 546
rect 6816 478 6874 512
rect 6816 444 6828 478
rect 6862 444 6874 478
rect 6816 410 6874 444
rect 6816 376 6828 410
rect 6862 376 6874 410
rect 6816 361 6874 376
rect 7010 546 7068 561
rect 7010 512 7022 546
rect 7056 512 7068 546
rect 7010 478 7068 512
rect 7010 444 7022 478
rect 7056 444 7068 478
rect 7010 410 7068 444
rect 7010 376 7022 410
rect 7056 376 7068 410
rect 7010 361 7068 376
rect 7268 546 7326 561
rect 7268 512 7280 546
rect 7314 512 7326 546
rect 7268 478 7326 512
rect 7268 444 7280 478
rect 7314 444 7326 478
rect 7268 410 7326 444
rect 7268 376 7280 410
rect 7314 376 7326 410
rect 7268 361 7326 376
rect 7526 546 7584 561
rect 7526 512 7538 546
rect 7572 512 7584 546
rect 7526 478 7584 512
rect 7526 444 7538 478
rect 7572 444 7584 478
rect 7526 410 7584 444
rect 7526 376 7538 410
rect 7572 376 7584 410
rect 7526 361 7584 376
rect 7784 546 7842 561
rect 7784 512 7796 546
rect 7830 512 7842 546
rect 7784 478 7842 512
rect 7784 444 7796 478
rect 7830 444 7842 478
rect 7784 410 7842 444
rect 7784 376 7796 410
rect 7830 376 7842 410
rect 7784 361 7842 376
rect 7978 546 8036 561
rect 7978 512 7990 546
rect 8024 512 8036 546
rect 7978 478 8036 512
rect 7978 444 7990 478
rect 8024 444 8036 478
rect 7978 410 8036 444
rect 7978 376 7990 410
rect 8024 376 8036 410
rect 7978 361 8036 376
rect 8236 546 8294 561
rect 8236 512 8248 546
rect 8282 512 8294 546
rect 8236 478 8294 512
rect 8236 444 8248 478
rect 8282 444 8294 478
rect 8236 410 8294 444
rect 8236 376 8248 410
rect 8282 376 8294 410
rect 8236 361 8294 376
rect 8494 546 8552 561
rect 8494 512 8506 546
rect 8540 512 8552 546
rect 8494 478 8552 512
rect 8494 444 8506 478
rect 8540 444 8552 478
rect 8494 410 8552 444
rect 8494 376 8506 410
rect 8540 376 8552 410
rect 8494 361 8552 376
rect 8752 546 8810 561
rect 8752 512 8764 546
rect 8798 512 8810 546
rect 8752 478 8810 512
rect 8752 444 8764 478
rect 8798 444 8810 478
rect 8752 410 8810 444
rect 8752 376 8764 410
rect 8798 376 8810 410
rect 8752 361 8810 376
rect 9010 546 9068 561
rect 9010 512 9022 546
rect 9056 512 9068 546
rect 9010 478 9068 512
rect 9010 444 9022 478
rect 9056 444 9068 478
rect 9010 410 9068 444
rect 9010 376 9022 410
rect 9056 376 9068 410
rect 9010 361 9068 376
rect 9204 546 9262 561
rect 9204 512 9216 546
rect 9250 512 9262 546
rect 9204 478 9262 512
rect 9204 444 9216 478
rect 9250 444 9262 478
rect 9204 410 9262 444
rect 9204 376 9216 410
rect 9250 376 9262 410
rect 9204 361 9262 376
rect 9462 546 9520 561
rect 9462 512 9474 546
rect 9508 512 9520 546
rect 9462 478 9520 512
rect 9462 444 9474 478
rect 9508 444 9520 478
rect 9462 410 9520 444
rect 9462 376 9474 410
rect 9508 376 9520 410
rect 9462 361 9520 376
rect 975 -398 1033 -383
rect 975 -432 987 -398
rect 1021 -432 1033 -398
rect 975 -466 1033 -432
rect 975 -500 987 -466
rect 1021 -500 1033 -466
rect 975 -534 1033 -500
rect 975 -568 987 -534
rect 1021 -568 1033 -534
rect 975 -583 1033 -568
rect 1233 -398 1291 -383
rect 1233 -432 1245 -398
rect 1279 -432 1291 -398
rect 1233 -466 1291 -432
rect 1233 -500 1245 -466
rect 1279 -500 1291 -466
rect 1233 -534 1291 -500
rect 1233 -568 1245 -534
rect 1279 -568 1291 -534
rect 1233 -583 1291 -568
rect 1427 -398 1485 -383
rect 1427 -432 1439 -398
rect 1473 -432 1485 -398
rect 1427 -466 1485 -432
rect 1427 -500 1439 -466
rect 1473 -500 1485 -466
rect 1427 -534 1485 -500
rect 1427 -568 1439 -534
rect 1473 -568 1485 -534
rect 1427 -583 1485 -568
rect 1685 -398 1743 -383
rect 1685 -432 1697 -398
rect 1731 -432 1743 -398
rect 1685 -466 1743 -432
rect 1685 -500 1697 -466
rect 1731 -500 1743 -466
rect 1685 -534 1743 -500
rect 1685 -568 1697 -534
rect 1731 -568 1743 -534
rect 1685 -583 1743 -568
rect 1943 -398 2001 -383
rect 1943 -432 1955 -398
rect 1989 -432 2001 -398
rect 1943 -466 2001 -432
rect 1943 -500 1955 -466
rect 1989 -500 2001 -466
rect 1943 -534 2001 -500
rect 1943 -568 1955 -534
rect 1989 -568 2001 -534
rect 1943 -583 2001 -568
rect 2201 -398 2259 -383
rect 2201 -432 2213 -398
rect 2247 -432 2259 -398
rect 2201 -466 2259 -432
rect 2201 -500 2213 -466
rect 2247 -500 2259 -466
rect 2201 -534 2259 -500
rect 2201 -568 2213 -534
rect 2247 -568 2259 -534
rect 2201 -583 2259 -568
rect 2459 -398 2517 -383
rect 2459 -432 2471 -398
rect 2505 -432 2517 -398
rect 2459 -466 2517 -432
rect 2459 -500 2471 -466
rect 2505 -500 2517 -466
rect 2459 -534 2517 -500
rect 2459 -568 2471 -534
rect 2505 -568 2517 -534
rect 2459 -583 2517 -568
rect 2653 -398 2711 -383
rect 2653 -432 2665 -398
rect 2699 -432 2711 -398
rect 2653 -466 2711 -432
rect 2653 -500 2665 -466
rect 2699 -500 2711 -466
rect 2653 -534 2711 -500
rect 2653 -568 2665 -534
rect 2699 -568 2711 -534
rect 2653 -583 2711 -568
rect 2911 -398 2969 -383
rect 2911 -432 2923 -398
rect 2957 -432 2969 -398
rect 2911 -466 2969 -432
rect 2911 -500 2923 -466
rect 2957 -500 2969 -466
rect 2911 -534 2969 -500
rect 2911 -568 2923 -534
rect 2957 -568 2969 -534
rect 2911 -583 2969 -568
rect 3169 -398 3227 -383
rect 3169 -432 3181 -398
rect 3215 -432 3227 -398
rect 3169 -466 3227 -432
rect 3169 -500 3181 -466
rect 3215 -500 3227 -466
rect 3169 -534 3227 -500
rect 3169 -568 3181 -534
rect 3215 -568 3227 -534
rect 3169 -583 3227 -568
rect 3427 -398 3485 -383
rect 3427 -432 3439 -398
rect 3473 -432 3485 -398
rect 3427 -466 3485 -432
rect 3427 -500 3439 -466
rect 3473 -500 3485 -466
rect 3427 -534 3485 -500
rect 3427 -568 3439 -534
rect 3473 -568 3485 -534
rect 3427 -583 3485 -568
rect 3621 -398 3679 -383
rect 3621 -432 3633 -398
rect 3667 -432 3679 -398
rect 3621 -466 3679 -432
rect 3621 -500 3633 -466
rect 3667 -500 3679 -466
rect 3621 -534 3679 -500
rect 3621 -568 3633 -534
rect 3667 -568 3679 -534
rect 3621 -583 3679 -568
rect 3879 -398 3937 -383
rect 3879 -432 3891 -398
rect 3925 -432 3937 -398
rect 3879 -466 3937 -432
rect 3879 -500 3891 -466
rect 3925 -500 3937 -466
rect 3879 -534 3937 -500
rect 3879 -568 3891 -534
rect 3925 -568 3937 -534
rect 3879 -583 3937 -568
rect 4137 -398 4195 -383
rect 4137 -432 4149 -398
rect 4183 -432 4195 -398
rect 4137 -466 4195 -432
rect 4137 -500 4149 -466
rect 4183 -500 4195 -466
rect 4137 -534 4195 -500
rect 4137 -568 4149 -534
rect 4183 -568 4195 -534
rect 4137 -583 4195 -568
rect 4395 -398 4453 -383
rect 4395 -432 4407 -398
rect 4441 -432 4453 -398
rect 4395 -466 4453 -432
rect 4395 -500 4407 -466
rect 4441 -500 4453 -466
rect 4395 -534 4453 -500
rect 4395 -568 4407 -534
rect 4441 -568 4453 -534
rect 4395 -583 4453 -568
rect 4653 -398 4711 -383
rect 4653 -432 4665 -398
rect 4699 -432 4711 -398
rect 4653 -466 4711 -432
rect 4653 -500 4665 -466
rect 4699 -500 4711 -466
rect 4653 -534 4711 -500
rect 4653 -568 4665 -534
rect 4699 -568 4711 -534
rect 4653 -583 4711 -568
rect 4847 -398 4905 -383
rect 4847 -432 4859 -398
rect 4893 -432 4905 -398
rect 4847 -466 4905 -432
rect 4847 -500 4859 -466
rect 4893 -500 4905 -466
rect 4847 -534 4905 -500
rect 4847 -568 4859 -534
rect 4893 -568 4905 -534
rect 4847 -583 4905 -568
rect 5105 -398 5163 -383
rect 5105 -432 5117 -398
rect 5151 -432 5163 -398
rect 5105 -466 5163 -432
rect 5105 -500 5117 -466
rect 5151 -500 5163 -466
rect 5105 -534 5163 -500
rect 5105 -568 5117 -534
rect 5151 -568 5163 -534
rect 5105 -583 5163 -568
rect 5333 -398 5391 -383
rect 5333 -432 5345 -398
rect 5379 -432 5391 -398
rect 5333 -466 5391 -432
rect 5333 -500 5345 -466
rect 5379 -500 5391 -466
rect 5333 -534 5391 -500
rect 5333 -568 5345 -534
rect 5379 -568 5391 -534
rect 5333 -583 5391 -568
rect 5591 -398 5649 -383
rect 5591 -432 5603 -398
rect 5637 -432 5649 -398
rect 5591 -466 5649 -432
rect 5591 -500 5603 -466
rect 5637 -500 5649 -466
rect 5591 -534 5649 -500
rect 5591 -568 5603 -534
rect 5637 -568 5649 -534
rect 5591 -583 5649 -568
rect 5784 -398 5842 -383
rect 5784 -432 5796 -398
rect 5830 -432 5842 -398
rect 5784 -466 5842 -432
rect 5784 -500 5796 -466
rect 5830 -500 5842 -466
rect 5784 -534 5842 -500
rect 5784 -568 5796 -534
rect 5830 -568 5842 -534
rect 5784 -583 5842 -568
rect 6042 -398 6100 -383
rect 6042 -432 6054 -398
rect 6088 -432 6100 -398
rect 6042 -466 6100 -432
rect 6042 -500 6054 -466
rect 6088 -500 6100 -466
rect 6042 -534 6100 -500
rect 6042 -568 6054 -534
rect 6088 -568 6100 -534
rect 6042 -583 6100 -568
rect 6300 -398 6358 -383
rect 6300 -432 6312 -398
rect 6346 -432 6358 -398
rect 6300 -466 6358 -432
rect 6300 -500 6312 -466
rect 6346 -500 6358 -466
rect 6300 -534 6358 -500
rect 6300 -568 6312 -534
rect 6346 -568 6358 -534
rect 6300 -583 6358 -568
rect 6558 -398 6616 -383
rect 6558 -432 6570 -398
rect 6604 -432 6616 -398
rect 6558 -466 6616 -432
rect 6558 -500 6570 -466
rect 6604 -500 6616 -466
rect 6558 -534 6616 -500
rect 6558 -568 6570 -534
rect 6604 -568 6616 -534
rect 6558 -583 6616 -568
rect 6816 -398 6874 -383
rect 6816 -432 6828 -398
rect 6862 -432 6874 -398
rect 6816 -466 6874 -432
rect 6816 -500 6828 -466
rect 6862 -500 6874 -466
rect 6816 -534 6874 -500
rect 6816 -568 6828 -534
rect 6862 -568 6874 -534
rect 6816 -583 6874 -568
rect 7010 -398 7068 -383
rect 7010 -432 7022 -398
rect 7056 -432 7068 -398
rect 7010 -466 7068 -432
rect 7010 -500 7022 -466
rect 7056 -500 7068 -466
rect 7010 -534 7068 -500
rect 7010 -568 7022 -534
rect 7056 -568 7068 -534
rect 7010 -583 7068 -568
rect 7268 -398 7326 -383
rect 7268 -432 7280 -398
rect 7314 -432 7326 -398
rect 7268 -466 7326 -432
rect 7268 -500 7280 -466
rect 7314 -500 7326 -466
rect 7268 -534 7326 -500
rect 7268 -568 7280 -534
rect 7314 -568 7326 -534
rect 7268 -583 7326 -568
rect 7526 -398 7584 -383
rect 7526 -432 7538 -398
rect 7572 -432 7584 -398
rect 7526 -466 7584 -432
rect 7526 -500 7538 -466
rect 7572 -500 7584 -466
rect 7526 -534 7584 -500
rect 7526 -568 7538 -534
rect 7572 -568 7584 -534
rect 7526 -583 7584 -568
rect 7784 -398 7842 -383
rect 7784 -432 7796 -398
rect 7830 -432 7842 -398
rect 7784 -466 7842 -432
rect 7784 -500 7796 -466
rect 7830 -500 7842 -466
rect 7784 -534 7842 -500
rect 7784 -568 7796 -534
rect 7830 -568 7842 -534
rect 7784 -583 7842 -568
rect 7978 -398 8036 -383
rect 7978 -432 7990 -398
rect 8024 -432 8036 -398
rect 7978 -466 8036 -432
rect 7978 -500 7990 -466
rect 8024 -500 8036 -466
rect 7978 -534 8036 -500
rect 7978 -568 7990 -534
rect 8024 -568 8036 -534
rect 7978 -583 8036 -568
rect 8236 -398 8294 -383
rect 8236 -432 8248 -398
rect 8282 -432 8294 -398
rect 8236 -466 8294 -432
rect 8236 -500 8248 -466
rect 8282 -500 8294 -466
rect 8236 -534 8294 -500
rect 8236 -568 8248 -534
rect 8282 -568 8294 -534
rect 8236 -583 8294 -568
rect 8494 -398 8552 -383
rect 8494 -432 8506 -398
rect 8540 -432 8552 -398
rect 8494 -466 8552 -432
rect 8494 -500 8506 -466
rect 8540 -500 8552 -466
rect 8494 -534 8552 -500
rect 8494 -568 8506 -534
rect 8540 -568 8552 -534
rect 8494 -583 8552 -568
rect 8752 -398 8810 -383
rect 8752 -432 8764 -398
rect 8798 -432 8810 -398
rect 8752 -466 8810 -432
rect 8752 -500 8764 -466
rect 8798 -500 8810 -466
rect 8752 -534 8810 -500
rect 8752 -568 8764 -534
rect 8798 -568 8810 -534
rect 8752 -583 8810 -568
rect 9010 -398 9068 -383
rect 9010 -432 9022 -398
rect 9056 -432 9068 -398
rect 9010 -466 9068 -432
rect 9010 -500 9022 -466
rect 9056 -500 9068 -466
rect 9010 -534 9068 -500
rect 9010 -568 9022 -534
rect 9056 -568 9068 -534
rect 9010 -583 9068 -568
rect 9204 -398 9262 -383
rect 9204 -432 9216 -398
rect 9250 -432 9262 -398
rect 9204 -466 9262 -432
rect 9204 -500 9216 -466
rect 9250 -500 9262 -466
rect 9204 -534 9262 -500
rect 9204 -568 9216 -534
rect 9250 -568 9262 -534
rect 9204 -583 9262 -568
rect 9462 -398 9520 -383
rect 9462 -432 9474 -398
rect 9508 -432 9520 -398
rect 9462 -466 9520 -432
rect 9462 -500 9474 -466
rect 9508 -500 9520 -466
rect 9462 -534 9520 -500
rect 9462 -568 9474 -534
rect 9508 -568 9520 -534
rect 9462 -583 9520 -568
rect 975 -1089 1033 -1074
rect 975 -1123 987 -1089
rect 1021 -1123 1033 -1089
rect 975 -1157 1033 -1123
rect 975 -1191 987 -1157
rect 1021 -1191 1033 -1157
rect 975 -1225 1033 -1191
rect 975 -1259 987 -1225
rect 1021 -1259 1033 -1225
rect 975 -1274 1033 -1259
rect 1233 -1089 1291 -1074
rect 1233 -1123 1245 -1089
rect 1279 -1123 1291 -1089
rect 1233 -1157 1291 -1123
rect 1233 -1191 1245 -1157
rect 1279 -1191 1291 -1157
rect 1233 -1225 1291 -1191
rect 1233 -1259 1245 -1225
rect 1279 -1259 1291 -1225
rect 1233 -1274 1291 -1259
rect 1427 -1089 1485 -1074
rect 1427 -1123 1439 -1089
rect 1473 -1123 1485 -1089
rect 1427 -1157 1485 -1123
rect 1427 -1191 1439 -1157
rect 1473 -1191 1485 -1157
rect 1427 -1225 1485 -1191
rect 1427 -1259 1439 -1225
rect 1473 -1259 1485 -1225
rect 1427 -1274 1485 -1259
rect 1685 -1089 1743 -1074
rect 1685 -1123 1697 -1089
rect 1731 -1123 1743 -1089
rect 1685 -1157 1743 -1123
rect 1685 -1191 1697 -1157
rect 1731 -1191 1743 -1157
rect 1685 -1225 1743 -1191
rect 1685 -1259 1697 -1225
rect 1731 -1259 1743 -1225
rect 1685 -1274 1743 -1259
rect 1943 -1089 2001 -1074
rect 1943 -1123 1955 -1089
rect 1989 -1123 2001 -1089
rect 1943 -1157 2001 -1123
rect 1943 -1191 1955 -1157
rect 1989 -1191 2001 -1157
rect 1943 -1225 2001 -1191
rect 1943 -1259 1955 -1225
rect 1989 -1259 2001 -1225
rect 1943 -1274 2001 -1259
rect 2201 -1089 2259 -1074
rect 2201 -1123 2213 -1089
rect 2247 -1123 2259 -1089
rect 2201 -1157 2259 -1123
rect 2201 -1191 2213 -1157
rect 2247 -1191 2259 -1157
rect 2201 -1225 2259 -1191
rect 2201 -1259 2213 -1225
rect 2247 -1259 2259 -1225
rect 2201 -1274 2259 -1259
rect 2459 -1089 2517 -1074
rect 2459 -1123 2471 -1089
rect 2505 -1123 2517 -1089
rect 2459 -1157 2517 -1123
rect 2459 -1191 2471 -1157
rect 2505 -1191 2517 -1157
rect 2459 -1225 2517 -1191
rect 2459 -1259 2471 -1225
rect 2505 -1259 2517 -1225
rect 2459 -1274 2517 -1259
rect 2653 -1089 2711 -1074
rect 2653 -1123 2665 -1089
rect 2699 -1123 2711 -1089
rect 2653 -1157 2711 -1123
rect 2653 -1191 2665 -1157
rect 2699 -1191 2711 -1157
rect 2653 -1225 2711 -1191
rect 2653 -1259 2665 -1225
rect 2699 -1259 2711 -1225
rect 2653 -1274 2711 -1259
rect 2911 -1089 2969 -1074
rect 2911 -1123 2923 -1089
rect 2957 -1123 2969 -1089
rect 2911 -1157 2969 -1123
rect 2911 -1191 2923 -1157
rect 2957 -1191 2969 -1157
rect 2911 -1225 2969 -1191
rect 2911 -1259 2923 -1225
rect 2957 -1259 2969 -1225
rect 2911 -1274 2969 -1259
rect 3169 -1089 3227 -1074
rect 3169 -1123 3181 -1089
rect 3215 -1123 3227 -1089
rect 3169 -1157 3227 -1123
rect 3169 -1191 3181 -1157
rect 3215 -1191 3227 -1157
rect 3169 -1225 3227 -1191
rect 3169 -1259 3181 -1225
rect 3215 -1259 3227 -1225
rect 3169 -1274 3227 -1259
rect 3427 -1089 3485 -1074
rect 3427 -1123 3439 -1089
rect 3473 -1123 3485 -1089
rect 3427 -1157 3485 -1123
rect 3427 -1191 3439 -1157
rect 3473 -1191 3485 -1157
rect 3427 -1225 3485 -1191
rect 3427 -1259 3439 -1225
rect 3473 -1259 3485 -1225
rect 3427 -1274 3485 -1259
rect 3621 -1089 3679 -1074
rect 3621 -1123 3633 -1089
rect 3667 -1123 3679 -1089
rect 3621 -1157 3679 -1123
rect 3621 -1191 3633 -1157
rect 3667 -1191 3679 -1157
rect 3621 -1225 3679 -1191
rect 3621 -1259 3633 -1225
rect 3667 -1259 3679 -1225
rect 3621 -1274 3679 -1259
rect 3879 -1089 3937 -1074
rect 3879 -1123 3891 -1089
rect 3925 -1123 3937 -1089
rect 3879 -1157 3937 -1123
rect 3879 -1191 3891 -1157
rect 3925 -1191 3937 -1157
rect 3879 -1225 3937 -1191
rect 3879 -1259 3891 -1225
rect 3925 -1259 3937 -1225
rect 3879 -1274 3937 -1259
rect 4137 -1089 4195 -1074
rect 4137 -1123 4149 -1089
rect 4183 -1123 4195 -1089
rect 4137 -1157 4195 -1123
rect 4137 -1191 4149 -1157
rect 4183 -1191 4195 -1157
rect 4137 -1225 4195 -1191
rect 4137 -1259 4149 -1225
rect 4183 -1259 4195 -1225
rect 4137 -1274 4195 -1259
rect 4395 -1089 4453 -1074
rect 4395 -1123 4407 -1089
rect 4441 -1123 4453 -1089
rect 4395 -1157 4453 -1123
rect 4395 -1191 4407 -1157
rect 4441 -1191 4453 -1157
rect 4395 -1225 4453 -1191
rect 4395 -1259 4407 -1225
rect 4441 -1259 4453 -1225
rect 4395 -1274 4453 -1259
rect 4653 -1089 4711 -1074
rect 4653 -1123 4665 -1089
rect 4699 -1123 4711 -1089
rect 4653 -1157 4711 -1123
rect 4653 -1191 4665 -1157
rect 4699 -1191 4711 -1157
rect 4653 -1225 4711 -1191
rect 4653 -1259 4665 -1225
rect 4699 -1259 4711 -1225
rect 4653 -1274 4711 -1259
rect 4847 -1089 4905 -1074
rect 4847 -1123 4859 -1089
rect 4893 -1123 4905 -1089
rect 4847 -1157 4905 -1123
rect 4847 -1191 4859 -1157
rect 4893 -1191 4905 -1157
rect 4847 -1225 4905 -1191
rect 4847 -1259 4859 -1225
rect 4893 -1259 4905 -1225
rect 4847 -1274 4905 -1259
rect 5105 -1089 5163 -1074
rect 5105 -1123 5117 -1089
rect 5151 -1123 5163 -1089
rect 5105 -1157 5163 -1123
rect 5105 -1191 5117 -1157
rect 5151 -1191 5163 -1157
rect 5105 -1225 5163 -1191
rect 5105 -1259 5117 -1225
rect 5151 -1259 5163 -1225
rect 5105 -1274 5163 -1259
rect 5333 -1089 5391 -1074
rect 5333 -1123 5345 -1089
rect 5379 -1123 5391 -1089
rect 5333 -1157 5391 -1123
rect 5333 -1191 5345 -1157
rect 5379 -1191 5391 -1157
rect 5333 -1225 5391 -1191
rect 5333 -1259 5345 -1225
rect 5379 -1259 5391 -1225
rect 5333 -1274 5391 -1259
rect 5591 -1089 5649 -1074
rect 5591 -1123 5603 -1089
rect 5637 -1123 5649 -1089
rect 5591 -1157 5649 -1123
rect 5591 -1191 5603 -1157
rect 5637 -1191 5649 -1157
rect 5591 -1225 5649 -1191
rect 5591 -1259 5603 -1225
rect 5637 -1259 5649 -1225
rect 5591 -1274 5649 -1259
rect 5784 -1089 5842 -1074
rect 5784 -1123 5796 -1089
rect 5830 -1123 5842 -1089
rect 5784 -1157 5842 -1123
rect 5784 -1191 5796 -1157
rect 5830 -1191 5842 -1157
rect 5784 -1225 5842 -1191
rect 5784 -1259 5796 -1225
rect 5830 -1259 5842 -1225
rect 5784 -1274 5842 -1259
rect 6042 -1089 6100 -1074
rect 6042 -1123 6054 -1089
rect 6088 -1123 6100 -1089
rect 6042 -1157 6100 -1123
rect 6042 -1191 6054 -1157
rect 6088 -1191 6100 -1157
rect 6042 -1225 6100 -1191
rect 6042 -1259 6054 -1225
rect 6088 -1259 6100 -1225
rect 6042 -1274 6100 -1259
rect 6300 -1089 6358 -1074
rect 6300 -1123 6312 -1089
rect 6346 -1123 6358 -1089
rect 6300 -1157 6358 -1123
rect 6300 -1191 6312 -1157
rect 6346 -1191 6358 -1157
rect 6300 -1225 6358 -1191
rect 6300 -1259 6312 -1225
rect 6346 -1259 6358 -1225
rect 6300 -1274 6358 -1259
rect 6558 -1089 6616 -1074
rect 6558 -1123 6570 -1089
rect 6604 -1123 6616 -1089
rect 6558 -1157 6616 -1123
rect 6558 -1191 6570 -1157
rect 6604 -1191 6616 -1157
rect 6558 -1225 6616 -1191
rect 6558 -1259 6570 -1225
rect 6604 -1259 6616 -1225
rect 6558 -1274 6616 -1259
rect 6816 -1089 6874 -1074
rect 6816 -1123 6828 -1089
rect 6862 -1123 6874 -1089
rect 6816 -1157 6874 -1123
rect 6816 -1191 6828 -1157
rect 6862 -1191 6874 -1157
rect 6816 -1225 6874 -1191
rect 6816 -1259 6828 -1225
rect 6862 -1259 6874 -1225
rect 6816 -1274 6874 -1259
rect 7010 -1089 7068 -1074
rect 7010 -1123 7022 -1089
rect 7056 -1123 7068 -1089
rect 7010 -1157 7068 -1123
rect 7010 -1191 7022 -1157
rect 7056 -1191 7068 -1157
rect 7010 -1225 7068 -1191
rect 7010 -1259 7022 -1225
rect 7056 -1259 7068 -1225
rect 7010 -1274 7068 -1259
rect 7268 -1089 7326 -1074
rect 7268 -1123 7280 -1089
rect 7314 -1123 7326 -1089
rect 7268 -1157 7326 -1123
rect 7268 -1191 7280 -1157
rect 7314 -1191 7326 -1157
rect 7268 -1225 7326 -1191
rect 7268 -1259 7280 -1225
rect 7314 -1259 7326 -1225
rect 7268 -1274 7326 -1259
rect 7526 -1089 7584 -1074
rect 7526 -1123 7538 -1089
rect 7572 -1123 7584 -1089
rect 7526 -1157 7584 -1123
rect 7526 -1191 7538 -1157
rect 7572 -1191 7584 -1157
rect 7526 -1225 7584 -1191
rect 7526 -1259 7538 -1225
rect 7572 -1259 7584 -1225
rect 7526 -1274 7584 -1259
rect 7784 -1089 7842 -1074
rect 7784 -1123 7796 -1089
rect 7830 -1123 7842 -1089
rect 7784 -1157 7842 -1123
rect 7784 -1191 7796 -1157
rect 7830 -1191 7842 -1157
rect 7784 -1225 7842 -1191
rect 7784 -1259 7796 -1225
rect 7830 -1259 7842 -1225
rect 7784 -1274 7842 -1259
rect 7978 -1089 8036 -1074
rect 7978 -1123 7990 -1089
rect 8024 -1123 8036 -1089
rect 7978 -1157 8036 -1123
rect 7978 -1191 7990 -1157
rect 8024 -1191 8036 -1157
rect 7978 -1225 8036 -1191
rect 7978 -1259 7990 -1225
rect 8024 -1259 8036 -1225
rect 7978 -1274 8036 -1259
rect 8236 -1089 8294 -1074
rect 8236 -1123 8248 -1089
rect 8282 -1123 8294 -1089
rect 8236 -1157 8294 -1123
rect 8236 -1191 8248 -1157
rect 8282 -1191 8294 -1157
rect 8236 -1225 8294 -1191
rect 8236 -1259 8248 -1225
rect 8282 -1259 8294 -1225
rect 8236 -1274 8294 -1259
rect 8494 -1089 8552 -1074
rect 8494 -1123 8506 -1089
rect 8540 -1123 8552 -1089
rect 8494 -1157 8552 -1123
rect 8494 -1191 8506 -1157
rect 8540 -1191 8552 -1157
rect 8494 -1225 8552 -1191
rect 8494 -1259 8506 -1225
rect 8540 -1259 8552 -1225
rect 8494 -1274 8552 -1259
rect 8752 -1089 8810 -1074
rect 8752 -1123 8764 -1089
rect 8798 -1123 8810 -1089
rect 8752 -1157 8810 -1123
rect 8752 -1191 8764 -1157
rect 8798 -1191 8810 -1157
rect 8752 -1225 8810 -1191
rect 8752 -1259 8764 -1225
rect 8798 -1259 8810 -1225
rect 8752 -1274 8810 -1259
rect 9010 -1089 9068 -1074
rect 9010 -1123 9022 -1089
rect 9056 -1123 9068 -1089
rect 9010 -1157 9068 -1123
rect 9010 -1191 9022 -1157
rect 9056 -1191 9068 -1157
rect 9010 -1225 9068 -1191
rect 9010 -1259 9022 -1225
rect 9056 -1259 9068 -1225
rect 9010 -1274 9068 -1259
rect 9204 -1089 9262 -1074
rect 9204 -1123 9216 -1089
rect 9250 -1123 9262 -1089
rect 9204 -1157 9262 -1123
rect 9204 -1191 9216 -1157
rect 9250 -1191 9262 -1157
rect 9204 -1225 9262 -1191
rect 9204 -1259 9216 -1225
rect 9250 -1259 9262 -1225
rect 9204 -1274 9262 -1259
rect 9462 -1089 9520 -1074
rect 9462 -1123 9474 -1089
rect 9508 -1123 9520 -1089
rect 9462 -1157 9520 -1123
rect 9462 -1191 9474 -1157
rect 9508 -1191 9520 -1157
rect 9462 -1225 9520 -1191
rect 9462 -1259 9474 -1225
rect 9508 -1259 9520 -1225
rect 9462 -1274 9520 -1259
rect 975 -2045 1033 -2030
rect 975 -2079 987 -2045
rect 1021 -2079 1033 -2045
rect 975 -2113 1033 -2079
rect 975 -2147 987 -2113
rect 1021 -2147 1033 -2113
rect 975 -2181 1033 -2147
rect 975 -2215 987 -2181
rect 1021 -2215 1033 -2181
rect 975 -2230 1033 -2215
rect 1233 -2045 1291 -2030
rect 1233 -2079 1245 -2045
rect 1279 -2079 1291 -2045
rect 1233 -2113 1291 -2079
rect 1233 -2147 1245 -2113
rect 1279 -2147 1291 -2113
rect 1233 -2181 1291 -2147
rect 1233 -2215 1245 -2181
rect 1279 -2215 1291 -2181
rect 1233 -2230 1291 -2215
rect 1427 -2045 1485 -2030
rect 1427 -2079 1439 -2045
rect 1473 -2079 1485 -2045
rect 1427 -2113 1485 -2079
rect 1427 -2147 1439 -2113
rect 1473 -2147 1485 -2113
rect 1427 -2181 1485 -2147
rect 1427 -2215 1439 -2181
rect 1473 -2215 1485 -2181
rect 1427 -2230 1485 -2215
rect 1685 -2045 1743 -2030
rect 1685 -2079 1697 -2045
rect 1731 -2079 1743 -2045
rect 1685 -2113 1743 -2079
rect 1685 -2147 1697 -2113
rect 1731 -2147 1743 -2113
rect 1685 -2181 1743 -2147
rect 1685 -2215 1697 -2181
rect 1731 -2215 1743 -2181
rect 1685 -2230 1743 -2215
rect 1943 -2045 2001 -2030
rect 1943 -2079 1955 -2045
rect 1989 -2079 2001 -2045
rect 1943 -2113 2001 -2079
rect 1943 -2147 1955 -2113
rect 1989 -2147 2001 -2113
rect 1943 -2181 2001 -2147
rect 1943 -2215 1955 -2181
rect 1989 -2215 2001 -2181
rect 1943 -2230 2001 -2215
rect 2201 -2045 2259 -2030
rect 2201 -2079 2213 -2045
rect 2247 -2079 2259 -2045
rect 2201 -2113 2259 -2079
rect 2201 -2147 2213 -2113
rect 2247 -2147 2259 -2113
rect 2201 -2181 2259 -2147
rect 2201 -2215 2213 -2181
rect 2247 -2215 2259 -2181
rect 2201 -2230 2259 -2215
rect 2459 -2045 2517 -2030
rect 2459 -2079 2471 -2045
rect 2505 -2079 2517 -2045
rect 2459 -2113 2517 -2079
rect 2459 -2147 2471 -2113
rect 2505 -2147 2517 -2113
rect 2459 -2181 2517 -2147
rect 2459 -2215 2471 -2181
rect 2505 -2215 2517 -2181
rect 2459 -2230 2517 -2215
rect 2653 -2045 2711 -2030
rect 2653 -2079 2665 -2045
rect 2699 -2079 2711 -2045
rect 2653 -2113 2711 -2079
rect 2653 -2147 2665 -2113
rect 2699 -2147 2711 -2113
rect 2653 -2181 2711 -2147
rect 2653 -2215 2665 -2181
rect 2699 -2215 2711 -2181
rect 2653 -2230 2711 -2215
rect 2911 -2045 2969 -2030
rect 2911 -2079 2923 -2045
rect 2957 -2079 2969 -2045
rect 2911 -2113 2969 -2079
rect 2911 -2147 2923 -2113
rect 2957 -2147 2969 -2113
rect 2911 -2181 2969 -2147
rect 2911 -2215 2923 -2181
rect 2957 -2215 2969 -2181
rect 2911 -2230 2969 -2215
rect 3169 -2045 3227 -2030
rect 3169 -2079 3181 -2045
rect 3215 -2079 3227 -2045
rect 3169 -2113 3227 -2079
rect 3169 -2147 3181 -2113
rect 3215 -2147 3227 -2113
rect 3169 -2181 3227 -2147
rect 3169 -2215 3181 -2181
rect 3215 -2215 3227 -2181
rect 3169 -2230 3227 -2215
rect 3427 -2045 3485 -2030
rect 3427 -2079 3439 -2045
rect 3473 -2079 3485 -2045
rect 3427 -2113 3485 -2079
rect 3427 -2147 3439 -2113
rect 3473 -2147 3485 -2113
rect 3427 -2181 3485 -2147
rect 3427 -2215 3439 -2181
rect 3473 -2215 3485 -2181
rect 3427 -2230 3485 -2215
rect 3621 -2045 3679 -2030
rect 3621 -2079 3633 -2045
rect 3667 -2079 3679 -2045
rect 3621 -2113 3679 -2079
rect 3621 -2147 3633 -2113
rect 3667 -2147 3679 -2113
rect 3621 -2181 3679 -2147
rect 3621 -2215 3633 -2181
rect 3667 -2215 3679 -2181
rect 3621 -2230 3679 -2215
rect 3879 -2045 3937 -2030
rect 3879 -2079 3891 -2045
rect 3925 -2079 3937 -2045
rect 3879 -2113 3937 -2079
rect 3879 -2147 3891 -2113
rect 3925 -2147 3937 -2113
rect 3879 -2181 3937 -2147
rect 3879 -2215 3891 -2181
rect 3925 -2215 3937 -2181
rect 3879 -2230 3937 -2215
rect 4137 -2045 4195 -2030
rect 4137 -2079 4149 -2045
rect 4183 -2079 4195 -2045
rect 4137 -2113 4195 -2079
rect 4137 -2147 4149 -2113
rect 4183 -2147 4195 -2113
rect 4137 -2181 4195 -2147
rect 4137 -2215 4149 -2181
rect 4183 -2215 4195 -2181
rect 4137 -2230 4195 -2215
rect 4395 -2045 4453 -2030
rect 4395 -2079 4407 -2045
rect 4441 -2079 4453 -2045
rect 4395 -2113 4453 -2079
rect 4395 -2147 4407 -2113
rect 4441 -2147 4453 -2113
rect 4395 -2181 4453 -2147
rect 4395 -2215 4407 -2181
rect 4441 -2215 4453 -2181
rect 4395 -2230 4453 -2215
rect 4653 -2045 4711 -2030
rect 4653 -2079 4665 -2045
rect 4699 -2079 4711 -2045
rect 4653 -2113 4711 -2079
rect 4653 -2147 4665 -2113
rect 4699 -2147 4711 -2113
rect 4653 -2181 4711 -2147
rect 4653 -2215 4665 -2181
rect 4699 -2215 4711 -2181
rect 4653 -2230 4711 -2215
rect 4847 -2045 4905 -2030
rect 4847 -2079 4859 -2045
rect 4893 -2079 4905 -2045
rect 4847 -2113 4905 -2079
rect 4847 -2147 4859 -2113
rect 4893 -2147 4905 -2113
rect 4847 -2181 4905 -2147
rect 4847 -2215 4859 -2181
rect 4893 -2215 4905 -2181
rect 4847 -2230 4905 -2215
rect 5105 -2045 5163 -2030
rect 5105 -2079 5117 -2045
rect 5151 -2079 5163 -2045
rect 5105 -2113 5163 -2079
rect 5105 -2147 5117 -2113
rect 5151 -2147 5163 -2113
rect 5105 -2181 5163 -2147
rect 5105 -2215 5117 -2181
rect 5151 -2215 5163 -2181
rect 5105 -2230 5163 -2215
rect 5333 -2045 5391 -2030
rect 5333 -2079 5345 -2045
rect 5379 -2079 5391 -2045
rect 5333 -2113 5391 -2079
rect 5333 -2147 5345 -2113
rect 5379 -2147 5391 -2113
rect 5333 -2181 5391 -2147
rect 5333 -2215 5345 -2181
rect 5379 -2215 5391 -2181
rect 5333 -2230 5391 -2215
rect 5591 -2045 5649 -2030
rect 5591 -2079 5603 -2045
rect 5637 -2079 5649 -2045
rect 5591 -2113 5649 -2079
rect 5591 -2147 5603 -2113
rect 5637 -2147 5649 -2113
rect 5591 -2181 5649 -2147
rect 5591 -2215 5603 -2181
rect 5637 -2215 5649 -2181
rect 5591 -2230 5649 -2215
rect 5784 -2045 5842 -2030
rect 5784 -2079 5796 -2045
rect 5830 -2079 5842 -2045
rect 5784 -2113 5842 -2079
rect 5784 -2147 5796 -2113
rect 5830 -2147 5842 -2113
rect 5784 -2181 5842 -2147
rect 5784 -2215 5796 -2181
rect 5830 -2215 5842 -2181
rect 5784 -2230 5842 -2215
rect 6042 -2045 6100 -2030
rect 6042 -2079 6054 -2045
rect 6088 -2079 6100 -2045
rect 6042 -2113 6100 -2079
rect 6042 -2147 6054 -2113
rect 6088 -2147 6100 -2113
rect 6042 -2181 6100 -2147
rect 6042 -2215 6054 -2181
rect 6088 -2215 6100 -2181
rect 6042 -2230 6100 -2215
rect 6300 -2045 6358 -2030
rect 6300 -2079 6312 -2045
rect 6346 -2079 6358 -2045
rect 6300 -2113 6358 -2079
rect 6300 -2147 6312 -2113
rect 6346 -2147 6358 -2113
rect 6300 -2181 6358 -2147
rect 6300 -2215 6312 -2181
rect 6346 -2215 6358 -2181
rect 6300 -2230 6358 -2215
rect 6558 -2045 6616 -2030
rect 6558 -2079 6570 -2045
rect 6604 -2079 6616 -2045
rect 6558 -2113 6616 -2079
rect 6558 -2147 6570 -2113
rect 6604 -2147 6616 -2113
rect 6558 -2181 6616 -2147
rect 6558 -2215 6570 -2181
rect 6604 -2215 6616 -2181
rect 6558 -2230 6616 -2215
rect 6816 -2045 6874 -2030
rect 6816 -2079 6828 -2045
rect 6862 -2079 6874 -2045
rect 6816 -2113 6874 -2079
rect 6816 -2147 6828 -2113
rect 6862 -2147 6874 -2113
rect 6816 -2181 6874 -2147
rect 6816 -2215 6828 -2181
rect 6862 -2215 6874 -2181
rect 6816 -2230 6874 -2215
rect 7010 -2045 7068 -2030
rect 7010 -2079 7022 -2045
rect 7056 -2079 7068 -2045
rect 7010 -2113 7068 -2079
rect 7010 -2147 7022 -2113
rect 7056 -2147 7068 -2113
rect 7010 -2181 7068 -2147
rect 7010 -2215 7022 -2181
rect 7056 -2215 7068 -2181
rect 7010 -2230 7068 -2215
rect 7268 -2045 7326 -2030
rect 7268 -2079 7280 -2045
rect 7314 -2079 7326 -2045
rect 7268 -2113 7326 -2079
rect 7268 -2147 7280 -2113
rect 7314 -2147 7326 -2113
rect 7268 -2181 7326 -2147
rect 7268 -2215 7280 -2181
rect 7314 -2215 7326 -2181
rect 7268 -2230 7326 -2215
rect 7526 -2045 7584 -2030
rect 7526 -2079 7538 -2045
rect 7572 -2079 7584 -2045
rect 7526 -2113 7584 -2079
rect 7526 -2147 7538 -2113
rect 7572 -2147 7584 -2113
rect 7526 -2181 7584 -2147
rect 7526 -2215 7538 -2181
rect 7572 -2215 7584 -2181
rect 7526 -2230 7584 -2215
rect 7784 -2045 7842 -2030
rect 7784 -2079 7796 -2045
rect 7830 -2079 7842 -2045
rect 7784 -2113 7842 -2079
rect 7784 -2147 7796 -2113
rect 7830 -2147 7842 -2113
rect 7784 -2181 7842 -2147
rect 7784 -2215 7796 -2181
rect 7830 -2215 7842 -2181
rect 7784 -2230 7842 -2215
rect 7978 -2045 8036 -2030
rect 7978 -2079 7990 -2045
rect 8024 -2079 8036 -2045
rect 7978 -2113 8036 -2079
rect 7978 -2147 7990 -2113
rect 8024 -2147 8036 -2113
rect 7978 -2181 8036 -2147
rect 7978 -2215 7990 -2181
rect 8024 -2215 8036 -2181
rect 7978 -2230 8036 -2215
rect 8236 -2045 8294 -2030
rect 8236 -2079 8248 -2045
rect 8282 -2079 8294 -2045
rect 8236 -2113 8294 -2079
rect 8236 -2147 8248 -2113
rect 8282 -2147 8294 -2113
rect 8236 -2181 8294 -2147
rect 8236 -2215 8248 -2181
rect 8282 -2215 8294 -2181
rect 8236 -2230 8294 -2215
rect 8494 -2045 8552 -2030
rect 8494 -2079 8506 -2045
rect 8540 -2079 8552 -2045
rect 8494 -2113 8552 -2079
rect 8494 -2147 8506 -2113
rect 8540 -2147 8552 -2113
rect 8494 -2181 8552 -2147
rect 8494 -2215 8506 -2181
rect 8540 -2215 8552 -2181
rect 8494 -2230 8552 -2215
rect 8752 -2045 8810 -2030
rect 8752 -2079 8764 -2045
rect 8798 -2079 8810 -2045
rect 8752 -2113 8810 -2079
rect 8752 -2147 8764 -2113
rect 8798 -2147 8810 -2113
rect 8752 -2181 8810 -2147
rect 8752 -2215 8764 -2181
rect 8798 -2215 8810 -2181
rect 8752 -2230 8810 -2215
rect 9010 -2045 9068 -2030
rect 9010 -2079 9022 -2045
rect 9056 -2079 9068 -2045
rect 9010 -2113 9068 -2079
rect 9010 -2147 9022 -2113
rect 9056 -2147 9068 -2113
rect 9010 -2181 9068 -2147
rect 9010 -2215 9022 -2181
rect 9056 -2215 9068 -2181
rect 9010 -2230 9068 -2215
rect 9204 -2045 9262 -2030
rect 9204 -2079 9216 -2045
rect 9250 -2079 9262 -2045
rect 9204 -2113 9262 -2079
rect 9204 -2147 9216 -2113
rect 9250 -2147 9262 -2113
rect 9204 -2181 9262 -2147
rect 9204 -2215 9216 -2181
rect 9250 -2215 9262 -2181
rect 9204 -2230 9262 -2215
rect 9462 -2045 9520 -2030
rect 9462 -2079 9474 -2045
rect 9508 -2079 9520 -2045
rect 9462 -2113 9520 -2079
rect 9462 -2147 9474 -2113
rect 9508 -2147 9520 -2113
rect 9462 -2181 9520 -2147
rect 9462 -2215 9474 -2181
rect 9508 -2215 9520 -2181
rect 9462 -2230 9520 -2215
rect 975 -2736 1033 -2721
rect 975 -2770 987 -2736
rect 1021 -2770 1033 -2736
rect 975 -2804 1033 -2770
rect 975 -2838 987 -2804
rect 1021 -2838 1033 -2804
rect 975 -2872 1033 -2838
rect 975 -2906 987 -2872
rect 1021 -2906 1033 -2872
rect 975 -2921 1033 -2906
rect 1233 -2736 1291 -2721
rect 1233 -2770 1245 -2736
rect 1279 -2770 1291 -2736
rect 1233 -2804 1291 -2770
rect 1233 -2838 1245 -2804
rect 1279 -2838 1291 -2804
rect 1233 -2872 1291 -2838
rect 1233 -2906 1245 -2872
rect 1279 -2906 1291 -2872
rect 1233 -2921 1291 -2906
rect 1427 -2736 1485 -2721
rect 1427 -2770 1439 -2736
rect 1473 -2770 1485 -2736
rect 1427 -2804 1485 -2770
rect 1427 -2838 1439 -2804
rect 1473 -2838 1485 -2804
rect 1427 -2872 1485 -2838
rect 1427 -2906 1439 -2872
rect 1473 -2906 1485 -2872
rect 1427 -2921 1485 -2906
rect 1685 -2736 1743 -2721
rect 1685 -2770 1697 -2736
rect 1731 -2770 1743 -2736
rect 1685 -2804 1743 -2770
rect 1685 -2838 1697 -2804
rect 1731 -2838 1743 -2804
rect 1685 -2872 1743 -2838
rect 1685 -2906 1697 -2872
rect 1731 -2906 1743 -2872
rect 1685 -2921 1743 -2906
rect 1943 -2736 2001 -2721
rect 1943 -2770 1955 -2736
rect 1989 -2770 2001 -2736
rect 1943 -2804 2001 -2770
rect 1943 -2838 1955 -2804
rect 1989 -2838 2001 -2804
rect 1943 -2872 2001 -2838
rect 1943 -2906 1955 -2872
rect 1989 -2906 2001 -2872
rect 1943 -2921 2001 -2906
rect 2201 -2736 2259 -2721
rect 2201 -2770 2213 -2736
rect 2247 -2770 2259 -2736
rect 2201 -2804 2259 -2770
rect 2201 -2838 2213 -2804
rect 2247 -2838 2259 -2804
rect 2201 -2872 2259 -2838
rect 2201 -2906 2213 -2872
rect 2247 -2906 2259 -2872
rect 2201 -2921 2259 -2906
rect 2459 -2736 2517 -2721
rect 2459 -2770 2471 -2736
rect 2505 -2770 2517 -2736
rect 2459 -2804 2517 -2770
rect 2459 -2838 2471 -2804
rect 2505 -2838 2517 -2804
rect 2459 -2872 2517 -2838
rect 2459 -2906 2471 -2872
rect 2505 -2906 2517 -2872
rect 2459 -2921 2517 -2906
rect 2653 -2736 2711 -2721
rect 2653 -2770 2665 -2736
rect 2699 -2770 2711 -2736
rect 2653 -2804 2711 -2770
rect 2653 -2838 2665 -2804
rect 2699 -2838 2711 -2804
rect 2653 -2872 2711 -2838
rect 2653 -2906 2665 -2872
rect 2699 -2906 2711 -2872
rect 2653 -2921 2711 -2906
rect 2911 -2736 2969 -2721
rect 2911 -2770 2923 -2736
rect 2957 -2770 2969 -2736
rect 2911 -2804 2969 -2770
rect 2911 -2838 2923 -2804
rect 2957 -2838 2969 -2804
rect 2911 -2872 2969 -2838
rect 2911 -2906 2923 -2872
rect 2957 -2906 2969 -2872
rect 2911 -2921 2969 -2906
rect 3169 -2736 3227 -2721
rect 3169 -2770 3181 -2736
rect 3215 -2770 3227 -2736
rect 3169 -2804 3227 -2770
rect 3169 -2838 3181 -2804
rect 3215 -2838 3227 -2804
rect 3169 -2872 3227 -2838
rect 3169 -2906 3181 -2872
rect 3215 -2906 3227 -2872
rect 3169 -2921 3227 -2906
rect 3427 -2736 3485 -2721
rect 3427 -2770 3439 -2736
rect 3473 -2770 3485 -2736
rect 3427 -2804 3485 -2770
rect 3427 -2838 3439 -2804
rect 3473 -2838 3485 -2804
rect 3427 -2872 3485 -2838
rect 3427 -2906 3439 -2872
rect 3473 -2906 3485 -2872
rect 3427 -2921 3485 -2906
rect 3621 -2736 3679 -2721
rect 3621 -2770 3633 -2736
rect 3667 -2770 3679 -2736
rect 3621 -2804 3679 -2770
rect 3621 -2838 3633 -2804
rect 3667 -2838 3679 -2804
rect 3621 -2872 3679 -2838
rect 3621 -2906 3633 -2872
rect 3667 -2906 3679 -2872
rect 3621 -2921 3679 -2906
rect 3879 -2736 3937 -2721
rect 3879 -2770 3891 -2736
rect 3925 -2770 3937 -2736
rect 3879 -2804 3937 -2770
rect 3879 -2838 3891 -2804
rect 3925 -2838 3937 -2804
rect 3879 -2872 3937 -2838
rect 3879 -2906 3891 -2872
rect 3925 -2906 3937 -2872
rect 3879 -2921 3937 -2906
rect 4137 -2736 4195 -2721
rect 4137 -2770 4149 -2736
rect 4183 -2770 4195 -2736
rect 4137 -2804 4195 -2770
rect 4137 -2838 4149 -2804
rect 4183 -2838 4195 -2804
rect 4137 -2872 4195 -2838
rect 4137 -2906 4149 -2872
rect 4183 -2906 4195 -2872
rect 4137 -2921 4195 -2906
rect 4395 -2736 4453 -2721
rect 4395 -2770 4407 -2736
rect 4441 -2770 4453 -2736
rect 4395 -2804 4453 -2770
rect 4395 -2838 4407 -2804
rect 4441 -2838 4453 -2804
rect 4395 -2872 4453 -2838
rect 4395 -2906 4407 -2872
rect 4441 -2906 4453 -2872
rect 4395 -2921 4453 -2906
rect 4653 -2736 4711 -2721
rect 4653 -2770 4665 -2736
rect 4699 -2770 4711 -2736
rect 4653 -2804 4711 -2770
rect 4653 -2838 4665 -2804
rect 4699 -2838 4711 -2804
rect 4653 -2872 4711 -2838
rect 4653 -2906 4665 -2872
rect 4699 -2906 4711 -2872
rect 4653 -2921 4711 -2906
rect 4847 -2736 4905 -2721
rect 4847 -2770 4859 -2736
rect 4893 -2770 4905 -2736
rect 4847 -2804 4905 -2770
rect 4847 -2838 4859 -2804
rect 4893 -2838 4905 -2804
rect 4847 -2872 4905 -2838
rect 4847 -2906 4859 -2872
rect 4893 -2906 4905 -2872
rect 4847 -2921 4905 -2906
rect 5105 -2736 5163 -2721
rect 5105 -2770 5117 -2736
rect 5151 -2770 5163 -2736
rect 5105 -2804 5163 -2770
rect 5105 -2838 5117 -2804
rect 5151 -2838 5163 -2804
rect 5105 -2872 5163 -2838
rect 5105 -2906 5117 -2872
rect 5151 -2906 5163 -2872
rect 5105 -2921 5163 -2906
rect 5333 -2736 5391 -2721
rect 5333 -2770 5345 -2736
rect 5379 -2770 5391 -2736
rect 5333 -2804 5391 -2770
rect 5333 -2838 5345 -2804
rect 5379 -2838 5391 -2804
rect 5333 -2872 5391 -2838
rect 5333 -2906 5345 -2872
rect 5379 -2906 5391 -2872
rect 5333 -2921 5391 -2906
rect 5591 -2736 5649 -2721
rect 5591 -2770 5603 -2736
rect 5637 -2770 5649 -2736
rect 5591 -2804 5649 -2770
rect 5591 -2838 5603 -2804
rect 5637 -2838 5649 -2804
rect 5591 -2872 5649 -2838
rect 5591 -2906 5603 -2872
rect 5637 -2906 5649 -2872
rect 5591 -2921 5649 -2906
rect 5784 -2736 5842 -2721
rect 5784 -2770 5796 -2736
rect 5830 -2770 5842 -2736
rect 5784 -2804 5842 -2770
rect 5784 -2838 5796 -2804
rect 5830 -2838 5842 -2804
rect 5784 -2872 5842 -2838
rect 5784 -2906 5796 -2872
rect 5830 -2906 5842 -2872
rect 5784 -2921 5842 -2906
rect 6042 -2736 6100 -2721
rect 6042 -2770 6054 -2736
rect 6088 -2770 6100 -2736
rect 6042 -2804 6100 -2770
rect 6042 -2838 6054 -2804
rect 6088 -2838 6100 -2804
rect 6042 -2872 6100 -2838
rect 6042 -2906 6054 -2872
rect 6088 -2906 6100 -2872
rect 6042 -2921 6100 -2906
rect 6300 -2736 6358 -2721
rect 6300 -2770 6312 -2736
rect 6346 -2770 6358 -2736
rect 6300 -2804 6358 -2770
rect 6300 -2838 6312 -2804
rect 6346 -2838 6358 -2804
rect 6300 -2872 6358 -2838
rect 6300 -2906 6312 -2872
rect 6346 -2906 6358 -2872
rect 6300 -2921 6358 -2906
rect 6558 -2736 6616 -2721
rect 6558 -2770 6570 -2736
rect 6604 -2770 6616 -2736
rect 6558 -2804 6616 -2770
rect 6558 -2838 6570 -2804
rect 6604 -2838 6616 -2804
rect 6558 -2872 6616 -2838
rect 6558 -2906 6570 -2872
rect 6604 -2906 6616 -2872
rect 6558 -2921 6616 -2906
rect 6816 -2736 6874 -2721
rect 6816 -2770 6828 -2736
rect 6862 -2770 6874 -2736
rect 6816 -2804 6874 -2770
rect 6816 -2838 6828 -2804
rect 6862 -2838 6874 -2804
rect 6816 -2872 6874 -2838
rect 6816 -2906 6828 -2872
rect 6862 -2906 6874 -2872
rect 6816 -2921 6874 -2906
rect 7010 -2736 7068 -2721
rect 7010 -2770 7022 -2736
rect 7056 -2770 7068 -2736
rect 7010 -2804 7068 -2770
rect 7010 -2838 7022 -2804
rect 7056 -2838 7068 -2804
rect 7010 -2872 7068 -2838
rect 7010 -2906 7022 -2872
rect 7056 -2906 7068 -2872
rect 7010 -2921 7068 -2906
rect 7268 -2736 7326 -2721
rect 7268 -2770 7280 -2736
rect 7314 -2770 7326 -2736
rect 7268 -2804 7326 -2770
rect 7268 -2838 7280 -2804
rect 7314 -2838 7326 -2804
rect 7268 -2872 7326 -2838
rect 7268 -2906 7280 -2872
rect 7314 -2906 7326 -2872
rect 7268 -2921 7326 -2906
rect 7526 -2736 7584 -2721
rect 7526 -2770 7538 -2736
rect 7572 -2770 7584 -2736
rect 7526 -2804 7584 -2770
rect 7526 -2838 7538 -2804
rect 7572 -2838 7584 -2804
rect 7526 -2872 7584 -2838
rect 7526 -2906 7538 -2872
rect 7572 -2906 7584 -2872
rect 7526 -2921 7584 -2906
rect 7784 -2736 7842 -2721
rect 7784 -2770 7796 -2736
rect 7830 -2770 7842 -2736
rect 7784 -2804 7842 -2770
rect 7784 -2838 7796 -2804
rect 7830 -2838 7842 -2804
rect 7784 -2872 7842 -2838
rect 7784 -2906 7796 -2872
rect 7830 -2906 7842 -2872
rect 7784 -2921 7842 -2906
rect 7978 -2736 8036 -2721
rect 7978 -2770 7990 -2736
rect 8024 -2770 8036 -2736
rect 7978 -2804 8036 -2770
rect 7978 -2838 7990 -2804
rect 8024 -2838 8036 -2804
rect 7978 -2872 8036 -2838
rect 7978 -2906 7990 -2872
rect 8024 -2906 8036 -2872
rect 7978 -2921 8036 -2906
rect 8236 -2736 8294 -2721
rect 8236 -2770 8248 -2736
rect 8282 -2770 8294 -2736
rect 8236 -2804 8294 -2770
rect 8236 -2838 8248 -2804
rect 8282 -2838 8294 -2804
rect 8236 -2872 8294 -2838
rect 8236 -2906 8248 -2872
rect 8282 -2906 8294 -2872
rect 8236 -2921 8294 -2906
rect 8494 -2736 8552 -2721
rect 8494 -2770 8506 -2736
rect 8540 -2770 8552 -2736
rect 8494 -2804 8552 -2770
rect 8494 -2838 8506 -2804
rect 8540 -2838 8552 -2804
rect 8494 -2872 8552 -2838
rect 8494 -2906 8506 -2872
rect 8540 -2906 8552 -2872
rect 8494 -2921 8552 -2906
rect 8752 -2736 8810 -2721
rect 8752 -2770 8764 -2736
rect 8798 -2770 8810 -2736
rect 8752 -2804 8810 -2770
rect 8752 -2838 8764 -2804
rect 8798 -2838 8810 -2804
rect 8752 -2872 8810 -2838
rect 8752 -2906 8764 -2872
rect 8798 -2906 8810 -2872
rect 8752 -2921 8810 -2906
rect 9010 -2736 9068 -2721
rect 9010 -2770 9022 -2736
rect 9056 -2770 9068 -2736
rect 9010 -2804 9068 -2770
rect 9010 -2838 9022 -2804
rect 9056 -2838 9068 -2804
rect 9010 -2872 9068 -2838
rect 9010 -2906 9022 -2872
rect 9056 -2906 9068 -2872
rect 9010 -2921 9068 -2906
rect 9204 -2736 9262 -2721
rect 9204 -2770 9216 -2736
rect 9250 -2770 9262 -2736
rect 9204 -2804 9262 -2770
rect 9204 -2838 9216 -2804
rect 9250 -2838 9262 -2804
rect 9204 -2872 9262 -2838
rect 9204 -2906 9216 -2872
rect 9250 -2906 9262 -2872
rect 9204 -2921 9262 -2906
rect 9462 -2736 9520 -2721
rect 9462 -2770 9474 -2736
rect 9508 -2770 9520 -2736
rect 9462 -2804 9520 -2770
rect 9462 -2838 9474 -2804
rect 9508 -2838 9520 -2804
rect 9462 -2872 9520 -2838
rect 9462 -2906 9474 -2872
rect 9508 -2906 9520 -2872
rect 9462 -2921 9520 -2906
rect 975 -3726 1033 -3711
rect 975 -3760 987 -3726
rect 1021 -3760 1033 -3726
rect 975 -3794 1033 -3760
rect 975 -3828 987 -3794
rect 1021 -3828 1033 -3794
rect 975 -3862 1033 -3828
rect 975 -3896 987 -3862
rect 1021 -3896 1033 -3862
rect 975 -3911 1033 -3896
rect 1233 -3726 1291 -3711
rect 1233 -3760 1245 -3726
rect 1279 -3760 1291 -3726
rect 1233 -3794 1291 -3760
rect 1233 -3828 1245 -3794
rect 1279 -3828 1291 -3794
rect 1233 -3862 1291 -3828
rect 1233 -3896 1245 -3862
rect 1279 -3896 1291 -3862
rect 1233 -3911 1291 -3896
rect 1427 -3726 1485 -3711
rect 1427 -3760 1439 -3726
rect 1473 -3760 1485 -3726
rect 1427 -3794 1485 -3760
rect 1427 -3828 1439 -3794
rect 1473 -3828 1485 -3794
rect 1427 -3862 1485 -3828
rect 1427 -3896 1439 -3862
rect 1473 -3896 1485 -3862
rect 1427 -3911 1485 -3896
rect 1685 -3726 1743 -3711
rect 1685 -3760 1697 -3726
rect 1731 -3760 1743 -3726
rect 1685 -3794 1743 -3760
rect 1685 -3828 1697 -3794
rect 1731 -3828 1743 -3794
rect 1685 -3862 1743 -3828
rect 1685 -3896 1697 -3862
rect 1731 -3896 1743 -3862
rect 1685 -3911 1743 -3896
rect 1943 -3726 2001 -3711
rect 1943 -3760 1955 -3726
rect 1989 -3760 2001 -3726
rect 1943 -3794 2001 -3760
rect 1943 -3828 1955 -3794
rect 1989 -3828 2001 -3794
rect 1943 -3862 2001 -3828
rect 1943 -3896 1955 -3862
rect 1989 -3896 2001 -3862
rect 1943 -3911 2001 -3896
rect 2201 -3726 2259 -3711
rect 2201 -3760 2213 -3726
rect 2247 -3760 2259 -3726
rect 2201 -3794 2259 -3760
rect 2201 -3828 2213 -3794
rect 2247 -3828 2259 -3794
rect 2201 -3862 2259 -3828
rect 2201 -3896 2213 -3862
rect 2247 -3896 2259 -3862
rect 2201 -3911 2259 -3896
rect 2459 -3726 2517 -3711
rect 2459 -3760 2471 -3726
rect 2505 -3760 2517 -3726
rect 2459 -3794 2517 -3760
rect 2459 -3828 2471 -3794
rect 2505 -3828 2517 -3794
rect 2459 -3862 2517 -3828
rect 2459 -3896 2471 -3862
rect 2505 -3896 2517 -3862
rect 2459 -3911 2517 -3896
rect 2653 -3726 2711 -3711
rect 2653 -3760 2665 -3726
rect 2699 -3760 2711 -3726
rect 2653 -3794 2711 -3760
rect 2653 -3828 2665 -3794
rect 2699 -3828 2711 -3794
rect 2653 -3862 2711 -3828
rect 2653 -3896 2665 -3862
rect 2699 -3896 2711 -3862
rect 2653 -3911 2711 -3896
rect 2911 -3726 2969 -3711
rect 2911 -3760 2923 -3726
rect 2957 -3760 2969 -3726
rect 2911 -3794 2969 -3760
rect 2911 -3828 2923 -3794
rect 2957 -3828 2969 -3794
rect 2911 -3862 2969 -3828
rect 2911 -3896 2923 -3862
rect 2957 -3896 2969 -3862
rect 2911 -3911 2969 -3896
rect 3169 -3726 3227 -3711
rect 3169 -3760 3181 -3726
rect 3215 -3760 3227 -3726
rect 3169 -3794 3227 -3760
rect 3169 -3828 3181 -3794
rect 3215 -3828 3227 -3794
rect 3169 -3862 3227 -3828
rect 3169 -3896 3181 -3862
rect 3215 -3896 3227 -3862
rect 3169 -3911 3227 -3896
rect 3427 -3726 3485 -3711
rect 3427 -3760 3439 -3726
rect 3473 -3760 3485 -3726
rect 3427 -3794 3485 -3760
rect 3427 -3828 3439 -3794
rect 3473 -3828 3485 -3794
rect 3427 -3862 3485 -3828
rect 3427 -3896 3439 -3862
rect 3473 -3896 3485 -3862
rect 3427 -3911 3485 -3896
rect 3621 -3726 3679 -3711
rect 3621 -3760 3633 -3726
rect 3667 -3760 3679 -3726
rect 3621 -3794 3679 -3760
rect 3621 -3828 3633 -3794
rect 3667 -3828 3679 -3794
rect 3621 -3862 3679 -3828
rect 3621 -3896 3633 -3862
rect 3667 -3896 3679 -3862
rect 3621 -3911 3679 -3896
rect 3879 -3726 3937 -3711
rect 3879 -3760 3891 -3726
rect 3925 -3760 3937 -3726
rect 3879 -3794 3937 -3760
rect 3879 -3828 3891 -3794
rect 3925 -3828 3937 -3794
rect 3879 -3862 3937 -3828
rect 3879 -3896 3891 -3862
rect 3925 -3896 3937 -3862
rect 3879 -3911 3937 -3896
rect 4137 -3726 4195 -3711
rect 4137 -3760 4149 -3726
rect 4183 -3760 4195 -3726
rect 4137 -3794 4195 -3760
rect 4137 -3828 4149 -3794
rect 4183 -3828 4195 -3794
rect 4137 -3862 4195 -3828
rect 4137 -3896 4149 -3862
rect 4183 -3896 4195 -3862
rect 4137 -3911 4195 -3896
rect 4395 -3726 4453 -3711
rect 4395 -3760 4407 -3726
rect 4441 -3760 4453 -3726
rect 4395 -3794 4453 -3760
rect 4395 -3828 4407 -3794
rect 4441 -3828 4453 -3794
rect 4395 -3862 4453 -3828
rect 4395 -3896 4407 -3862
rect 4441 -3896 4453 -3862
rect 4395 -3911 4453 -3896
rect 4653 -3726 4711 -3711
rect 4653 -3760 4665 -3726
rect 4699 -3760 4711 -3726
rect 4653 -3794 4711 -3760
rect 4653 -3828 4665 -3794
rect 4699 -3828 4711 -3794
rect 4653 -3862 4711 -3828
rect 4653 -3896 4665 -3862
rect 4699 -3896 4711 -3862
rect 4653 -3911 4711 -3896
rect 4847 -3726 4905 -3711
rect 4847 -3760 4859 -3726
rect 4893 -3760 4905 -3726
rect 4847 -3794 4905 -3760
rect 4847 -3828 4859 -3794
rect 4893 -3828 4905 -3794
rect 4847 -3862 4905 -3828
rect 4847 -3896 4859 -3862
rect 4893 -3896 4905 -3862
rect 4847 -3911 4905 -3896
rect 5105 -3726 5163 -3711
rect 5105 -3760 5117 -3726
rect 5151 -3760 5163 -3726
rect 5105 -3794 5163 -3760
rect 5105 -3828 5117 -3794
rect 5151 -3828 5163 -3794
rect 5105 -3862 5163 -3828
rect 5105 -3896 5117 -3862
rect 5151 -3896 5163 -3862
rect 5105 -3911 5163 -3896
rect 5333 -3726 5391 -3711
rect 5333 -3760 5345 -3726
rect 5379 -3760 5391 -3726
rect 5333 -3794 5391 -3760
rect 5333 -3828 5345 -3794
rect 5379 -3828 5391 -3794
rect 5333 -3862 5391 -3828
rect 5333 -3896 5345 -3862
rect 5379 -3896 5391 -3862
rect 5333 -3911 5391 -3896
rect 5591 -3726 5649 -3711
rect 5591 -3760 5603 -3726
rect 5637 -3760 5649 -3726
rect 5591 -3794 5649 -3760
rect 5591 -3828 5603 -3794
rect 5637 -3828 5649 -3794
rect 5591 -3862 5649 -3828
rect 5591 -3896 5603 -3862
rect 5637 -3896 5649 -3862
rect 5591 -3911 5649 -3896
rect 5784 -3726 5842 -3711
rect 5784 -3760 5796 -3726
rect 5830 -3760 5842 -3726
rect 5784 -3794 5842 -3760
rect 5784 -3828 5796 -3794
rect 5830 -3828 5842 -3794
rect 5784 -3862 5842 -3828
rect 5784 -3896 5796 -3862
rect 5830 -3896 5842 -3862
rect 5784 -3911 5842 -3896
rect 6042 -3726 6100 -3711
rect 6042 -3760 6054 -3726
rect 6088 -3760 6100 -3726
rect 6042 -3794 6100 -3760
rect 6042 -3828 6054 -3794
rect 6088 -3828 6100 -3794
rect 6042 -3862 6100 -3828
rect 6042 -3896 6054 -3862
rect 6088 -3896 6100 -3862
rect 6042 -3911 6100 -3896
rect 6300 -3726 6358 -3711
rect 6300 -3760 6312 -3726
rect 6346 -3760 6358 -3726
rect 6300 -3794 6358 -3760
rect 6300 -3828 6312 -3794
rect 6346 -3828 6358 -3794
rect 6300 -3862 6358 -3828
rect 6300 -3896 6312 -3862
rect 6346 -3896 6358 -3862
rect 6300 -3911 6358 -3896
rect 6558 -3726 6616 -3711
rect 6558 -3760 6570 -3726
rect 6604 -3760 6616 -3726
rect 6558 -3794 6616 -3760
rect 6558 -3828 6570 -3794
rect 6604 -3828 6616 -3794
rect 6558 -3862 6616 -3828
rect 6558 -3896 6570 -3862
rect 6604 -3896 6616 -3862
rect 6558 -3911 6616 -3896
rect 6816 -3726 6874 -3711
rect 6816 -3760 6828 -3726
rect 6862 -3760 6874 -3726
rect 6816 -3794 6874 -3760
rect 6816 -3828 6828 -3794
rect 6862 -3828 6874 -3794
rect 6816 -3862 6874 -3828
rect 6816 -3896 6828 -3862
rect 6862 -3896 6874 -3862
rect 6816 -3911 6874 -3896
rect 7010 -3726 7068 -3711
rect 7010 -3760 7022 -3726
rect 7056 -3760 7068 -3726
rect 7010 -3794 7068 -3760
rect 7010 -3828 7022 -3794
rect 7056 -3828 7068 -3794
rect 7010 -3862 7068 -3828
rect 7010 -3896 7022 -3862
rect 7056 -3896 7068 -3862
rect 7010 -3911 7068 -3896
rect 7268 -3726 7326 -3711
rect 7268 -3760 7280 -3726
rect 7314 -3760 7326 -3726
rect 7268 -3794 7326 -3760
rect 7268 -3828 7280 -3794
rect 7314 -3828 7326 -3794
rect 7268 -3862 7326 -3828
rect 7268 -3896 7280 -3862
rect 7314 -3896 7326 -3862
rect 7268 -3911 7326 -3896
rect 7526 -3726 7584 -3711
rect 7526 -3760 7538 -3726
rect 7572 -3760 7584 -3726
rect 7526 -3794 7584 -3760
rect 7526 -3828 7538 -3794
rect 7572 -3828 7584 -3794
rect 7526 -3862 7584 -3828
rect 7526 -3896 7538 -3862
rect 7572 -3896 7584 -3862
rect 7526 -3911 7584 -3896
rect 7784 -3726 7842 -3711
rect 7784 -3760 7796 -3726
rect 7830 -3760 7842 -3726
rect 7784 -3794 7842 -3760
rect 7784 -3828 7796 -3794
rect 7830 -3828 7842 -3794
rect 7784 -3862 7842 -3828
rect 7784 -3896 7796 -3862
rect 7830 -3896 7842 -3862
rect 7784 -3911 7842 -3896
rect 7978 -3726 8036 -3711
rect 7978 -3760 7990 -3726
rect 8024 -3760 8036 -3726
rect 7978 -3794 8036 -3760
rect 7978 -3828 7990 -3794
rect 8024 -3828 8036 -3794
rect 7978 -3862 8036 -3828
rect 7978 -3896 7990 -3862
rect 8024 -3896 8036 -3862
rect 7978 -3911 8036 -3896
rect 8236 -3726 8294 -3711
rect 8236 -3760 8248 -3726
rect 8282 -3760 8294 -3726
rect 8236 -3794 8294 -3760
rect 8236 -3828 8248 -3794
rect 8282 -3828 8294 -3794
rect 8236 -3862 8294 -3828
rect 8236 -3896 8248 -3862
rect 8282 -3896 8294 -3862
rect 8236 -3911 8294 -3896
rect 8494 -3726 8552 -3711
rect 8494 -3760 8506 -3726
rect 8540 -3760 8552 -3726
rect 8494 -3794 8552 -3760
rect 8494 -3828 8506 -3794
rect 8540 -3828 8552 -3794
rect 8494 -3862 8552 -3828
rect 8494 -3896 8506 -3862
rect 8540 -3896 8552 -3862
rect 8494 -3911 8552 -3896
rect 8752 -3726 8810 -3711
rect 8752 -3760 8764 -3726
rect 8798 -3760 8810 -3726
rect 8752 -3794 8810 -3760
rect 8752 -3828 8764 -3794
rect 8798 -3828 8810 -3794
rect 8752 -3862 8810 -3828
rect 8752 -3896 8764 -3862
rect 8798 -3896 8810 -3862
rect 8752 -3911 8810 -3896
rect 9010 -3726 9068 -3711
rect 9010 -3760 9022 -3726
rect 9056 -3760 9068 -3726
rect 9010 -3794 9068 -3760
rect 9010 -3828 9022 -3794
rect 9056 -3828 9068 -3794
rect 9010 -3862 9068 -3828
rect 9010 -3896 9022 -3862
rect 9056 -3896 9068 -3862
rect 9010 -3911 9068 -3896
rect 9204 -3726 9262 -3711
rect 9204 -3760 9216 -3726
rect 9250 -3760 9262 -3726
rect 9204 -3794 9262 -3760
rect 9204 -3828 9216 -3794
rect 9250 -3828 9262 -3794
rect 9204 -3862 9262 -3828
rect 9204 -3896 9216 -3862
rect 9250 -3896 9262 -3862
rect 9204 -3911 9262 -3896
rect 9462 -3726 9520 -3711
rect 9462 -3760 9474 -3726
rect 9508 -3760 9520 -3726
rect 9462 -3794 9520 -3760
rect 9462 -3828 9474 -3794
rect 9508 -3828 9520 -3794
rect 9462 -3862 9520 -3828
rect 9462 -3896 9474 -3862
rect 9508 -3896 9520 -3862
rect 9462 -3911 9520 -3896
rect 975 -4282 1033 -4267
rect 975 -4316 987 -4282
rect 1021 -4316 1033 -4282
rect 975 -4350 1033 -4316
rect 975 -4384 987 -4350
rect 1021 -4384 1033 -4350
rect 975 -4418 1033 -4384
rect 975 -4452 987 -4418
rect 1021 -4452 1033 -4418
rect 975 -4467 1033 -4452
rect 1233 -4282 1291 -4267
rect 1233 -4316 1245 -4282
rect 1279 -4316 1291 -4282
rect 1233 -4350 1291 -4316
rect 1233 -4384 1245 -4350
rect 1279 -4384 1291 -4350
rect 1233 -4418 1291 -4384
rect 1233 -4452 1245 -4418
rect 1279 -4452 1291 -4418
rect 1233 -4467 1291 -4452
rect 1427 -4282 1485 -4267
rect 1427 -4316 1439 -4282
rect 1473 -4316 1485 -4282
rect 1427 -4350 1485 -4316
rect 1427 -4384 1439 -4350
rect 1473 -4384 1485 -4350
rect 1427 -4418 1485 -4384
rect 1427 -4452 1439 -4418
rect 1473 -4452 1485 -4418
rect 1427 -4467 1485 -4452
rect 1685 -4282 1743 -4267
rect 1685 -4316 1697 -4282
rect 1731 -4316 1743 -4282
rect 1685 -4350 1743 -4316
rect 1685 -4384 1697 -4350
rect 1731 -4384 1743 -4350
rect 1685 -4418 1743 -4384
rect 1685 -4452 1697 -4418
rect 1731 -4452 1743 -4418
rect 1685 -4467 1743 -4452
rect 1943 -4282 2001 -4267
rect 1943 -4316 1955 -4282
rect 1989 -4316 2001 -4282
rect 1943 -4350 2001 -4316
rect 1943 -4384 1955 -4350
rect 1989 -4384 2001 -4350
rect 1943 -4418 2001 -4384
rect 1943 -4452 1955 -4418
rect 1989 -4452 2001 -4418
rect 1943 -4467 2001 -4452
rect 2201 -4282 2259 -4267
rect 2201 -4316 2213 -4282
rect 2247 -4316 2259 -4282
rect 2201 -4350 2259 -4316
rect 2201 -4384 2213 -4350
rect 2247 -4384 2259 -4350
rect 2201 -4418 2259 -4384
rect 2201 -4452 2213 -4418
rect 2247 -4452 2259 -4418
rect 2201 -4467 2259 -4452
rect 2459 -4282 2517 -4267
rect 2459 -4316 2471 -4282
rect 2505 -4316 2517 -4282
rect 2459 -4350 2517 -4316
rect 2459 -4384 2471 -4350
rect 2505 -4384 2517 -4350
rect 2459 -4418 2517 -4384
rect 2459 -4452 2471 -4418
rect 2505 -4452 2517 -4418
rect 2459 -4467 2517 -4452
rect 2653 -4282 2711 -4267
rect 2653 -4316 2665 -4282
rect 2699 -4316 2711 -4282
rect 2653 -4350 2711 -4316
rect 2653 -4384 2665 -4350
rect 2699 -4384 2711 -4350
rect 2653 -4418 2711 -4384
rect 2653 -4452 2665 -4418
rect 2699 -4452 2711 -4418
rect 2653 -4467 2711 -4452
rect 2911 -4282 2969 -4267
rect 2911 -4316 2923 -4282
rect 2957 -4316 2969 -4282
rect 2911 -4350 2969 -4316
rect 2911 -4384 2923 -4350
rect 2957 -4384 2969 -4350
rect 2911 -4418 2969 -4384
rect 2911 -4452 2923 -4418
rect 2957 -4452 2969 -4418
rect 2911 -4467 2969 -4452
rect 3169 -4282 3227 -4267
rect 3169 -4316 3181 -4282
rect 3215 -4316 3227 -4282
rect 3169 -4350 3227 -4316
rect 3169 -4384 3181 -4350
rect 3215 -4384 3227 -4350
rect 3169 -4418 3227 -4384
rect 3169 -4452 3181 -4418
rect 3215 -4452 3227 -4418
rect 3169 -4467 3227 -4452
rect 3427 -4282 3485 -4267
rect 3427 -4316 3439 -4282
rect 3473 -4316 3485 -4282
rect 3427 -4350 3485 -4316
rect 3427 -4384 3439 -4350
rect 3473 -4384 3485 -4350
rect 3427 -4418 3485 -4384
rect 3427 -4452 3439 -4418
rect 3473 -4452 3485 -4418
rect 3427 -4467 3485 -4452
rect 3621 -4282 3679 -4267
rect 3621 -4316 3633 -4282
rect 3667 -4316 3679 -4282
rect 3621 -4350 3679 -4316
rect 3621 -4384 3633 -4350
rect 3667 -4384 3679 -4350
rect 3621 -4418 3679 -4384
rect 3621 -4452 3633 -4418
rect 3667 -4452 3679 -4418
rect 3621 -4467 3679 -4452
rect 3879 -4282 3937 -4267
rect 3879 -4316 3891 -4282
rect 3925 -4316 3937 -4282
rect 3879 -4350 3937 -4316
rect 3879 -4384 3891 -4350
rect 3925 -4384 3937 -4350
rect 3879 -4418 3937 -4384
rect 3879 -4452 3891 -4418
rect 3925 -4452 3937 -4418
rect 3879 -4467 3937 -4452
rect 4137 -4282 4195 -4267
rect 4137 -4316 4149 -4282
rect 4183 -4316 4195 -4282
rect 4137 -4350 4195 -4316
rect 4137 -4384 4149 -4350
rect 4183 -4384 4195 -4350
rect 4137 -4418 4195 -4384
rect 4137 -4452 4149 -4418
rect 4183 -4452 4195 -4418
rect 4137 -4467 4195 -4452
rect 4395 -4282 4453 -4267
rect 4395 -4316 4407 -4282
rect 4441 -4316 4453 -4282
rect 4395 -4350 4453 -4316
rect 4395 -4384 4407 -4350
rect 4441 -4384 4453 -4350
rect 4395 -4418 4453 -4384
rect 4395 -4452 4407 -4418
rect 4441 -4452 4453 -4418
rect 4395 -4467 4453 -4452
rect 4653 -4282 4711 -4267
rect 4653 -4316 4665 -4282
rect 4699 -4316 4711 -4282
rect 4653 -4350 4711 -4316
rect 4653 -4384 4665 -4350
rect 4699 -4384 4711 -4350
rect 4653 -4418 4711 -4384
rect 4653 -4452 4665 -4418
rect 4699 -4452 4711 -4418
rect 4653 -4467 4711 -4452
rect 4847 -4282 4905 -4267
rect 4847 -4316 4859 -4282
rect 4893 -4316 4905 -4282
rect 4847 -4350 4905 -4316
rect 4847 -4384 4859 -4350
rect 4893 -4384 4905 -4350
rect 4847 -4418 4905 -4384
rect 4847 -4452 4859 -4418
rect 4893 -4452 4905 -4418
rect 4847 -4467 4905 -4452
rect 5105 -4282 5163 -4267
rect 5105 -4316 5117 -4282
rect 5151 -4316 5163 -4282
rect 5105 -4350 5163 -4316
rect 5105 -4384 5117 -4350
rect 5151 -4384 5163 -4350
rect 5105 -4418 5163 -4384
rect 5105 -4452 5117 -4418
rect 5151 -4452 5163 -4418
rect 5105 -4467 5163 -4452
rect 5333 -4282 5391 -4267
rect 5333 -4316 5345 -4282
rect 5379 -4316 5391 -4282
rect 5333 -4350 5391 -4316
rect 5333 -4384 5345 -4350
rect 5379 -4384 5391 -4350
rect 5333 -4418 5391 -4384
rect 5333 -4452 5345 -4418
rect 5379 -4452 5391 -4418
rect 5333 -4467 5391 -4452
rect 5591 -4282 5649 -4267
rect 5591 -4316 5603 -4282
rect 5637 -4316 5649 -4282
rect 5591 -4350 5649 -4316
rect 5591 -4384 5603 -4350
rect 5637 -4384 5649 -4350
rect 5591 -4418 5649 -4384
rect 5591 -4452 5603 -4418
rect 5637 -4452 5649 -4418
rect 5591 -4467 5649 -4452
rect 5784 -4282 5842 -4267
rect 5784 -4316 5796 -4282
rect 5830 -4316 5842 -4282
rect 5784 -4350 5842 -4316
rect 5784 -4384 5796 -4350
rect 5830 -4384 5842 -4350
rect 5784 -4418 5842 -4384
rect 5784 -4452 5796 -4418
rect 5830 -4452 5842 -4418
rect 5784 -4467 5842 -4452
rect 6042 -4282 6100 -4267
rect 6042 -4316 6054 -4282
rect 6088 -4316 6100 -4282
rect 6042 -4350 6100 -4316
rect 6042 -4384 6054 -4350
rect 6088 -4384 6100 -4350
rect 6042 -4418 6100 -4384
rect 6042 -4452 6054 -4418
rect 6088 -4452 6100 -4418
rect 6042 -4467 6100 -4452
rect 6300 -4282 6358 -4267
rect 6300 -4316 6312 -4282
rect 6346 -4316 6358 -4282
rect 6300 -4350 6358 -4316
rect 6300 -4384 6312 -4350
rect 6346 -4384 6358 -4350
rect 6300 -4418 6358 -4384
rect 6300 -4452 6312 -4418
rect 6346 -4452 6358 -4418
rect 6300 -4467 6358 -4452
rect 6558 -4282 6616 -4267
rect 6558 -4316 6570 -4282
rect 6604 -4316 6616 -4282
rect 6558 -4350 6616 -4316
rect 6558 -4384 6570 -4350
rect 6604 -4384 6616 -4350
rect 6558 -4418 6616 -4384
rect 6558 -4452 6570 -4418
rect 6604 -4452 6616 -4418
rect 6558 -4467 6616 -4452
rect 6816 -4282 6874 -4267
rect 6816 -4316 6828 -4282
rect 6862 -4316 6874 -4282
rect 6816 -4350 6874 -4316
rect 6816 -4384 6828 -4350
rect 6862 -4384 6874 -4350
rect 6816 -4418 6874 -4384
rect 6816 -4452 6828 -4418
rect 6862 -4452 6874 -4418
rect 6816 -4467 6874 -4452
rect 7010 -4282 7068 -4267
rect 7010 -4316 7022 -4282
rect 7056 -4316 7068 -4282
rect 7010 -4350 7068 -4316
rect 7010 -4384 7022 -4350
rect 7056 -4384 7068 -4350
rect 7010 -4418 7068 -4384
rect 7010 -4452 7022 -4418
rect 7056 -4452 7068 -4418
rect 7010 -4467 7068 -4452
rect 7268 -4282 7326 -4267
rect 7268 -4316 7280 -4282
rect 7314 -4316 7326 -4282
rect 7268 -4350 7326 -4316
rect 7268 -4384 7280 -4350
rect 7314 -4384 7326 -4350
rect 7268 -4418 7326 -4384
rect 7268 -4452 7280 -4418
rect 7314 -4452 7326 -4418
rect 7268 -4467 7326 -4452
rect 7526 -4282 7584 -4267
rect 7526 -4316 7538 -4282
rect 7572 -4316 7584 -4282
rect 7526 -4350 7584 -4316
rect 7526 -4384 7538 -4350
rect 7572 -4384 7584 -4350
rect 7526 -4418 7584 -4384
rect 7526 -4452 7538 -4418
rect 7572 -4452 7584 -4418
rect 7526 -4467 7584 -4452
rect 7784 -4282 7842 -4267
rect 7784 -4316 7796 -4282
rect 7830 -4316 7842 -4282
rect 7784 -4350 7842 -4316
rect 7784 -4384 7796 -4350
rect 7830 -4384 7842 -4350
rect 7784 -4418 7842 -4384
rect 7784 -4452 7796 -4418
rect 7830 -4452 7842 -4418
rect 7784 -4467 7842 -4452
rect 7978 -4282 8036 -4267
rect 7978 -4316 7990 -4282
rect 8024 -4316 8036 -4282
rect 7978 -4350 8036 -4316
rect 7978 -4384 7990 -4350
rect 8024 -4384 8036 -4350
rect 7978 -4418 8036 -4384
rect 7978 -4452 7990 -4418
rect 8024 -4452 8036 -4418
rect 7978 -4467 8036 -4452
rect 8236 -4282 8294 -4267
rect 8236 -4316 8248 -4282
rect 8282 -4316 8294 -4282
rect 8236 -4350 8294 -4316
rect 8236 -4384 8248 -4350
rect 8282 -4384 8294 -4350
rect 8236 -4418 8294 -4384
rect 8236 -4452 8248 -4418
rect 8282 -4452 8294 -4418
rect 8236 -4467 8294 -4452
rect 8494 -4282 8552 -4267
rect 8494 -4316 8506 -4282
rect 8540 -4316 8552 -4282
rect 8494 -4350 8552 -4316
rect 8494 -4384 8506 -4350
rect 8540 -4384 8552 -4350
rect 8494 -4418 8552 -4384
rect 8494 -4452 8506 -4418
rect 8540 -4452 8552 -4418
rect 8494 -4467 8552 -4452
rect 8752 -4282 8810 -4267
rect 8752 -4316 8764 -4282
rect 8798 -4316 8810 -4282
rect 8752 -4350 8810 -4316
rect 8752 -4384 8764 -4350
rect 8798 -4384 8810 -4350
rect 8752 -4418 8810 -4384
rect 8752 -4452 8764 -4418
rect 8798 -4452 8810 -4418
rect 8752 -4467 8810 -4452
rect 9010 -4282 9068 -4267
rect 9010 -4316 9022 -4282
rect 9056 -4316 9068 -4282
rect 9010 -4350 9068 -4316
rect 9010 -4384 9022 -4350
rect 9056 -4384 9068 -4350
rect 9010 -4418 9068 -4384
rect 9010 -4452 9022 -4418
rect 9056 -4452 9068 -4418
rect 9010 -4467 9068 -4452
rect 9204 -4282 9262 -4267
rect 9204 -4316 9216 -4282
rect 9250 -4316 9262 -4282
rect 9204 -4350 9262 -4316
rect 9204 -4384 9216 -4350
rect 9250 -4384 9262 -4350
rect 9204 -4418 9262 -4384
rect 9204 -4452 9216 -4418
rect 9250 -4452 9262 -4418
rect 9204 -4467 9262 -4452
rect 9462 -4282 9520 -4267
rect 9462 -4316 9474 -4282
rect 9508 -4316 9520 -4282
rect 9462 -4350 9520 -4316
rect 9462 -4384 9474 -4350
rect 9508 -4384 9520 -4350
rect 9462 -4418 9520 -4384
rect 9462 -4452 9474 -4418
rect 9508 -4452 9520 -4418
rect 9462 -4467 9520 -4452
rect 975 -5272 1033 -5257
rect 975 -5306 987 -5272
rect 1021 -5306 1033 -5272
rect 975 -5340 1033 -5306
rect 975 -5374 987 -5340
rect 1021 -5374 1033 -5340
rect 975 -5408 1033 -5374
rect 975 -5442 987 -5408
rect 1021 -5442 1033 -5408
rect 975 -5457 1033 -5442
rect 1233 -5272 1291 -5257
rect 1233 -5306 1245 -5272
rect 1279 -5306 1291 -5272
rect 1233 -5340 1291 -5306
rect 1233 -5374 1245 -5340
rect 1279 -5374 1291 -5340
rect 1233 -5408 1291 -5374
rect 1233 -5442 1245 -5408
rect 1279 -5442 1291 -5408
rect 1233 -5457 1291 -5442
rect 1427 -5272 1485 -5257
rect 1427 -5306 1439 -5272
rect 1473 -5306 1485 -5272
rect 1427 -5340 1485 -5306
rect 1427 -5374 1439 -5340
rect 1473 -5374 1485 -5340
rect 1427 -5408 1485 -5374
rect 1427 -5442 1439 -5408
rect 1473 -5442 1485 -5408
rect 1427 -5457 1485 -5442
rect 1685 -5272 1743 -5257
rect 1685 -5306 1697 -5272
rect 1731 -5306 1743 -5272
rect 1685 -5340 1743 -5306
rect 1685 -5374 1697 -5340
rect 1731 -5374 1743 -5340
rect 1685 -5408 1743 -5374
rect 1685 -5442 1697 -5408
rect 1731 -5442 1743 -5408
rect 1685 -5457 1743 -5442
rect 1943 -5272 2001 -5257
rect 1943 -5306 1955 -5272
rect 1989 -5306 2001 -5272
rect 1943 -5340 2001 -5306
rect 1943 -5374 1955 -5340
rect 1989 -5374 2001 -5340
rect 1943 -5408 2001 -5374
rect 1943 -5442 1955 -5408
rect 1989 -5442 2001 -5408
rect 1943 -5457 2001 -5442
rect 2201 -5272 2259 -5257
rect 2201 -5306 2213 -5272
rect 2247 -5306 2259 -5272
rect 2201 -5340 2259 -5306
rect 2201 -5374 2213 -5340
rect 2247 -5374 2259 -5340
rect 2201 -5408 2259 -5374
rect 2201 -5442 2213 -5408
rect 2247 -5442 2259 -5408
rect 2201 -5457 2259 -5442
rect 2459 -5272 2517 -5257
rect 2459 -5306 2471 -5272
rect 2505 -5306 2517 -5272
rect 2459 -5340 2517 -5306
rect 2459 -5374 2471 -5340
rect 2505 -5374 2517 -5340
rect 2459 -5408 2517 -5374
rect 2459 -5442 2471 -5408
rect 2505 -5442 2517 -5408
rect 2459 -5457 2517 -5442
rect 2653 -5272 2711 -5257
rect 2653 -5306 2665 -5272
rect 2699 -5306 2711 -5272
rect 2653 -5340 2711 -5306
rect 2653 -5374 2665 -5340
rect 2699 -5374 2711 -5340
rect 2653 -5408 2711 -5374
rect 2653 -5442 2665 -5408
rect 2699 -5442 2711 -5408
rect 2653 -5457 2711 -5442
rect 2911 -5272 2969 -5257
rect 2911 -5306 2923 -5272
rect 2957 -5306 2969 -5272
rect 2911 -5340 2969 -5306
rect 2911 -5374 2923 -5340
rect 2957 -5374 2969 -5340
rect 2911 -5408 2969 -5374
rect 2911 -5442 2923 -5408
rect 2957 -5442 2969 -5408
rect 2911 -5457 2969 -5442
rect 3169 -5272 3227 -5257
rect 3169 -5306 3181 -5272
rect 3215 -5306 3227 -5272
rect 3169 -5340 3227 -5306
rect 3169 -5374 3181 -5340
rect 3215 -5374 3227 -5340
rect 3169 -5408 3227 -5374
rect 3169 -5442 3181 -5408
rect 3215 -5442 3227 -5408
rect 3169 -5457 3227 -5442
rect 3427 -5272 3485 -5257
rect 3427 -5306 3439 -5272
rect 3473 -5306 3485 -5272
rect 3427 -5340 3485 -5306
rect 3427 -5374 3439 -5340
rect 3473 -5374 3485 -5340
rect 3427 -5408 3485 -5374
rect 3427 -5442 3439 -5408
rect 3473 -5442 3485 -5408
rect 3427 -5457 3485 -5442
rect 3621 -5272 3679 -5257
rect 3621 -5306 3633 -5272
rect 3667 -5306 3679 -5272
rect 3621 -5340 3679 -5306
rect 3621 -5374 3633 -5340
rect 3667 -5374 3679 -5340
rect 3621 -5408 3679 -5374
rect 3621 -5442 3633 -5408
rect 3667 -5442 3679 -5408
rect 3621 -5457 3679 -5442
rect 3879 -5272 3937 -5257
rect 3879 -5306 3891 -5272
rect 3925 -5306 3937 -5272
rect 3879 -5340 3937 -5306
rect 3879 -5374 3891 -5340
rect 3925 -5374 3937 -5340
rect 3879 -5408 3937 -5374
rect 3879 -5442 3891 -5408
rect 3925 -5442 3937 -5408
rect 3879 -5457 3937 -5442
rect 4137 -5272 4195 -5257
rect 4137 -5306 4149 -5272
rect 4183 -5306 4195 -5272
rect 4137 -5340 4195 -5306
rect 4137 -5374 4149 -5340
rect 4183 -5374 4195 -5340
rect 4137 -5408 4195 -5374
rect 4137 -5442 4149 -5408
rect 4183 -5442 4195 -5408
rect 4137 -5457 4195 -5442
rect 4395 -5272 4453 -5257
rect 4395 -5306 4407 -5272
rect 4441 -5306 4453 -5272
rect 4395 -5340 4453 -5306
rect 4395 -5374 4407 -5340
rect 4441 -5374 4453 -5340
rect 4395 -5408 4453 -5374
rect 4395 -5442 4407 -5408
rect 4441 -5442 4453 -5408
rect 4395 -5457 4453 -5442
rect 4653 -5272 4711 -5257
rect 4653 -5306 4665 -5272
rect 4699 -5306 4711 -5272
rect 4653 -5340 4711 -5306
rect 4653 -5374 4665 -5340
rect 4699 -5374 4711 -5340
rect 4653 -5408 4711 -5374
rect 4653 -5442 4665 -5408
rect 4699 -5442 4711 -5408
rect 4653 -5457 4711 -5442
rect 4847 -5272 4905 -5257
rect 4847 -5306 4859 -5272
rect 4893 -5306 4905 -5272
rect 4847 -5340 4905 -5306
rect 4847 -5374 4859 -5340
rect 4893 -5374 4905 -5340
rect 4847 -5408 4905 -5374
rect 4847 -5442 4859 -5408
rect 4893 -5442 4905 -5408
rect 4847 -5457 4905 -5442
rect 5105 -5272 5163 -5257
rect 5105 -5306 5117 -5272
rect 5151 -5306 5163 -5272
rect 5105 -5340 5163 -5306
rect 5105 -5374 5117 -5340
rect 5151 -5374 5163 -5340
rect 5105 -5408 5163 -5374
rect 5105 -5442 5117 -5408
rect 5151 -5442 5163 -5408
rect 5105 -5457 5163 -5442
rect 5333 -5272 5391 -5257
rect 5333 -5306 5345 -5272
rect 5379 -5306 5391 -5272
rect 5333 -5340 5391 -5306
rect 5333 -5374 5345 -5340
rect 5379 -5374 5391 -5340
rect 5333 -5408 5391 -5374
rect 5333 -5442 5345 -5408
rect 5379 -5442 5391 -5408
rect 5333 -5457 5391 -5442
rect 5591 -5272 5649 -5257
rect 5591 -5306 5603 -5272
rect 5637 -5306 5649 -5272
rect 5591 -5340 5649 -5306
rect 5591 -5374 5603 -5340
rect 5637 -5374 5649 -5340
rect 5591 -5408 5649 -5374
rect 5591 -5442 5603 -5408
rect 5637 -5442 5649 -5408
rect 5591 -5457 5649 -5442
rect 5784 -5272 5842 -5257
rect 5784 -5306 5796 -5272
rect 5830 -5306 5842 -5272
rect 5784 -5340 5842 -5306
rect 5784 -5374 5796 -5340
rect 5830 -5374 5842 -5340
rect 5784 -5408 5842 -5374
rect 5784 -5442 5796 -5408
rect 5830 -5442 5842 -5408
rect 5784 -5457 5842 -5442
rect 6042 -5272 6100 -5257
rect 6042 -5306 6054 -5272
rect 6088 -5306 6100 -5272
rect 6042 -5340 6100 -5306
rect 6042 -5374 6054 -5340
rect 6088 -5374 6100 -5340
rect 6042 -5408 6100 -5374
rect 6042 -5442 6054 -5408
rect 6088 -5442 6100 -5408
rect 6042 -5457 6100 -5442
rect 6300 -5272 6358 -5257
rect 6300 -5306 6312 -5272
rect 6346 -5306 6358 -5272
rect 6300 -5340 6358 -5306
rect 6300 -5374 6312 -5340
rect 6346 -5374 6358 -5340
rect 6300 -5408 6358 -5374
rect 6300 -5442 6312 -5408
rect 6346 -5442 6358 -5408
rect 6300 -5457 6358 -5442
rect 6558 -5272 6616 -5257
rect 6558 -5306 6570 -5272
rect 6604 -5306 6616 -5272
rect 6558 -5340 6616 -5306
rect 6558 -5374 6570 -5340
rect 6604 -5374 6616 -5340
rect 6558 -5408 6616 -5374
rect 6558 -5442 6570 -5408
rect 6604 -5442 6616 -5408
rect 6558 -5457 6616 -5442
rect 6816 -5272 6874 -5257
rect 6816 -5306 6828 -5272
rect 6862 -5306 6874 -5272
rect 6816 -5340 6874 -5306
rect 6816 -5374 6828 -5340
rect 6862 -5374 6874 -5340
rect 6816 -5408 6874 -5374
rect 6816 -5442 6828 -5408
rect 6862 -5442 6874 -5408
rect 6816 -5457 6874 -5442
rect 7010 -5272 7068 -5257
rect 7010 -5306 7022 -5272
rect 7056 -5306 7068 -5272
rect 7010 -5340 7068 -5306
rect 7010 -5374 7022 -5340
rect 7056 -5374 7068 -5340
rect 7010 -5408 7068 -5374
rect 7010 -5442 7022 -5408
rect 7056 -5442 7068 -5408
rect 7010 -5457 7068 -5442
rect 7268 -5272 7326 -5257
rect 7268 -5306 7280 -5272
rect 7314 -5306 7326 -5272
rect 7268 -5340 7326 -5306
rect 7268 -5374 7280 -5340
rect 7314 -5374 7326 -5340
rect 7268 -5408 7326 -5374
rect 7268 -5442 7280 -5408
rect 7314 -5442 7326 -5408
rect 7268 -5457 7326 -5442
rect 7526 -5272 7584 -5257
rect 7526 -5306 7538 -5272
rect 7572 -5306 7584 -5272
rect 7526 -5340 7584 -5306
rect 7526 -5374 7538 -5340
rect 7572 -5374 7584 -5340
rect 7526 -5408 7584 -5374
rect 7526 -5442 7538 -5408
rect 7572 -5442 7584 -5408
rect 7526 -5457 7584 -5442
rect 7784 -5272 7842 -5257
rect 7784 -5306 7796 -5272
rect 7830 -5306 7842 -5272
rect 7784 -5340 7842 -5306
rect 7784 -5374 7796 -5340
rect 7830 -5374 7842 -5340
rect 7784 -5408 7842 -5374
rect 7784 -5442 7796 -5408
rect 7830 -5442 7842 -5408
rect 7784 -5457 7842 -5442
rect 7978 -5272 8036 -5257
rect 7978 -5306 7990 -5272
rect 8024 -5306 8036 -5272
rect 7978 -5340 8036 -5306
rect 7978 -5374 7990 -5340
rect 8024 -5374 8036 -5340
rect 7978 -5408 8036 -5374
rect 7978 -5442 7990 -5408
rect 8024 -5442 8036 -5408
rect 7978 -5457 8036 -5442
rect 8236 -5272 8294 -5257
rect 8236 -5306 8248 -5272
rect 8282 -5306 8294 -5272
rect 8236 -5340 8294 -5306
rect 8236 -5374 8248 -5340
rect 8282 -5374 8294 -5340
rect 8236 -5408 8294 -5374
rect 8236 -5442 8248 -5408
rect 8282 -5442 8294 -5408
rect 8236 -5457 8294 -5442
rect 8494 -5272 8552 -5257
rect 8494 -5306 8506 -5272
rect 8540 -5306 8552 -5272
rect 8494 -5340 8552 -5306
rect 8494 -5374 8506 -5340
rect 8540 -5374 8552 -5340
rect 8494 -5408 8552 -5374
rect 8494 -5442 8506 -5408
rect 8540 -5442 8552 -5408
rect 8494 -5457 8552 -5442
rect 8752 -5272 8810 -5257
rect 8752 -5306 8764 -5272
rect 8798 -5306 8810 -5272
rect 8752 -5340 8810 -5306
rect 8752 -5374 8764 -5340
rect 8798 -5374 8810 -5340
rect 8752 -5408 8810 -5374
rect 8752 -5442 8764 -5408
rect 8798 -5442 8810 -5408
rect 8752 -5457 8810 -5442
rect 9010 -5272 9068 -5257
rect 9010 -5306 9022 -5272
rect 9056 -5306 9068 -5272
rect 9010 -5340 9068 -5306
rect 9010 -5374 9022 -5340
rect 9056 -5374 9068 -5340
rect 9010 -5408 9068 -5374
rect 9010 -5442 9022 -5408
rect 9056 -5442 9068 -5408
rect 9010 -5457 9068 -5442
rect 9204 -5272 9262 -5257
rect 9204 -5306 9216 -5272
rect 9250 -5306 9262 -5272
rect 9204 -5340 9262 -5306
rect 9204 -5374 9216 -5340
rect 9250 -5374 9262 -5340
rect 9204 -5408 9262 -5374
rect 9204 -5442 9216 -5408
rect 9250 -5442 9262 -5408
rect 9204 -5457 9262 -5442
rect 9462 -5272 9520 -5257
rect 9462 -5306 9474 -5272
rect 9508 -5306 9520 -5272
rect 9462 -5340 9520 -5306
rect 9462 -5374 9474 -5340
rect 9508 -5374 9520 -5340
rect 9462 -5408 9520 -5374
rect 9462 -5442 9474 -5408
rect 9508 -5442 9520 -5408
rect 9462 -5457 9520 -5442
rect 975 -5962 1033 -5947
rect 975 -5996 987 -5962
rect 1021 -5996 1033 -5962
rect 975 -6030 1033 -5996
rect 975 -6064 987 -6030
rect 1021 -6064 1033 -6030
rect 975 -6098 1033 -6064
rect 975 -6132 987 -6098
rect 1021 -6132 1033 -6098
rect 975 -6147 1033 -6132
rect 1233 -5962 1291 -5947
rect 1233 -5996 1245 -5962
rect 1279 -5996 1291 -5962
rect 1233 -6030 1291 -5996
rect 1233 -6064 1245 -6030
rect 1279 -6064 1291 -6030
rect 1233 -6098 1291 -6064
rect 1233 -6132 1245 -6098
rect 1279 -6132 1291 -6098
rect 1233 -6147 1291 -6132
rect 1427 -5962 1485 -5947
rect 1427 -5996 1439 -5962
rect 1473 -5996 1485 -5962
rect 1427 -6030 1485 -5996
rect 1427 -6064 1439 -6030
rect 1473 -6064 1485 -6030
rect 1427 -6098 1485 -6064
rect 1427 -6132 1439 -6098
rect 1473 -6132 1485 -6098
rect 1427 -6147 1485 -6132
rect 1685 -5962 1743 -5947
rect 1685 -5996 1697 -5962
rect 1731 -5996 1743 -5962
rect 1685 -6030 1743 -5996
rect 1685 -6064 1697 -6030
rect 1731 -6064 1743 -6030
rect 1685 -6098 1743 -6064
rect 1685 -6132 1697 -6098
rect 1731 -6132 1743 -6098
rect 1685 -6147 1743 -6132
rect 1943 -5962 2001 -5947
rect 1943 -5996 1955 -5962
rect 1989 -5996 2001 -5962
rect 1943 -6030 2001 -5996
rect 1943 -6064 1955 -6030
rect 1989 -6064 2001 -6030
rect 1943 -6098 2001 -6064
rect 1943 -6132 1955 -6098
rect 1989 -6132 2001 -6098
rect 1943 -6147 2001 -6132
rect 2201 -5962 2259 -5947
rect 2201 -5996 2213 -5962
rect 2247 -5996 2259 -5962
rect 2201 -6030 2259 -5996
rect 2201 -6064 2213 -6030
rect 2247 -6064 2259 -6030
rect 2201 -6098 2259 -6064
rect 2201 -6132 2213 -6098
rect 2247 -6132 2259 -6098
rect 2201 -6147 2259 -6132
rect 2459 -5962 2517 -5947
rect 2459 -5996 2471 -5962
rect 2505 -5996 2517 -5962
rect 2459 -6030 2517 -5996
rect 2459 -6064 2471 -6030
rect 2505 -6064 2517 -6030
rect 2459 -6098 2517 -6064
rect 2459 -6132 2471 -6098
rect 2505 -6132 2517 -6098
rect 2459 -6147 2517 -6132
rect 2653 -5962 2711 -5947
rect 2653 -5996 2665 -5962
rect 2699 -5996 2711 -5962
rect 2653 -6030 2711 -5996
rect 2653 -6064 2665 -6030
rect 2699 -6064 2711 -6030
rect 2653 -6098 2711 -6064
rect 2653 -6132 2665 -6098
rect 2699 -6132 2711 -6098
rect 2653 -6147 2711 -6132
rect 2911 -5962 2969 -5947
rect 2911 -5996 2923 -5962
rect 2957 -5996 2969 -5962
rect 2911 -6030 2969 -5996
rect 2911 -6064 2923 -6030
rect 2957 -6064 2969 -6030
rect 2911 -6098 2969 -6064
rect 2911 -6132 2923 -6098
rect 2957 -6132 2969 -6098
rect 2911 -6147 2969 -6132
rect 3169 -5962 3227 -5947
rect 3169 -5996 3181 -5962
rect 3215 -5996 3227 -5962
rect 3169 -6030 3227 -5996
rect 3169 -6064 3181 -6030
rect 3215 -6064 3227 -6030
rect 3169 -6098 3227 -6064
rect 3169 -6132 3181 -6098
rect 3215 -6132 3227 -6098
rect 3169 -6147 3227 -6132
rect 3427 -5962 3485 -5947
rect 3427 -5996 3439 -5962
rect 3473 -5996 3485 -5962
rect 3427 -6030 3485 -5996
rect 3427 -6064 3439 -6030
rect 3473 -6064 3485 -6030
rect 3427 -6098 3485 -6064
rect 3427 -6132 3439 -6098
rect 3473 -6132 3485 -6098
rect 3427 -6147 3485 -6132
rect 3621 -5962 3679 -5947
rect 3621 -5996 3633 -5962
rect 3667 -5996 3679 -5962
rect 3621 -6030 3679 -5996
rect 3621 -6064 3633 -6030
rect 3667 -6064 3679 -6030
rect 3621 -6098 3679 -6064
rect 3621 -6132 3633 -6098
rect 3667 -6132 3679 -6098
rect 3621 -6147 3679 -6132
rect 3879 -5962 3937 -5947
rect 3879 -5996 3891 -5962
rect 3925 -5996 3937 -5962
rect 3879 -6030 3937 -5996
rect 3879 -6064 3891 -6030
rect 3925 -6064 3937 -6030
rect 3879 -6098 3937 -6064
rect 3879 -6132 3891 -6098
rect 3925 -6132 3937 -6098
rect 3879 -6147 3937 -6132
rect 4137 -5962 4195 -5947
rect 4137 -5996 4149 -5962
rect 4183 -5996 4195 -5962
rect 4137 -6030 4195 -5996
rect 4137 -6064 4149 -6030
rect 4183 -6064 4195 -6030
rect 4137 -6098 4195 -6064
rect 4137 -6132 4149 -6098
rect 4183 -6132 4195 -6098
rect 4137 -6147 4195 -6132
rect 4395 -5962 4453 -5947
rect 4395 -5996 4407 -5962
rect 4441 -5996 4453 -5962
rect 4395 -6030 4453 -5996
rect 4395 -6064 4407 -6030
rect 4441 -6064 4453 -6030
rect 4395 -6098 4453 -6064
rect 4395 -6132 4407 -6098
rect 4441 -6132 4453 -6098
rect 4395 -6147 4453 -6132
rect 4653 -5962 4711 -5947
rect 4653 -5996 4665 -5962
rect 4699 -5996 4711 -5962
rect 4653 -6030 4711 -5996
rect 4653 -6064 4665 -6030
rect 4699 -6064 4711 -6030
rect 4653 -6098 4711 -6064
rect 4653 -6132 4665 -6098
rect 4699 -6132 4711 -6098
rect 4653 -6147 4711 -6132
rect 4847 -5962 4905 -5947
rect 4847 -5996 4859 -5962
rect 4893 -5996 4905 -5962
rect 4847 -6030 4905 -5996
rect 4847 -6064 4859 -6030
rect 4893 -6064 4905 -6030
rect 4847 -6098 4905 -6064
rect 4847 -6132 4859 -6098
rect 4893 -6132 4905 -6098
rect 4847 -6147 4905 -6132
rect 5105 -5962 5163 -5947
rect 5105 -5996 5117 -5962
rect 5151 -5996 5163 -5962
rect 5105 -6030 5163 -5996
rect 5105 -6064 5117 -6030
rect 5151 -6064 5163 -6030
rect 5105 -6098 5163 -6064
rect 5105 -6132 5117 -6098
rect 5151 -6132 5163 -6098
rect 5105 -6147 5163 -6132
rect 5333 -5962 5391 -5947
rect 5333 -5996 5345 -5962
rect 5379 -5996 5391 -5962
rect 5333 -6030 5391 -5996
rect 5333 -6064 5345 -6030
rect 5379 -6064 5391 -6030
rect 5333 -6098 5391 -6064
rect 5333 -6132 5345 -6098
rect 5379 -6132 5391 -6098
rect 5333 -6147 5391 -6132
rect 5591 -5962 5649 -5947
rect 5591 -5996 5603 -5962
rect 5637 -5996 5649 -5962
rect 5591 -6030 5649 -5996
rect 5591 -6064 5603 -6030
rect 5637 -6064 5649 -6030
rect 5591 -6098 5649 -6064
rect 5591 -6132 5603 -6098
rect 5637 -6132 5649 -6098
rect 5591 -6147 5649 -6132
rect 5784 -5962 5842 -5947
rect 5784 -5996 5796 -5962
rect 5830 -5996 5842 -5962
rect 5784 -6030 5842 -5996
rect 5784 -6064 5796 -6030
rect 5830 -6064 5842 -6030
rect 5784 -6098 5842 -6064
rect 5784 -6132 5796 -6098
rect 5830 -6132 5842 -6098
rect 5784 -6147 5842 -6132
rect 6042 -5962 6100 -5947
rect 6042 -5996 6054 -5962
rect 6088 -5996 6100 -5962
rect 6042 -6030 6100 -5996
rect 6042 -6064 6054 -6030
rect 6088 -6064 6100 -6030
rect 6042 -6098 6100 -6064
rect 6042 -6132 6054 -6098
rect 6088 -6132 6100 -6098
rect 6042 -6147 6100 -6132
rect 6300 -5962 6358 -5947
rect 6300 -5996 6312 -5962
rect 6346 -5996 6358 -5962
rect 6300 -6030 6358 -5996
rect 6300 -6064 6312 -6030
rect 6346 -6064 6358 -6030
rect 6300 -6098 6358 -6064
rect 6300 -6132 6312 -6098
rect 6346 -6132 6358 -6098
rect 6300 -6147 6358 -6132
rect 6558 -5962 6616 -5947
rect 6558 -5996 6570 -5962
rect 6604 -5996 6616 -5962
rect 6558 -6030 6616 -5996
rect 6558 -6064 6570 -6030
rect 6604 -6064 6616 -6030
rect 6558 -6098 6616 -6064
rect 6558 -6132 6570 -6098
rect 6604 -6132 6616 -6098
rect 6558 -6147 6616 -6132
rect 6816 -5962 6874 -5947
rect 6816 -5996 6828 -5962
rect 6862 -5996 6874 -5962
rect 6816 -6030 6874 -5996
rect 6816 -6064 6828 -6030
rect 6862 -6064 6874 -6030
rect 6816 -6098 6874 -6064
rect 6816 -6132 6828 -6098
rect 6862 -6132 6874 -6098
rect 6816 -6147 6874 -6132
rect 7010 -5962 7068 -5947
rect 7010 -5996 7022 -5962
rect 7056 -5996 7068 -5962
rect 7010 -6030 7068 -5996
rect 7010 -6064 7022 -6030
rect 7056 -6064 7068 -6030
rect 7010 -6098 7068 -6064
rect 7010 -6132 7022 -6098
rect 7056 -6132 7068 -6098
rect 7010 -6147 7068 -6132
rect 7268 -5962 7326 -5947
rect 7268 -5996 7280 -5962
rect 7314 -5996 7326 -5962
rect 7268 -6030 7326 -5996
rect 7268 -6064 7280 -6030
rect 7314 -6064 7326 -6030
rect 7268 -6098 7326 -6064
rect 7268 -6132 7280 -6098
rect 7314 -6132 7326 -6098
rect 7268 -6147 7326 -6132
rect 7526 -5962 7584 -5947
rect 7526 -5996 7538 -5962
rect 7572 -5996 7584 -5962
rect 7526 -6030 7584 -5996
rect 7526 -6064 7538 -6030
rect 7572 -6064 7584 -6030
rect 7526 -6098 7584 -6064
rect 7526 -6132 7538 -6098
rect 7572 -6132 7584 -6098
rect 7526 -6147 7584 -6132
rect 7784 -5962 7842 -5947
rect 7784 -5996 7796 -5962
rect 7830 -5996 7842 -5962
rect 7784 -6030 7842 -5996
rect 7784 -6064 7796 -6030
rect 7830 -6064 7842 -6030
rect 7784 -6098 7842 -6064
rect 7784 -6132 7796 -6098
rect 7830 -6132 7842 -6098
rect 7784 -6147 7842 -6132
rect 7978 -5962 8036 -5947
rect 7978 -5996 7990 -5962
rect 8024 -5996 8036 -5962
rect 7978 -6030 8036 -5996
rect 7978 -6064 7990 -6030
rect 8024 -6064 8036 -6030
rect 7978 -6098 8036 -6064
rect 7978 -6132 7990 -6098
rect 8024 -6132 8036 -6098
rect 7978 -6147 8036 -6132
rect 8236 -5962 8294 -5947
rect 8236 -5996 8248 -5962
rect 8282 -5996 8294 -5962
rect 8236 -6030 8294 -5996
rect 8236 -6064 8248 -6030
rect 8282 -6064 8294 -6030
rect 8236 -6098 8294 -6064
rect 8236 -6132 8248 -6098
rect 8282 -6132 8294 -6098
rect 8236 -6147 8294 -6132
rect 8494 -5962 8552 -5947
rect 8494 -5996 8506 -5962
rect 8540 -5996 8552 -5962
rect 8494 -6030 8552 -5996
rect 8494 -6064 8506 -6030
rect 8540 -6064 8552 -6030
rect 8494 -6098 8552 -6064
rect 8494 -6132 8506 -6098
rect 8540 -6132 8552 -6098
rect 8494 -6147 8552 -6132
rect 8752 -5962 8810 -5947
rect 8752 -5996 8764 -5962
rect 8798 -5996 8810 -5962
rect 8752 -6030 8810 -5996
rect 8752 -6064 8764 -6030
rect 8798 -6064 8810 -6030
rect 8752 -6098 8810 -6064
rect 8752 -6132 8764 -6098
rect 8798 -6132 8810 -6098
rect 8752 -6147 8810 -6132
rect 9010 -5962 9068 -5947
rect 9010 -5996 9022 -5962
rect 9056 -5996 9068 -5962
rect 9010 -6030 9068 -5996
rect 9010 -6064 9022 -6030
rect 9056 -6064 9068 -6030
rect 9010 -6098 9068 -6064
rect 9010 -6132 9022 -6098
rect 9056 -6132 9068 -6098
rect 9010 -6147 9068 -6132
rect 9204 -5962 9262 -5947
rect 9204 -5996 9216 -5962
rect 9250 -5996 9262 -5962
rect 9204 -6030 9262 -5996
rect 9204 -6064 9216 -6030
rect 9250 -6064 9262 -6030
rect 9204 -6098 9262 -6064
rect 9204 -6132 9216 -6098
rect 9250 -6132 9262 -6098
rect 9204 -6147 9262 -6132
rect 9462 -5962 9520 -5947
rect 9462 -5996 9474 -5962
rect 9508 -5996 9520 -5962
rect 9462 -6030 9520 -5996
rect 9462 -6064 9474 -6030
rect 9508 -6064 9520 -6030
rect 9462 -6098 9520 -6064
rect 9462 -6132 9474 -6098
rect 9508 -6132 9520 -6098
rect 9462 -6147 9520 -6132
rect 975 -6919 1033 -6904
rect 975 -6953 987 -6919
rect 1021 -6953 1033 -6919
rect 975 -6987 1033 -6953
rect 975 -7021 987 -6987
rect 1021 -7021 1033 -6987
rect 975 -7055 1033 -7021
rect 975 -7089 987 -7055
rect 1021 -7089 1033 -7055
rect 975 -7104 1033 -7089
rect 1233 -6919 1291 -6904
rect 1233 -6953 1245 -6919
rect 1279 -6953 1291 -6919
rect 1233 -6987 1291 -6953
rect 1233 -7021 1245 -6987
rect 1279 -7021 1291 -6987
rect 1233 -7055 1291 -7021
rect 1233 -7089 1245 -7055
rect 1279 -7089 1291 -7055
rect 1233 -7104 1291 -7089
rect 1427 -6919 1485 -6904
rect 1427 -6953 1439 -6919
rect 1473 -6953 1485 -6919
rect 1427 -6987 1485 -6953
rect 1427 -7021 1439 -6987
rect 1473 -7021 1485 -6987
rect 1427 -7055 1485 -7021
rect 1427 -7089 1439 -7055
rect 1473 -7089 1485 -7055
rect 1427 -7104 1485 -7089
rect 1685 -6919 1743 -6904
rect 1685 -6953 1697 -6919
rect 1731 -6953 1743 -6919
rect 1685 -6987 1743 -6953
rect 1685 -7021 1697 -6987
rect 1731 -7021 1743 -6987
rect 1685 -7055 1743 -7021
rect 1685 -7089 1697 -7055
rect 1731 -7089 1743 -7055
rect 1685 -7104 1743 -7089
rect 1943 -6919 2001 -6904
rect 1943 -6953 1955 -6919
rect 1989 -6953 2001 -6919
rect 1943 -6987 2001 -6953
rect 1943 -7021 1955 -6987
rect 1989 -7021 2001 -6987
rect 1943 -7055 2001 -7021
rect 1943 -7089 1955 -7055
rect 1989 -7089 2001 -7055
rect 1943 -7104 2001 -7089
rect 2201 -6919 2259 -6904
rect 2201 -6953 2213 -6919
rect 2247 -6953 2259 -6919
rect 2201 -6987 2259 -6953
rect 2201 -7021 2213 -6987
rect 2247 -7021 2259 -6987
rect 2201 -7055 2259 -7021
rect 2201 -7089 2213 -7055
rect 2247 -7089 2259 -7055
rect 2201 -7104 2259 -7089
rect 2459 -6919 2517 -6904
rect 2459 -6953 2471 -6919
rect 2505 -6953 2517 -6919
rect 2459 -6987 2517 -6953
rect 2459 -7021 2471 -6987
rect 2505 -7021 2517 -6987
rect 2459 -7055 2517 -7021
rect 2459 -7089 2471 -7055
rect 2505 -7089 2517 -7055
rect 2459 -7104 2517 -7089
rect 2653 -6919 2711 -6904
rect 2653 -6953 2665 -6919
rect 2699 -6953 2711 -6919
rect 2653 -6987 2711 -6953
rect 2653 -7021 2665 -6987
rect 2699 -7021 2711 -6987
rect 2653 -7055 2711 -7021
rect 2653 -7089 2665 -7055
rect 2699 -7089 2711 -7055
rect 2653 -7104 2711 -7089
rect 2911 -6919 2969 -6904
rect 2911 -6953 2923 -6919
rect 2957 -6953 2969 -6919
rect 2911 -6987 2969 -6953
rect 2911 -7021 2923 -6987
rect 2957 -7021 2969 -6987
rect 2911 -7055 2969 -7021
rect 2911 -7089 2923 -7055
rect 2957 -7089 2969 -7055
rect 2911 -7104 2969 -7089
rect 3169 -6919 3227 -6904
rect 3169 -6953 3181 -6919
rect 3215 -6953 3227 -6919
rect 3169 -6987 3227 -6953
rect 3169 -7021 3181 -6987
rect 3215 -7021 3227 -6987
rect 3169 -7055 3227 -7021
rect 3169 -7089 3181 -7055
rect 3215 -7089 3227 -7055
rect 3169 -7104 3227 -7089
rect 3427 -6919 3485 -6904
rect 3427 -6953 3439 -6919
rect 3473 -6953 3485 -6919
rect 3427 -6987 3485 -6953
rect 3427 -7021 3439 -6987
rect 3473 -7021 3485 -6987
rect 3427 -7055 3485 -7021
rect 3427 -7089 3439 -7055
rect 3473 -7089 3485 -7055
rect 3427 -7104 3485 -7089
rect 3621 -6919 3679 -6904
rect 3621 -6953 3633 -6919
rect 3667 -6953 3679 -6919
rect 3621 -6987 3679 -6953
rect 3621 -7021 3633 -6987
rect 3667 -7021 3679 -6987
rect 3621 -7055 3679 -7021
rect 3621 -7089 3633 -7055
rect 3667 -7089 3679 -7055
rect 3621 -7104 3679 -7089
rect 3879 -6919 3937 -6904
rect 3879 -6953 3891 -6919
rect 3925 -6953 3937 -6919
rect 3879 -6987 3937 -6953
rect 3879 -7021 3891 -6987
rect 3925 -7021 3937 -6987
rect 3879 -7055 3937 -7021
rect 3879 -7089 3891 -7055
rect 3925 -7089 3937 -7055
rect 3879 -7104 3937 -7089
rect 4137 -6919 4195 -6904
rect 4137 -6953 4149 -6919
rect 4183 -6953 4195 -6919
rect 4137 -6987 4195 -6953
rect 4137 -7021 4149 -6987
rect 4183 -7021 4195 -6987
rect 4137 -7055 4195 -7021
rect 4137 -7089 4149 -7055
rect 4183 -7089 4195 -7055
rect 4137 -7104 4195 -7089
rect 4395 -6919 4453 -6904
rect 4395 -6953 4407 -6919
rect 4441 -6953 4453 -6919
rect 4395 -6987 4453 -6953
rect 4395 -7021 4407 -6987
rect 4441 -7021 4453 -6987
rect 4395 -7055 4453 -7021
rect 4395 -7089 4407 -7055
rect 4441 -7089 4453 -7055
rect 4395 -7104 4453 -7089
rect 4653 -6919 4711 -6904
rect 4653 -6953 4665 -6919
rect 4699 -6953 4711 -6919
rect 4653 -6987 4711 -6953
rect 4653 -7021 4665 -6987
rect 4699 -7021 4711 -6987
rect 4653 -7055 4711 -7021
rect 4653 -7089 4665 -7055
rect 4699 -7089 4711 -7055
rect 4653 -7104 4711 -7089
rect 4847 -6919 4905 -6904
rect 4847 -6953 4859 -6919
rect 4893 -6953 4905 -6919
rect 4847 -6987 4905 -6953
rect 4847 -7021 4859 -6987
rect 4893 -7021 4905 -6987
rect 4847 -7055 4905 -7021
rect 4847 -7089 4859 -7055
rect 4893 -7089 4905 -7055
rect 4847 -7104 4905 -7089
rect 5105 -6919 5163 -6904
rect 5105 -6953 5117 -6919
rect 5151 -6953 5163 -6919
rect 5105 -6987 5163 -6953
rect 5105 -7021 5117 -6987
rect 5151 -7021 5163 -6987
rect 5105 -7055 5163 -7021
rect 5105 -7089 5117 -7055
rect 5151 -7089 5163 -7055
rect 5105 -7104 5163 -7089
rect 5333 -6919 5391 -6904
rect 5333 -6953 5345 -6919
rect 5379 -6953 5391 -6919
rect 5333 -6987 5391 -6953
rect 5333 -7021 5345 -6987
rect 5379 -7021 5391 -6987
rect 5333 -7055 5391 -7021
rect 5333 -7089 5345 -7055
rect 5379 -7089 5391 -7055
rect 5333 -7104 5391 -7089
rect 5591 -6919 5649 -6904
rect 5591 -6953 5603 -6919
rect 5637 -6953 5649 -6919
rect 5591 -6987 5649 -6953
rect 5591 -7021 5603 -6987
rect 5637 -7021 5649 -6987
rect 5591 -7055 5649 -7021
rect 5591 -7089 5603 -7055
rect 5637 -7089 5649 -7055
rect 5591 -7104 5649 -7089
rect 5784 -6919 5842 -6904
rect 5784 -6953 5796 -6919
rect 5830 -6953 5842 -6919
rect 5784 -6987 5842 -6953
rect 5784 -7021 5796 -6987
rect 5830 -7021 5842 -6987
rect 5784 -7055 5842 -7021
rect 5784 -7089 5796 -7055
rect 5830 -7089 5842 -7055
rect 5784 -7104 5842 -7089
rect 6042 -6919 6100 -6904
rect 6042 -6953 6054 -6919
rect 6088 -6953 6100 -6919
rect 6042 -6987 6100 -6953
rect 6042 -7021 6054 -6987
rect 6088 -7021 6100 -6987
rect 6042 -7055 6100 -7021
rect 6042 -7089 6054 -7055
rect 6088 -7089 6100 -7055
rect 6042 -7104 6100 -7089
rect 6300 -6919 6358 -6904
rect 6300 -6953 6312 -6919
rect 6346 -6953 6358 -6919
rect 6300 -6987 6358 -6953
rect 6300 -7021 6312 -6987
rect 6346 -7021 6358 -6987
rect 6300 -7055 6358 -7021
rect 6300 -7089 6312 -7055
rect 6346 -7089 6358 -7055
rect 6300 -7104 6358 -7089
rect 6558 -6919 6616 -6904
rect 6558 -6953 6570 -6919
rect 6604 -6953 6616 -6919
rect 6558 -6987 6616 -6953
rect 6558 -7021 6570 -6987
rect 6604 -7021 6616 -6987
rect 6558 -7055 6616 -7021
rect 6558 -7089 6570 -7055
rect 6604 -7089 6616 -7055
rect 6558 -7104 6616 -7089
rect 6816 -6919 6874 -6904
rect 6816 -6953 6828 -6919
rect 6862 -6953 6874 -6919
rect 6816 -6987 6874 -6953
rect 6816 -7021 6828 -6987
rect 6862 -7021 6874 -6987
rect 6816 -7055 6874 -7021
rect 6816 -7089 6828 -7055
rect 6862 -7089 6874 -7055
rect 6816 -7104 6874 -7089
rect 7010 -6919 7068 -6904
rect 7010 -6953 7022 -6919
rect 7056 -6953 7068 -6919
rect 7010 -6987 7068 -6953
rect 7010 -7021 7022 -6987
rect 7056 -7021 7068 -6987
rect 7010 -7055 7068 -7021
rect 7010 -7089 7022 -7055
rect 7056 -7089 7068 -7055
rect 7010 -7104 7068 -7089
rect 7268 -6919 7326 -6904
rect 7268 -6953 7280 -6919
rect 7314 -6953 7326 -6919
rect 7268 -6987 7326 -6953
rect 7268 -7021 7280 -6987
rect 7314 -7021 7326 -6987
rect 7268 -7055 7326 -7021
rect 7268 -7089 7280 -7055
rect 7314 -7089 7326 -7055
rect 7268 -7104 7326 -7089
rect 7526 -6919 7584 -6904
rect 7526 -6953 7538 -6919
rect 7572 -6953 7584 -6919
rect 7526 -6987 7584 -6953
rect 7526 -7021 7538 -6987
rect 7572 -7021 7584 -6987
rect 7526 -7055 7584 -7021
rect 7526 -7089 7538 -7055
rect 7572 -7089 7584 -7055
rect 7526 -7104 7584 -7089
rect 7784 -6919 7842 -6904
rect 7784 -6953 7796 -6919
rect 7830 -6953 7842 -6919
rect 7784 -6987 7842 -6953
rect 7784 -7021 7796 -6987
rect 7830 -7021 7842 -6987
rect 7784 -7055 7842 -7021
rect 7784 -7089 7796 -7055
rect 7830 -7089 7842 -7055
rect 7784 -7104 7842 -7089
rect 7978 -6919 8036 -6904
rect 7978 -6953 7990 -6919
rect 8024 -6953 8036 -6919
rect 7978 -6987 8036 -6953
rect 7978 -7021 7990 -6987
rect 8024 -7021 8036 -6987
rect 7978 -7055 8036 -7021
rect 7978 -7089 7990 -7055
rect 8024 -7089 8036 -7055
rect 7978 -7104 8036 -7089
rect 8236 -6919 8294 -6904
rect 8236 -6953 8248 -6919
rect 8282 -6953 8294 -6919
rect 8236 -6987 8294 -6953
rect 8236 -7021 8248 -6987
rect 8282 -7021 8294 -6987
rect 8236 -7055 8294 -7021
rect 8236 -7089 8248 -7055
rect 8282 -7089 8294 -7055
rect 8236 -7104 8294 -7089
rect 8494 -6919 8552 -6904
rect 8494 -6953 8506 -6919
rect 8540 -6953 8552 -6919
rect 8494 -6987 8552 -6953
rect 8494 -7021 8506 -6987
rect 8540 -7021 8552 -6987
rect 8494 -7055 8552 -7021
rect 8494 -7089 8506 -7055
rect 8540 -7089 8552 -7055
rect 8494 -7104 8552 -7089
rect 8752 -6919 8810 -6904
rect 8752 -6953 8764 -6919
rect 8798 -6953 8810 -6919
rect 8752 -6987 8810 -6953
rect 8752 -7021 8764 -6987
rect 8798 -7021 8810 -6987
rect 8752 -7055 8810 -7021
rect 8752 -7089 8764 -7055
rect 8798 -7089 8810 -7055
rect 8752 -7104 8810 -7089
rect 9010 -6919 9068 -6904
rect 9010 -6953 9022 -6919
rect 9056 -6953 9068 -6919
rect 9010 -6987 9068 -6953
rect 9010 -7021 9022 -6987
rect 9056 -7021 9068 -6987
rect 9010 -7055 9068 -7021
rect 9010 -7089 9022 -7055
rect 9056 -7089 9068 -7055
rect 9010 -7104 9068 -7089
rect 9204 -6919 9262 -6904
rect 9204 -6953 9216 -6919
rect 9250 -6953 9262 -6919
rect 9204 -6987 9262 -6953
rect 9204 -7021 9216 -6987
rect 9250 -7021 9262 -6987
rect 9204 -7055 9262 -7021
rect 9204 -7089 9216 -7055
rect 9250 -7089 9262 -7055
rect 9204 -7104 9262 -7089
rect 9462 -6919 9520 -6904
rect 9462 -6953 9474 -6919
rect 9508 -6953 9520 -6919
rect 9462 -6987 9520 -6953
rect 9462 -7021 9474 -6987
rect 9508 -7021 9520 -6987
rect 9462 -7055 9520 -7021
rect 9462 -7089 9474 -7055
rect 9508 -7089 9520 -7055
rect 9462 -7104 9520 -7089
rect 975 -7609 1033 -7594
rect 975 -7643 987 -7609
rect 1021 -7643 1033 -7609
rect 975 -7677 1033 -7643
rect 975 -7711 987 -7677
rect 1021 -7711 1033 -7677
rect 975 -7745 1033 -7711
rect 975 -7779 987 -7745
rect 1021 -7779 1033 -7745
rect 975 -7794 1033 -7779
rect 1233 -7609 1291 -7594
rect 1233 -7643 1245 -7609
rect 1279 -7643 1291 -7609
rect 1233 -7677 1291 -7643
rect 1233 -7711 1245 -7677
rect 1279 -7711 1291 -7677
rect 1233 -7745 1291 -7711
rect 1233 -7779 1245 -7745
rect 1279 -7779 1291 -7745
rect 1233 -7794 1291 -7779
rect 1427 -7609 1485 -7594
rect 1427 -7643 1439 -7609
rect 1473 -7643 1485 -7609
rect 1427 -7677 1485 -7643
rect 1427 -7711 1439 -7677
rect 1473 -7711 1485 -7677
rect 1427 -7745 1485 -7711
rect 1427 -7779 1439 -7745
rect 1473 -7779 1485 -7745
rect 1427 -7794 1485 -7779
rect 1685 -7609 1743 -7594
rect 1685 -7643 1697 -7609
rect 1731 -7643 1743 -7609
rect 1685 -7677 1743 -7643
rect 1685 -7711 1697 -7677
rect 1731 -7711 1743 -7677
rect 1685 -7745 1743 -7711
rect 1685 -7779 1697 -7745
rect 1731 -7779 1743 -7745
rect 1685 -7794 1743 -7779
rect 1943 -7609 2001 -7594
rect 1943 -7643 1955 -7609
rect 1989 -7643 2001 -7609
rect 1943 -7677 2001 -7643
rect 1943 -7711 1955 -7677
rect 1989 -7711 2001 -7677
rect 1943 -7745 2001 -7711
rect 1943 -7779 1955 -7745
rect 1989 -7779 2001 -7745
rect 1943 -7794 2001 -7779
rect 2201 -7609 2259 -7594
rect 2201 -7643 2213 -7609
rect 2247 -7643 2259 -7609
rect 2201 -7677 2259 -7643
rect 2201 -7711 2213 -7677
rect 2247 -7711 2259 -7677
rect 2201 -7745 2259 -7711
rect 2201 -7779 2213 -7745
rect 2247 -7779 2259 -7745
rect 2201 -7794 2259 -7779
rect 2459 -7609 2517 -7594
rect 2459 -7643 2471 -7609
rect 2505 -7643 2517 -7609
rect 2459 -7677 2517 -7643
rect 2459 -7711 2471 -7677
rect 2505 -7711 2517 -7677
rect 2459 -7745 2517 -7711
rect 2459 -7779 2471 -7745
rect 2505 -7779 2517 -7745
rect 2459 -7794 2517 -7779
rect 2653 -7609 2711 -7594
rect 2653 -7643 2665 -7609
rect 2699 -7643 2711 -7609
rect 2653 -7677 2711 -7643
rect 2653 -7711 2665 -7677
rect 2699 -7711 2711 -7677
rect 2653 -7745 2711 -7711
rect 2653 -7779 2665 -7745
rect 2699 -7779 2711 -7745
rect 2653 -7794 2711 -7779
rect 2911 -7609 2969 -7594
rect 2911 -7643 2923 -7609
rect 2957 -7643 2969 -7609
rect 2911 -7677 2969 -7643
rect 2911 -7711 2923 -7677
rect 2957 -7711 2969 -7677
rect 2911 -7745 2969 -7711
rect 2911 -7779 2923 -7745
rect 2957 -7779 2969 -7745
rect 2911 -7794 2969 -7779
rect 3169 -7609 3227 -7594
rect 3169 -7643 3181 -7609
rect 3215 -7643 3227 -7609
rect 3169 -7677 3227 -7643
rect 3169 -7711 3181 -7677
rect 3215 -7711 3227 -7677
rect 3169 -7745 3227 -7711
rect 3169 -7779 3181 -7745
rect 3215 -7779 3227 -7745
rect 3169 -7794 3227 -7779
rect 3427 -7609 3485 -7594
rect 3427 -7643 3439 -7609
rect 3473 -7643 3485 -7609
rect 3427 -7677 3485 -7643
rect 3427 -7711 3439 -7677
rect 3473 -7711 3485 -7677
rect 3427 -7745 3485 -7711
rect 3427 -7779 3439 -7745
rect 3473 -7779 3485 -7745
rect 3427 -7794 3485 -7779
rect 3621 -7609 3679 -7594
rect 3621 -7643 3633 -7609
rect 3667 -7643 3679 -7609
rect 3621 -7677 3679 -7643
rect 3621 -7711 3633 -7677
rect 3667 -7711 3679 -7677
rect 3621 -7745 3679 -7711
rect 3621 -7779 3633 -7745
rect 3667 -7779 3679 -7745
rect 3621 -7794 3679 -7779
rect 3879 -7609 3937 -7594
rect 3879 -7643 3891 -7609
rect 3925 -7643 3937 -7609
rect 3879 -7677 3937 -7643
rect 3879 -7711 3891 -7677
rect 3925 -7711 3937 -7677
rect 3879 -7745 3937 -7711
rect 3879 -7779 3891 -7745
rect 3925 -7779 3937 -7745
rect 3879 -7794 3937 -7779
rect 4137 -7609 4195 -7594
rect 4137 -7643 4149 -7609
rect 4183 -7643 4195 -7609
rect 4137 -7677 4195 -7643
rect 4137 -7711 4149 -7677
rect 4183 -7711 4195 -7677
rect 4137 -7745 4195 -7711
rect 4137 -7779 4149 -7745
rect 4183 -7779 4195 -7745
rect 4137 -7794 4195 -7779
rect 4395 -7609 4453 -7594
rect 4395 -7643 4407 -7609
rect 4441 -7643 4453 -7609
rect 4395 -7677 4453 -7643
rect 4395 -7711 4407 -7677
rect 4441 -7711 4453 -7677
rect 4395 -7745 4453 -7711
rect 4395 -7779 4407 -7745
rect 4441 -7779 4453 -7745
rect 4395 -7794 4453 -7779
rect 4653 -7609 4711 -7594
rect 4653 -7643 4665 -7609
rect 4699 -7643 4711 -7609
rect 4653 -7677 4711 -7643
rect 4653 -7711 4665 -7677
rect 4699 -7711 4711 -7677
rect 4653 -7745 4711 -7711
rect 4653 -7779 4665 -7745
rect 4699 -7779 4711 -7745
rect 4653 -7794 4711 -7779
rect 4847 -7609 4905 -7594
rect 4847 -7643 4859 -7609
rect 4893 -7643 4905 -7609
rect 4847 -7677 4905 -7643
rect 4847 -7711 4859 -7677
rect 4893 -7711 4905 -7677
rect 4847 -7745 4905 -7711
rect 4847 -7779 4859 -7745
rect 4893 -7779 4905 -7745
rect 4847 -7794 4905 -7779
rect 5105 -7609 5163 -7594
rect 5105 -7643 5117 -7609
rect 5151 -7643 5163 -7609
rect 5105 -7677 5163 -7643
rect 5105 -7711 5117 -7677
rect 5151 -7711 5163 -7677
rect 5105 -7745 5163 -7711
rect 5105 -7779 5117 -7745
rect 5151 -7779 5163 -7745
rect 5105 -7794 5163 -7779
rect 5333 -7609 5391 -7594
rect 5333 -7643 5345 -7609
rect 5379 -7643 5391 -7609
rect 5333 -7677 5391 -7643
rect 5333 -7711 5345 -7677
rect 5379 -7711 5391 -7677
rect 5333 -7745 5391 -7711
rect 5333 -7779 5345 -7745
rect 5379 -7779 5391 -7745
rect 5333 -7794 5391 -7779
rect 5591 -7609 5649 -7594
rect 5591 -7643 5603 -7609
rect 5637 -7643 5649 -7609
rect 5591 -7677 5649 -7643
rect 5591 -7711 5603 -7677
rect 5637 -7711 5649 -7677
rect 5591 -7745 5649 -7711
rect 5591 -7779 5603 -7745
rect 5637 -7779 5649 -7745
rect 5591 -7794 5649 -7779
rect 5784 -7609 5842 -7594
rect 5784 -7643 5796 -7609
rect 5830 -7643 5842 -7609
rect 5784 -7677 5842 -7643
rect 5784 -7711 5796 -7677
rect 5830 -7711 5842 -7677
rect 5784 -7745 5842 -7711
rect 5784 -7779 5796 -7745
rect 5830 -7779 5842 -7745
rect 5784 -7794 5842 -7779
rect 6042 -7609 6100 -7594
rect 6042 -7643 6054 -7609
rect 6088 -7643 6100 -7609
rect 6042 -7677 6100 -7643
rect 6042 -7711 6054 -7677
rect 6088 -7711 6100 -7677
rect 6042 -7745 6100 -7711
rect 6042 -7779 6054 -7745
rect 6088 -7779 6100 -7745
rect 6042 -7794 6100 -7779
rect 6300 -7609 6358 -7594
rect 6300 -7643 6312 -7609
rect 6346 -7643 6358 -7609
rect 6300 -7677 6358 -7643
rect 6300 -7711 6312 -7677
rect 6346 -7711 6358 -7677
rect 6300 -7745 6358 -7711
rect 6300 -7779 6312 -7745
rect 6346 -7779 6358 -7745
rect 6300 -7794 6358 -7779
rect 6558 -7609 6616 -7594
rect 6558 -7643 6570 -7609
rect 6604 -7643 6616 -7609
rect 6558 -7677 6616 -7643
rect 6558 -7711 6570 -7677
rect 6604 -7711 6616 -7677
rect 6558 -7745 6616 -7711
rect 6558 -7779 6570 -7745
rect 6604 -7779 6616 -7745
rect 6558 -7794 6616 -7779
rect 6816 -7609 6874 -7594
rect 6816 -7643 6828 -7609
rect 6862 -7643 6874 -7609
rect 6816 -7677 6874 -7643
rect 6816 -7711 6828 -7677
rect 6862 -7711 6874 -7677
rect 6816 -7745 6874 -7711
rect 6816 -7779 6828 -7745
rect 6862 -7779 6874 -7745
rect 6816 -7794 6874 -7779
rect 7010 -7609 7068 -7594
rect 7010 -7643 7022 -7609
rect 7056 -7643 7068 -7609
rect 7010 -7677 7068 -7643
rect 7010 -7711 7022 -7677
rect 7056 -7711 7068 -7677
rect 7010 -7745 7068 -7711
rect 7010 -7779 7022 -7745
rect 7056 -7779 7068 -7745
rect 7010 -7794 7068 -7779
rect 7268 -7609 7326 -7594
rect 7268 -7643 7280 -7609
rect 7314 -7643 7326 -7609
rect 7268 -7677 7326 -7643
rect 7268 -7711 7280 -7677
rect 7314 -7711 7326 -7677
rect 7268 -7745 7326 -7711
rect 7268 -7779 7280 -7745
rect 7314 -7779 7326 -7745
rect 7268 -7794 7326 -7779
rect 7526 -7609 7584 -7594
rect 7526 -7643 7538 -7609
rect 7572 -7643 7584 -7609
rect 7526 -7677 7584 -7643
rect 7526 -7711 7538 -7677
rect 7572 -7711 7584 -7677
rect 7526 -7745 7584 -7711
rect 7526 -7779 7538 -7745
rect 7572 -7779 7584 -7745
rect 7526 -7794 7584 -7779
rect 7784 -7609 7842 -7594
rect 7784 -7643 7796 -7609
rect 7830 -7643 7842 -7609
rect 7784 -7677 7842 -7643
rect 7784 -7711 7796 -7677
rect 7830 -7711 7842 -7677
rect 7784 -7745 7842 -7711
rect 7784 -7779 7796 -7745
rect 7830 -7779 7842 -7745
rect 7784 -7794 7842 -7779
rect 7978 -7609 8036 -7594
rect 7978 -7643 7990 -7609
rect 8024 -7643 8036 -7609
rect 7978 -7677 8036 -7643
rect 7978 -7711 7990 -7677
rect 8024 -7711 8036 -7677
rect 7978 -7745 8036 -7711
rect 7978 -7779 7990 -7745
rect 8024 -7779 8036 -7745
rect 7978 -7794 8036 -7779
rect 8236 -7609 8294 -7594
rect 8236 -7643 8248 -7609
rect 8282 -7643 8294 -7609
rect 8236 -7677 8294 -7643
rect 8236 -7711 8248 -7677
rect 8282 -7711 8294 -7677
rect 8236 -7745 8294 -7711
rect 8236 -7779 8248 -7745
rect 8282 -7779 8294 -7745
rect 8236 -7794 8294 -7779
rect 8494 -7609 8552 -7594
rect 8494 -7643 8506 -7609
rect 8540 -7643 8552 -7609
rect 8494 -7677 8552 -7643
rect 8494 -7711 8506 -7677
rect 8540 -7711 8552 -7677
rect 8494 -7745 8552 -7711
rect 8494 -7779 8506 -7745
rect 8540 -7779 8552 -7745
rect 8494 -7794 8552 -7779
rect 8752 -7609 8810 -7594
rect 8752 -7643 8764 -7609
rect 8798 -7643 8810 -7609
rect 8752 -7677 8810 -7643
rect 8752 -7711 8764 -7677
rect 8798 -7711 8810 -7677
rect 8752 -7745 8810 -7711
rect 8752 -7779 8764 -7745
rect 8798 -7779 8810 -7745
rect 8752 -7794 8810 -7779
rect 9010 -7609 9068 -7594
rect 9010 -7643 9022 -7609
rect 9056 -7643 9068 -7609
rect 9010 -7677 9068 -7643
rect 9010 -7711 9022 -7677
rect 9056 -7711 9068 -7677
rect 9010 -7745 9068 -7711
rect 9010 -7779 9022 -7745
rect 9056 -7779 9068 -7745
rect 9010 -7794 9068 -7779
rect 9204 -7609 9262 -7594
rect 9204 -7643 9216 -7609
rect 9250 -7643 9262 -7609
rect 9204 -7677 9262 -7643
rect 9204 -7711 9216 -7677
rect 9250 -7711 9262 -7677
rect 9204 -7745 9262 -7711
rect 9204 -7779 9216 -7745
rect 9250 -7779 9262 -7745
rect 9204 -7794 9262 -7779
rect 9462 -7609 9520 -7594
rect 9462 -7643 9474 -7609
rect 9508 -7643 9520 -7609
rect 9462 -7677 9520 -7643
rect 9462 -7711 9474 -7677
rect 9508 -7711 9520 -7677
rect 9462 -7745 9520 -7711
rect 9462 -7779 9474 -7745
rect 9508 -7779 9520 -7745
rect 9462 -7794 9520 -7779
rect 975 -8553 1033 -8538
rect 975 -8587 987 -8553
rect 1021 -8587 1033 -8553
rect 975 -8621 1033 -8587
rect 975 -8655 987 -8621
rect 1021 -8655 1033 -8621
rect 975 -8689 1033 -8655
rect 975 -8723 987 -8689
rect 1021 -8723 1033 -8689
rect 975 -8738 1033 -8723
rect 1233 -8553 1291 -8538
rect 1233 -8587 1245 -8553
rect 1279 -8587 1291 -8553
rect 1233 -8621 1291 -8587
rect 1233 -8655 1245 -8621
rect 1279 -8655 1291 -8621
rect 1233 -8689 1291 -8655
rect 1233 -8723 1245 -8689
rect 1279 -8723 1291 -8689
rect 1233 -8738 1291 -8723
rect 1427 -8553 1485 -8538
rect 1427 -8587 1439 -8553
rect 1473 -8587 1485 -8553
rect 1427 -8621 1485 -8587
rect 1427 -8655 1439 -8621
rect 1473 -8655 1485 -8621
rect 1427 -8689 1485 -8655
rect 1427 -8723 1439 -8689
rect 1473 -8723 1485 -8689
rect 1427 -8738 1485 -8723
rect 1685 -8553 1743 -8538
rect 1685 -8587 1697 -8553
rect 1731 -8587 1743 -8553
rect 1685 -8621 1743 -8587
rect 1685 -8655 1697 -8621
rect 1731 -8655 1743 -8621
rect 1685 -8689 1743 -8655
rect 1685 -8723 1697 -8689
rect 1731 -8723 1743 -8689
rect 1685 -8738 1743 -8723
rect 1943 -8553 2001 -8538
rect 1943 -8587 1955 -8553
rect 1989 -8587 2001 -8553
rect 1943 -8621 2001 -8587
rect 1943 -8655 1955 -8621
rect 1989 -8655 2001 -8621
rect 1943 -8689 2001 -8655
rect 1943 -8723 1955 -8689
rect 1989 -8723 2001 -8689
rect 1943 -8738 2001 -8723
rect 2201 -8553 2259 -8538
rect 2201 -8587 2213 -8553
rect 2247 -8587 2259 -8553
rect 2201 -8621 2259 -8587
rect 2201 -8655 2213 -8621
rect 2247 -8655 2259 -8621
rect 2201 -8689 2259 -8655
rect 2201 -8723 2213 -8689
rect 2247 -8723 2259 -8689
rect 2201 -8738 2259 -8723
rect 2459 -8553 2517 -8538
rect 2459 -8587 2471 -8553
rect 2505 -8587 2517 -8553
rect 2459 -8621 2517 -8587
rect 2459 -8655 2471 -8621
rect 2505 -8655 2517 -8621
rect 2459 -8689 2517 -8655
rect 2459 -8723 2471 -8689
rect 2505 -8723 2517 -8689
rect 2459 -8738 2517 -8723
rect 2653 -8553 2711 -8538
rect 2653 -8587 2665 -8553
rect 2699 -8587 2711 -8553
rect 2653 -8621 2711 -8587
rect 2653 -8655 2665 -8621
rect 2699 -8655 2711 -8621
rect 2653 -8689 2711 -8655
rect 2653 -8723 2665 -8689
rect 2699 -8723 2711 -8689
rect 2653 -8738 2711 -8723
rect 2911 -8553 2969 -8538
rect 2911 -8587 2923 -8553
rect 2957 -8587 2969 -8553
rect 2911 -8621 2969 -8587
rect 2911 -8655 2923 -8621
rect 2957 -8655 2969 -8621
rect 2911 -8689 2969 -8655
rect 2911 -8723 2923 -8689
rect 2957 -8723 2969 -8689
rect 2911 -8738 2969 -8723
rect 3169 -8553 3227 -8538
rect 3169 -8587 3181 -8553
rect 3215 -8587 3227 -8553
rect 3169 -8621 3227 -8587
rect 3169 -8655 3181 -8621
rect 3215 -8655 3227 -8621
rect 3169 -8689 3227 -8655
rect 3169 -8723 3181 -8689
rect 3215 -8723 3227 -8689
rect 3169 -8738 3227 -8723
rect 3427 -8553 3485 -8538
rect 3427 -8587 3439 -8553
rect 3473 -8587 3485 -8553
rect 3427 -8621 3485 -8587
rect 3427 -8655 3439 -8621
rect 3473 -8655 3485 -8621
rect 3427 -8689 3485 -8655
rect 3427 -8723 3439 -8689
rect 3473 -8723 3485 -8689
rect 3427 -8738 3485 -8723
rect 3621 -8553 3679 -8538
rect 3621 -8587 3633 -8553
rect 3667 -8587 3679 -8553
rect 3621 -8621 3679 -8587
rect 3621 -8655 3633 -8621
rect 3667 -8655 3679 -8621
rect 3621 -8689 3679 -8655
rect 3621 -8723 3633 -8689
rect 3667 -8723 3679 -8689
rect 3621 -8738 3679 -8723
rect 3879 -8553 3937 -8538
rect 3879 -8587 3891 -8553
rect 3925 -8587 3937 -8553
rect 3879 -8621 3937 -8587
rect 3879 -8655 3891 -8621
rect 3925 -8655 3937 -8621
rect 3879 -8689 3937 -8655
rect 3879 -8723 3891 -8689
rect 3925 -8723 3937 -8689
rect 3879 -8738 3937 -8723
rect 4137 -8553 4195 -8538
rect 4137 -8587 4149 -8553
rect 4183 -8587 4195 -8553
rect 4137 -8621 4195 -8587
rect 4137 -8655 4149 -8621
rect 4183 -8655 4195 -8621
rect 4137 -8689 4195 -8655
rect 4137 -8723 4149 -8689
rect 4183 -8723 4195 -8689
rect 4137 -8738 4195 -8723
rect 4395 -8553 4453 -8538
rect 4395 -8587 4407 -8553
rect 4441 -8587 4453 -8553
rect 4395 -8621 4453 -8587
rect 4395 -8655 4407 -8621
rect 4441 -8655 4453 -8621
rect 4395 -8689 4453 -8655
rect 4395 -8723 4407 -8689
rect 4441 -8723 4453 -8689
rect 4395 -8738 4453 -8723
rect 4653 -8553 4711 -8538
rect 4653 -8587 4665 -8553
rect 4699 -8587 4711 -8553
rect 4653 -8621 4711 -8587
rect 4653 -8655 4665 -8621
rect 4699 -8655 4711 -8621
rect 4653 -8689 4711 -8655
rect 4653 -8723 4665 -8689
rect 4699 -8723 4711 -8689
rect 4653 -8738 4711 -8723
rect 4847 -8553 4905 -8538
rect 4847 -8587 4859 -8553
rect 4893 -8587 4905 -8553
rect 4847 -8621 4905 -8587
rect 4847 -8655 4859 -8621
rect 4893 -8655 4905 -8621
rect 4847 -8689 4905 -8655
rect 4847 -8723 4859 -8689
rect 4893 -8723 4905 -8689
rect 4847 -8738 4905 -8723
rect 5105 -8553 5163 -8538
rect 5105 -8587 5117 -8553
rect 5151 -8587 5163 -8553
rect 5105 -8621 5163 -8587
rect 5105 -8655 5117 -8621
rect 5151 -8655 5163 -8621
rect 5105 -8689 5163 -8655
rect 5105 -8723 5117 -8689
rect 5151 -8723 5163 -8689
rect 5105 -8738 5163 -8723
rect 5333 -8553 5391 -8538
rect 5333 -8587 5345 -8553
rect 5379 -8587 5391 -8553
rect 5333 -8621 5391 -8587
rect 5333 -8655 5345 -8621
rect 5379 -8655 5391 -8621
rect 5333 -8689 5391 -8655
rect 5333 -8723 5345 -8689
rect 5379 -8723 5391 -8689
rect 5333 -8738 5391 -8723
rect 5591 -8553 5649 -8538
rect 5591 -8587 5603 -8553
rect 5637 -8587 5649 -8553
rect 5591 -8621 5649 -8587
rect 5591 -8655 5603 -8621
rect 5637 -8655 5649 -8621
rect 5591 -8689 5649 -8655
rect 5591 -8723 5603 -8689
rect 5637 -8723 5649 -8689
rect 5591 -8738 5649 -8723
rect 5784 -8553 5842 -8538
rect 5784 -8587 5796 -8553
rect 5830 -8587 5842 -8553
rect 5784 -8621 5842 -8587
rect 5784 -8655 5796 -8621
rect 5830 -8655 5842 -8621
rect 5784 -8689 5842 -8655
rect 5784 -8723 5796 -8689
rect 5830 -8723 5842 -8689
rect 5784 -8738 5842 -8723
rect 6042 -8553 6100 -8538
rect 6042 -8587 6054 -8553
rect 6088 -8587 6100 -8553
rect 6042 -8621 6100 -8587
rect 6042 -8655 6054 -8621
rect 6088 -8655 6100 -8621
rect 6042 -8689 6100 -8655
rect 6042 -8723 6054 -8689
rect 6088 -8723 6100 -8689
rect 6042 -8738 6100 -8723
rect 6300 -8553 6358 -8538
rect 6300 -8587 6312 -8553
rect 6346 -8587 6358 -8553
rect 6300 -8621 6358 -8587
rect 6300 -8655 6312 -8621
rect 6346 -8655 6358 -8621
rect 6300 -8689 6358 -8655
rect 6300 -8723 6312 -8689
rect 6346 -8723 6358 -8689
rect 6300 -8738 6358 -8723
rect 6558 -8553 6616 -8538
rect 6558 -8587 6570 -8553
rect 6604 -8587 6616 -8553
rect 6558 -8621 6616 -8587
rect 6558 -8655 6570 -8621
rect 6604 -8655 6616 -8621
rect 6558 -8689 6616 -8655
rect 6558 -8723 6570 -8689
rect 6604 -8723 6616 -8689
rect 6558 -8738 6616 -8723
rect 6816 -8553 6874 -8538
rect 6816 -8587 6828 -8553
rect 6862 -8587 6874 -8553
rect 6816 -8621 6874 -8587
rect 6816 -8655 6828 -8621
rect 6862 -8655 6874 -8621
rect 6816 -8689 6874 -8655
rect 6816 -8723 6828 -8689
rect 6862 -8723 6874 -8689
rect 6816 -8738 6874 -8723
rect 7010 -8553 7068 -8538
rect 7010 -8587 7022 -8553
rect 7056 -8587 7068 -8553
rect 7010 -8621 7068 -8587
rect 7010 -8655 7022 -8621
rect 7056 -8655 7068 -8621
rect 7010 -8689 7068 -8655
rect 7010 -8723 7022 -8689
rect 7056 -8723 7068 -8689
rect 7010 -8738 7068 -8723
rect 7268 -8553 7326 -8538
rect 7268 -8587 7280 -8553
rect 7314 -8587 7326 -8553
rect 7268 -8621 7326 -8587
rect 7268 -8655 7280 -8621
rect 7314 -8655 7326 -8621
rect 7268 -8689 7326 -8655
rect 7268 -8723 7280 -8689
rect 7314 -8723 7326 -8689
rect 7268 -8738 7326 -8723
rect 7526 -8553 7584 -8538
rect 7526 -8587 7538 -8553
rect 7572 -8587 7584 -8553
rect 7526 -8621 7584 -8587
rect 7526 -8655 7538 -8621
rect 7572 -8655 7584 -8621
rect 7526 -8689 7584 -8655
rect 7526 -8723 7538 -8689
rect 7572 -8723 7584 -8689
rect 7526 -8738 7584 -8723
rect 7784 -8553 7842 -8538
rect 7784 -8587 7796 -8553
rect 7830 -8587 7842 -8553
rect 7784 -8621 7842 -8587
rect 7784 -8655 7796 -8621
rect 7830 -8655 7842 -8621
rect 7784 -8689 7842 -8655
rect 7784 -8723 7796 -8689
rect 7830 -8723 7842 -8689
rect 7784 -8738 7842 -8723
rect 7978 -8553 8036 -8538
rect 7978 -8587 7990 -8553
rect 8024 -8587 8036 -8553
rect 7978 -8621 8036 -8587
rect 7978 -8655 7990 -8621
rect 8024 -8655 8036 -8621
rect 7978 -8689 8036 -8655
rect 7978 -8723 7990 -8689
rect 8024 -8723 8036 -8689
rect 7978 -8738 8036 -8723
rect 8236 -8553 8294 -8538
rect 8236 -8587 8248 -8553
rect 8282 -8587 8294 -8553
rect 8236 -8621 8294 -8587
rect 8236 -8655 8248 -8621
rect 8282 -8655 8294 -8621
rect 8236 -8689 8294 -8655
rect 8236 -8723 8248 -8689
rect 8282 -8723 8294 -8689
rect 8236 -8738 8294 -8723
rect 8494 -8553 8552 -8538
rect 8494 -8587 8506 -8553
rect 8540 -8587 8552 -8553
rect 8494 -8621 8552 -8587
rect 8494 -8655 8506 -8621
rect 8540 -8655 8552 -8621
rect 8494 -8689 8552 -8655
rect 8494 -8723 8506 -8689
rect 8540 -8723 8552 -8689
rect 8494 -8738 8552 -8723
rect 8752 -8553 8810 -8538
rect 8752 -8587 8764 -8553
rect 8798 -8587 8810 -8553
rect 8752 -8621 8810 -8587
rect 8752 -8655 8764 -8621
rect 8798 -8655 8810 -8621
rect 8752 -8689 8810 -8655
rect 8752 -8723 8764 -8689
rect 8798 -8723 8810 -8689
rect 8752 -8738 8810 -8723
rect 9010 -8553 9068 -8538
rect 9010 -8587 9022 -8553
rect 9056 -8587 9068 -8553
rect 9010 -8621 9068 -8587
rect 9010 -8655 9022 -8621
rect 9056 -8655 9068 -8621
rect 9010 -8689 9068 -8655
rect 9010 -8723 9022 -8689
rect 9056 -8723 9068 -8689
rect 9010 -8738 9068 -8723
rect 9204 -8553 9262 -8538
rect 9204 -8587 9216 -8553
rect 9250 -8587 9262 -8553
rect 9204 -8621 9262 -8587
rect 9204 -8655 9216 -8621
rect 9250 -8655 9262 -8621
rect 9204 -8689 9262 -8655
rect 9204 -8723 9216 -8689
rect 9250 -8723 9262 -8689
rect 9204 -8738 9262 -8723
rect 9462 -8553 9520 -8538
rect 9462 -8587 9474 -8553
rect 9508 -8587 9520 -8553
rect 9462 -8621 9520 -8587
rect 9462 -8655 9474 -8621
rect 9508 -8655 9520 -8621
rect 9462 -8689 9520 -8655
rect 9462 -8723 9474 -8689
rect 9508 -8723 9520 -8689
rect 9462 -8738 9520 -8723
<< pdiffc >>
rect 987 512 1021 546
rect 987 444 1021 478
rect 987 376 1021 410
rect 1245 512 1279 546
rect 1245 444 1279 478
rect 1245 376 1279 410
rect 1439 512 1473 546
rect 1439 444 1473 478
rect 1439 376 1473 410
rect 1697 512 1731 546
rect 1697 444 1731 478
rect 1697 376 1731 410
rect 1955 512 1989 546
rect 1955 444 1989 478
rect 1955 376 1989 410
rect 2213 512 2247 546
rect 2213 444 2247 478
rect 2213 376 2247 410
rect 2471 512 2505 546
rect 2471 444 2505 478
rect 2471 376 2505 410
rect 2665 512 2699 546
rect 2665 444 2699 478
rect 2665 376 2699 410
rect 2923 512 2957 546
rect 2923 444 2957 478
rect 2923 376 2957 410
rect 3181 512 3215 546
rect 3181 444 3215 478
rect 3181 376 3215 410
rect 3439 512 3473 546
rect 3439 444 3473 478
rect 3439 376 3473 410
rect 3633 512 3667 546
rect 3633 444 3667 478
rect 3633 376 3667 410
rect 3891 512 3925 546
rect 3891 444 3925 478
rect 3891 376 3925 410
rect 4149 512 4183 546
rect 4149 444 4183 478
rect 4149 376 4183 410
rect 4407 512 4441 546
rect 4407 444 4441 478
rect 4407 376 4441 410
rect 4665 512 4699 546
rect 4665 444 4699 478
rect 4665 376 4699 410
rect 4859 512 4893 546
rect 4859 444 4893 478
rect 4859 376 4893 410
rect 5117 512 5151 546
rect 5117 444 5151 478
rect 5117 376 5151 410
rect 5345 512 5379 546
rect 5345 444 5379 478
rect 5345 376 5379 410
rect 5603 512 5637 546
rect 5603 444 5637 478
rect 5603 376 5637 410
rect 5796 512 5830 546
rect 5796 444 5830 478
rect 5796 376 5830 410
rect 6054 512 6088 546
rect 6054 444 6088 478
rect 6054 376 6088 410
rect 6312 512 6346 546
rect 6312 444 6346 478
rect 6312 376 6346 410
rect 6570 512 6604 546
rect 6570 444 6604 478
rect 6570 376 6604 410
rect 6828 512 6862 546
rect 6828 444 6862 478
rect 6828 376 6862 410
rect 7022 512 7056 546
rect 7022 444 7056 478
rect 7022 376 7056 410
rect 7280 512 7314 546
rect 7280 444 7314 478
rect 7280 376 7314 410
rect 7538 512 7572 546
rect 7538 444 7572 478
rect 7538 376 7572 410
rect 7796 512 7830 546
rect 7796 444 7830 478
rect 7796 376 7830 410
rect 7990 512 8024 546
rect 7990 444 8024 478
rect 7990 376 8024 410
rect 8248 512 8282 546
rect 8248 444 8282 478
rect 8248 376 8282 410
rect 8506 512 8540 546
rect 8506 444 8540 478
rect 8506 376 8540 410
rect 8764 512 8798 546
rect 8764 444 8798 478
rect 8764 376 8798 410
rect 9022 512 9056 546
rect 9022 444 9056 478
rect 9022 376 9056 410
rect 9216 512 9250 546
rect 9216 444 9250 478
rect 9216 376 9250 410
rect 9474 512 9508 546
rect 9474 444 9508 478
rect 9474 376 9508 410
rect 987 -432 1021 -398
rect 987 -500 1021 -466
rect 987 -568 1021 -534
rect 1245 -432 1279 -398
rect 1245 -500 1279 -466
rect 1245 -568 1279 -534
rect 1439 -432 1473 -398
rect 1439 -500 1473 -466
rect 1439 -568 1473 -534
rect 1697 -432 1731 -398
rect 1697 -500 1731 -466
rect 1697 -568 1731 -534
rect 1955 -432 1989 -398
rect 1955 -500 1989 -466
rect 1955 -568 1989 -534
rect 2213 -432 2247 -398
rect 2213 -500 2247 -466
rect 2213 -568 2247 -534
rect 2471 -432 2505 -398
rect 2471 -500 2505 -466
rect 2471 -568 2505 -534
rect 2665 -432 2699 -398
rect 2665 -500 2699 -466
rect 2665 -568 2699 -534
rect 2923 -432 2957 -398
rect 2923 -500 2957 -466
rect 2923 -568 2957 -534
rect 3181 -432 3215 -398
rect 3181 -500 3215 -466
rect 3181 -568 3215 -534
rect 3439 -432 3473 -398
rect 3439 -500 3473 -466
rect 3439 -568 3473 -534
rect 3633 -432 3667 -398
rect 3633 -500 3667 -466
rect 3633 -568 3667 -534
rect 3891 -432 3925 -398
rect 3891 -500 3925 -466
rect 3891 -568 3925 -534
rect 4149 -432 4183 -398
rect 4149 -500 4183 -466
rect 4149 -568 4183 -534
rect 4407 -432 4441 -398
rect 4407 -500 4441 -466
rect 4407 -568 4441 -534
rect 4665 -432 4699 -398
rect 4665 -500 4699 -466
rect 4665 -568 4699 -534
rect 4859 -432 4893 -398
rect 4859 -500 4893 -466
rect 4859 -568 4893 -534
rect 5117 -432 5151 -398
rect 5117 -500 5151 -466
rect 5117 -568 5151 -534
rect 5345 -432 5379 -398
rect 5345 -500 5379 -466
rect 5345 -568 5379 -534
rect 5603 -432 5637 -398
rect 5603 -500 5637 -466
rect 5603 -568 5637 -534
rect 5796 -432 5830 -398
rect 5796 -500 5830 -466
rect 5796 -568 5830 -534
rect 6054 -432 6088 -398
rect 6054 -500 6088 -466
rect 6054 -568 6088 -534
rect 6312 -432 6346 -398
rect 6312 -500 6346 -466
rect 6312 -568 6346 -534
rect 6570 -432 6604 -398
rect 6570 -500 6604 -466
rect 6570 -568 6604 -534
rect 6828 -432 6862 -398
rect 6828 -500 6862 -466
rect 6828 -568 6862 -534
rect 7022 -432 7056 -398
rect 7022 -500 7056 -466
rect 7022 -568 7056 -534
rect 7280 -432 7314 -398
rect 7280 -500 7314 -466
rect 7280 -568 7314 -534
rect 7538 -432 7572 -398
rect 7538 -500 7572 -466
rect 7538 -568 7572 -534
rect 7796 -432 7830 -398
rect 7796 -500 7830 -466
rect 7796 -568 7830 -534
rect 7990 -432 8024 -398
rect 7990 -500 8024 -466
rect 7990 -568 8024 -534
rect 8248 -432 8282 -398
rect 8248 -500 8282 -466
rect 8248 -568 8282 -534
rect 8506 -432 8540 -398
rect 8506 -500 8540 -466
rect 8506 -568 8540 -534
rect 8764 -432 8798 -398
rect 8764 -500 8798 -466
rect 8764 -568 8798 -534
rect 9022 -432 9056 -398
rect 9022 -500 9056 -466
rect 9022 -568 9056 -534
rect 9216 -432 9250 -398
rect 9216 -500 9250 -466
rect 9216 -568 9250 -534
rect 9474 -432 9508 -398
rect 9474 -500 9508 -466
rect 9474 -568 9508 -534
rect 987 -1123 1021 -1089
rect 987 -1191 1021 -1157
rect 987 -1259 1021 -1225
rect 1245 -1123 1279 -1089
rect 1245 -1191 1279 -1157
rect 1245 -1259 1279 -1225
rect 1439 -1123 1473 -1089
rect 1439 -1191 1473 -1157
rect 1439 -1259 1473 -1225
rect 1697 -1123 1731 -1089
rect 1697 -1191 1731 -1157
rect 1697 -1259 1731 -1225
rect 1955 -1123 1989 -1089
rect 1955 -1191 1989 -1157
rect 1955 -1259 1989 -1225
rect 2213 -1123 2247 -1089
rect 2213 -1191 2247 -1157
rect 2213 -1259 2247 -1225
rect 2471 -1123 2505 -1089
rect 2471 -1191 2505 -1157
rect 2471 -1259 2505 -1225
rect 2665 -1123 2699 -1089
rect 2665 -1191 2699 -1157
rect 2665 -1259 2699 -1225
rect 2923 -1123 2957 -1089
rect 2923 -1191 2957 -1157
rect 2923 -1259 2957 -1225
rect 3181 -1123 3215 -1089
rect 3181 -1191 3215 -1157
rect 3181 -1259 3215 -1225
rect 3439 -1123 3473 -1089
rect 3439 -1191 3473 -1157
rect 3439 -1259 3473 -1225
rect 3633 -1123 3667 -1089
rect 3633 -1191 3667 -1157
rect 3633 -1259 3667 -1225
rect 3891 -1123 3925 -1089
rect 3891 -1191 3925 -1157
rect 3891 -1259 3925 -1225
rect 4149 -1123 4183 -1089
rect 4149 -1191 4183 -1157
rect 4149 -1259 4183 -1225
rect 4407 -1123 4441 -1089
rect 4407 -1191 4441 -1157
rect 4407 -1259 4441 -1225
rect 4665 -1123 4699 -1089
rect 4665 -1191 4699 -1157
rect 4665 -1259 4699 -1225
rect 4859 -1123 4893 -1089
rect 4859 -1191 4893 -1157
rect 4859 -1259 4893 -1225
rect 5117 -1123 5151 -1089
rect 5117 -1191 5151 -1157
rect 5117 -1259 5151 -1225
rect 5345 -1123 5379 -1089
rect 5345 -1191 5379 -1157
rect 5345 -1259 5379 -1225
rect 5603 -1123 5637 -1089
rect 5603 -1191 5637 -1157
rect 5603 -1259 5637 -1225
rect 5796 -1123 5830 -1089
rect 5796 -1191 5830 -1157
rect 5796 -1259 5830 -1225
rect 6054 -1123 6088 -1089
rect 6054 -1191 6088 -1157
rect 6054 -1259 6088 -1225
rect 6312 -1123 6346 -1089
rect 6312 -1191 6346 -1157
rect 6312 -1259 6346 -1225
rect 6570 -1123 6604 -1089
rect 6570 -1191 6604 -1157
rect 6570 -1259 6604 -1225
rect 6828 -1123 6862 -1089
rect 6828 -1191 6862 -1157
rect 6828 -1259 6862 -1225
rect 7022 -1123 7056 -1089
rect 7022 -1191 7056 -1157
rect 7022 -1259 7056 -1225
rect 7280 -1123 7314 -1089
rect 7280 -1191 7314 -1157
rect 7280 -1259 7314 -1225
rect 7538 -1123 7572 -1089
rect 7538 -1191 7572 -1157
rect 7538 -1259 7572 -1225
rect 7796 -1123 7830 -1089
rect 7796 -1191 7830 -1157
rect 7796 -1259 7830 -1225
rect 7990 -1123 8024 -1089
rect 7990 -1191 8024 -1157
rect 7990 -1259 8024 -1225
rect 8248 -1123 8282 -1089
rect 8248 -1191 8282 -1157
rect 8248 -1259 8282 -1225
rect 8506 -1123 8540 -1089
rect 8506 -1191 8540 -1157
rect 8506 -1259 8540 -1225
rect 8764 -1123 8798 -1089
rect 8764 -1191 8798 -1157
rect 8764 -1259 8798 -1225
rect 9022 -1123 9056 -1089
rect 9022 -1191 9056 -1157
rect 9022 -1259 9056 -1225
rect 9216 -1123 9250 -1089
rect 9216 -1191 9250 -1157
rect 9216 -1259 9250 -1225
rect 9474 -1123 9508 -1089
rect 9474 -1191 9508 -1157
rect 9474 -1259 9508 -1225
rect 987 -2079 1021 -2045
rect 987 -2147 1021 -2113
rect 987 -2215 1021 -2181
rect 1245 -2079 1279 -2045
rect 1245 -2147 1279 -2113
rect 1245 -2215 1279 -2181
rect 1439 -2079 1473 -2045
rect 1439 -2147 1473 -2113
rect 1439 -2215 1473 -2181
rect 1697 -2079 1731 -2045
rect 1697 -2147 1731 -2113
rect 1697 -2215 1731 -2181
rect 1955 -2079 1989 -2045
rect 1955 -2147 1989 -2113
rect 1955 -2215 1989 -2181
rect 2213 -2079 2247 -2045
rect 2213 -2147 2247 -2113
rect 2213 -2215 2247 -2181
rect 2471 -2079 2505 -2045
rect 2471 -2147 2505 -2113
rect 2471 -2215 2505 -2181
rect 2665 -2079 2699 -2045
rect 2665 -2147 2699 -2113
rect 2665 -2215 2699 -2181
rect 2923 -2079 2957 -2045
rect 2923 -2147 2957 -2113
rect 2923 -2215 2957 -2181
rect 3181 -2079 3215 -2045
rect 3181 -2147 3215 -2113
rect 3181 -2215 3215 -2181
rect 3439 -2079 3473 -2045
rect 3439 -2147 3473 -2113
rect 3439 -2215 3473 -2181
rect 3633 -2079 3667 -2045
rect 3633 -2147 3667 -2113
rect 3633 -2215 3667 -2181
rect 3891 -2079 3925 -2045
rect 3891 -2147 3925 -2113
rect 3891 -2215 3925 -2181
rect 4149 -2079 4183 -2045
rect 4149 -2147 4183 -2113
rect 4149 -2215 4183 -2181
rect 4407 -2079 4441 -2045
rect 4407 -2147 4441 -2113
rect 4407 -2215 4441 -2181
rect 4665 -2079 4699 -2045
rect 4665 -2147 4699 -2113
rect 4665 -2215 4699 -2181
rect 4859 -2079 4893 -2045
rect 4859 -2147 4893 -2113
rect 4859 -2215 4893 -2181
rect 5117 -2079 5151 -2045
rect 5117 -2147 5151 -2113
rect 5117 -2215 5151 -2181
rect 5345 -2079 5379 -2045
rect 5345 -2147 5379 -2113
rect 5345 -2215 5379 -2181
rect 5603 -2079 5637 -2045
rect 5603 -2147 5637 -2113
rect 5603 -2215 5637 -2181
rect 5796 -2079 5830 -2045
rect 5796 -2147 5830 -2113
rect 5796 -2215 5830 -2181
rect 6054 -2079 6088 -2045
rect 6054 -2147 6088 -2113
rect 6054 -2215 6088 -2181
rect 6312 -2079 6346 -2045
rect 6312 -2147 6346 -2113
rect 6312 -2215 6346 -2181
rect 6570 -2079 6604 -2045
rect 6570 -2147 6604 -2113
rect 6570 -2215 6604 -2181
rect 6828 -2079 6862 -2045
rect 6828 -2147 6862 -2113
rect 6828 -2215 6862 -2181
rect 7022 -2079 7056 -2045
rect 7022 -2147 7056 -2113
rect 7022 -2215 7056 -2181
rect 7280 -2079 7314 -2045
rect 7280 -2147 7314 -2113
rect 7280 -2215 7314 -2181
rect 7538 -2079 7572 -2045
rect 7538 -2147 7572 -2113
rect 7538 -2215 7572 -2181
rect 7796 -2079 7830 -2045
rect 7796 -2147 7830 -2113
rect 7796 -2215 7830 -2181
rect 7990 -2079 8024 -2045
rect 7990 -2147 8024 -2113
rect 7990 -2215 8024 -2181
rect 8248 -2079 8282 -2045
rect 8248 -2147 8282 -2113
rect 8248 -2215 8282 -2181
rect 8506 -2079 8540 -2045
rect 8506 -2147 8540 -2113
rect 8506 -2215 8540 -2181
rect 8764 -2079 8798 -2045
rect 8764 -2147 8798 -2113
rect 8764 -2215 8798 -2181
rect 9022 -2079 9056 -2045
rect 9022 -2147 9056 -2113
rect 9022 -2215 9056 -2181
rect 9216 -2079 9250 -2045
rect 9216 -2147 9250 -2113
rect 9216 -2215 9250 -2181
rect 9474 -2079 9508 -2045
rect 9474 -2147 9508 -2113
rect 9474 -2215 9508 -2181
rect 987 -2770 1021 -2736
rect 987 -2838 1021 -2804
rect 987 -2906 1021 -2872
rect 1245 -2770 1279 -2736
rect 1245 -2838 1279 -2804
rect 1245 -2906 1279 -2872
rect 1439 -2770 1473 -2736
rect 1439 -2838 1473 -2804
rect 1439 -2906 1473 -2872
rect 1697 -2770 1731 -2736
rect 1697 -2838 1731 -2804
rect 1697 -2906 1731 -2872
rect 1955 -2770 1989 -2736
rect 1955 -2838 1989 -2804
rect 1955 -2906 1989 -2872
rect 2213 -2770 2247 -2736
rect 2213 -2838 2247 -2804
rect 2213 -2906 2247 -2872
rect 2471 -2770 2505 -2736
rect 2471 -2838 2505 -2804
rect 2471 -2906 2505 -2872
rect 2665 -2770 2699 -2736
rect 2665 -2838 2699 -2804
rect 2665 -2906 2699 -2872
rect 2923 -2770 2957 -2736
rect 2923 -2838 2957 -2804
rect 2923 -2906 2957 -2872
rect 3181 -2770 3215 -2736
rect 3181 -2838 3215 -2804
rect 3181 -2906 3215 -2872
rect 3439 -2770 3473 -2736
rect 3439 -2838 3473 -2804
rect 3439 -2906 3473 -2872
rect 3633 -2770 3667 -2736
rect 3633 -2838 3667 -2804
rect 3633 -2906 3667 -2872
rect 3891 -2770 3925 -2736
rect 3891 -2838 3925 -2804
rect 3891 -2906 3925 -2872
rect 4149 -2770 4183 -2736
rect 4149 -2838 4183 -2804
rect 4149 -2906 4183 -2872
rect 4407 -2770 4441 -2736
rect 4407 -2838 4441 -2804
rect 4407 -2906 4441 -2872
rect 4665 -2770 4699 -2736
rect 4665 -2838 4699 -2804
rect 4665 -2906 4699 -2872
rect 4859 -2770 4893 -2736
rect 4859 -2838 4893 -2804
rect 4859 -2906 4893 -2872
rect 5117 -2770 5151 -2736
rect 5117 -2838 5151 -2804
rect 5117 -2906 5151 -2872
rect 5345 -2770 5379 -2736
rect 5345 -2838 5379 -2804
rect 5345 -2906 5379 -2872
rect 5603 -2770 5637 -2736
rect 5603 -2838 5637 -2804
rect 5603 -2906 5637 -2872
rect 5796 -2770 5830 -2736
rect 5796 -2838 5830 -2804
rect 5796 -2906 5830 -2872
rect 6054 -2770 6088 -2736
rect 6054 -2838 6088 -2804
rect 6054 -2906 6088 -2872
rect 6312 -2770 6346 -2736
rect 6312 -2838 6346 -2804
rect 6312 -2906 6346 -2872
rect 6570 -2770 6604 -2736
rect 6570 -2838 6604 -2804
rect 6570 -2906 6604 -2872
rect 6828 -2770 6862 -2736
rect 6828 -2838 6862 -2804
rect 6828 -2906 6862 -2872
rect 7022 -2770 7056 -2736
rect 7022 -2838 7056 -2804
rect 7022 -2906 7056 -2872
rect 7280 -2770 7314 -2736
rect 7280 -2838 7314 -2804
rect 7280 -2906 7314 -2872
rect 7538 -2770 7572 -2736
rect 7538 -2838 7572 -2804
rect 7538 -2906 7572 -2872
rect 7796 -2770 7830 -2736
rect 7796 -2838 7830 -2804
rect 7796 -2906 7830 -2872
rect 7990 -2770 8024 -2736
rect 7990 -2838 8024 -2804
rect 7990 -2906 8024 -2872
rect 8248 -2770 8282 -2736
rect 8248 -2838 8282 -2804
rect 8248 -2906 8282 -2872
rect 8506 -2770 8540 -2736
rect 8506 -2838 8540 -2804
rect 8506 -2906 8540 -2872
rect 8764 -2770 8798 -2736
rect 8764 -2838 8798 -2804
rect 8764 -2906 8798 -2872
rect 9022 -2770 9056 -2736
rect 9022 -2838 9056 -2804
rect 9022 -2906 9056 -2872
rect 9216 -2770 9250 -2736
rect 9216 -2838 9250 -2804
rect 9216 -2906 9250 -2872
rect 9474 -2770 9508 -2736
rect 9474 -2838 9508 -2804
rect 9474 -2906 9508 -2872
rect 987 -3760 1021 -3726
rect 987 -3828 1021 -3794
rect 987 -3896 1021 -3862
rect 1245 -3760 1279 -3726
rect 1245 -3828 1279 -3794
rect 1245 -3896 1279 -3862
rect 1439 -3760 1473 -3726
rect 1439 -3828 1473 -3794
rect 1439 -3896 1473 -3862
rect 1697 -3760 1731 -3726
rect 1697 -3828 1731 -3794
rect 1697 -3896 1731 -3862
rect 1955 -3760 1989 -3726
rect 1955 -3828 1989 -3794
rect 1955 -3896 1989 -3862
rect 2213 -3760 2247 -3726
rect 2213 -3828 2247 -3794
rect 2213 -3896 2247 -3862
rect 2471 -3760 2505 -3726
rect 2471 -3828 2505 -3794
rect 2471 -3896 2505 -3862
rect 2665 -3760 2699 -3726
rect 2665 -3828 2699 -3794
rect 2665 -3896 2699 -3862
rect 2923 -3760 2957 -3726
rect 2923 -3828 2957 -3794
rect 2923 -3896 2957 -3862
rect 3181 -3760 3215 -3726
rect 3181 -3828 3215 -3794
rect 3181 -3896 3215 -3862
rect 3439 -3760 3473 -3726
rect 3439 -3828 3473 -3794
rect 3439 -3896 3473 -3862
rect 3633 -3760 3667 -3726
rect 3633 -3828 3667 -3794
rect 3633 -3896 3667 -3862
rect 3891 -3760 3925 -3726
rect 3891 -3828 3925 -3794
rect 3891 -3896 3925 -3862
rect 4149 -3760 4183 -3726
rect 4149 -3828 4183 -3794
rect 4149 -3896 4183 -3862
rect 4407 -3760 4441 -3726
rect 4407 -3828 4441 -3794
rect 4407 -3896 4441 -3862
rect 4665 -3760 4699 -3726
rect 4665 -3828 4699 -3794
rect 4665 -3896 4699 -3862
rect 4859 -3760 4893 -3726
rect 4859 -3828 4893 -3794
rect 4859 -3896 4893 -3862
rect 5117 -3760 5151 -3726
rect 5117 -3828 5151 -3794
rect 5117 -3896 5151 -3862
rect 5345 -3760 5379 -3726
rect 5345 -3828 5379 -3794
rect 5345 -3896 5379 -3862
rect 5603 -3760 5637 -3726
rect 5603 -3828 5637 -3794
rect 5603 -3896 5637 -3862
rect 5796 -3760 5830 -3726
rect 5796 -3828 5830 -3794
rect 5796 -3896 5830 -3862
rect 6054 -3760 6088 -3726
rect 6054 -3828 6088 -3794
rect 6054 -3896 6088 -3862
rect 6312 -3760 6346 -3726
rect 6312 -3828 6346 -3794
rect 6312 -3896 6346 -3862
rect 6570 -3760 6604 -3726
rect 6570 -3828 6604 -3794
rect 6570 -3896 6604 -3862
rect 6828 -3760 6862 -3726
rect 6828 -3828 6862 -3794
rect 6828 -3896 6862 -3862
rect 7022 -3760 7056 -3726
rect 7022 -3828 7056 -3794
rect 7022 -3896 7056 -3862
rect 7280 -3760 7314 -3726
rect 7280 -3828 7314 -3794
rect 7280 -3896 7314 -3862
rect 7538 -3760 7572 -3726
rect 7538 -3828 7572 -3794
rect 7538 -3896 7572 -3862
rect 7796 -3760 7830 -3726
rect 7796 -3828 7830 -3794
rect 7796 -3896 7830 -3862
rect 7990 -3760 8024 -3726
rect 7990 -3828 8024 -3794
rect 7990 -3896 8024 -3862
rect 8248 -3760 8282 -3726
rect 8248 -3828 8282 -3794
rect 8248 -3896 8282 -3862
rect 8506 -3760 8540 -3726
rect 8506 -3828 8540 -3794
rect 8506 -3896 8540 -3862
rect 8764 -3760 8798 -3726
rect 8764 -3828 8798 -3794
rect 8764 -3896 8798 -3862
rect 9022 -3760 9056 -3726
rect 9022 -3828 9056 -3794
rect 9022 -3896 9056 -3862
rect 9216 -3760 9250 -3726
rect 9216 -3828 9250 -3794
rect 9216 -3896 9250 -3862
rect 9474 -3760 9508 -3726
rect 9474 -3828 9508 -3794
rect 9474 -3896 9508 -3862
rect 987 -4316 1021 -4282
rect 987 -4384 1021 -4350
rect 987 -4452 1021 -4418
rect 1245 -4316 1279 -4282
rect 1245 -4384 1279 -4350
rect 1245 -4452 1279 -4418
rect 1439 -4316 1473 -4282
rect 1439 -4384 1473 -4350
rect 1439 -4452 1473 -4418
rect 1697 -4316 1731 -4282
rect 1697 -4384 1731 -4350
rect 1697 -4452 1731 -4418
rect 1955 -4316 1989 -4282
rect 1955 -4384 1989 -4350
rect 1955 -4452 1989 -4418
rect 2213 -4316 2247 -4282
rect 2213 -4384 2247 -4350
rect 2213 -4452 2247 -4418
rect 2471 -4316 2505 -4282
rect 2471 -4384 2505 -4350
rect 2471 -4452 2505 -4418
rect 2665 -4316 2699 -4282
rect 2665 -4384 2699 -4350
rect 2665 -4452 2699 -4418
rect 2923 -4316 2957 -4282
rect 2923 -4384 2957 -4350
rect 2923 -4452 2957 -4418
rect 3181 -4316 3215 -4282
rect 3181 -4384 3215 -4350
rect 3181 -4452 3215 -4418
rect 3439 -4316 3473 -4282
rect 3439 -4384 3473 -4350
rect 3439 -4452 3473 -4418
rect 3633 -4316 3667 -4282
rect 3633 -4384 3667 -4350
rect 3633 -4452 3667 -4418
rect 3891 -4316 3925 -4282
rect 3891 -4384 3925 -4350
rect 3891 -4452 3925 -4418
rect 4149 -4316 4183 -4282
rect 4149 -4384 4183 -4350
rect 4149 -4452 4183 -4418
rect 4407 -4316 4441 -4282
rect 4407 -4384 4441 -4350
rect 4407 -4452 4441 -4418
rect 4665 -4316 4699 -4282
rect 4665 -4384 4699 -4350
rect 4665 -4452 4699 -4418
rect 4859 -4316 4893 -4282
rect 4859 -4384 4893 -4350
rect 4859 -4452 4893 -4418
rect 5117 -4316 5151 -4282
rect 5117 -4384 5151 -4350
rect 5117 -4452 5151 -4418
rect 5345 -4316 5379 -4282
rect 5345 -4384 5379 -4350
rect 5345 -4452 5379 -4418
rect 5603 -4316 5637 -4282
rect 5603 -4384 5637 -4350
rect 5603 -4452 5637 -4418
rect 5796 -4316 5830 -4282
rect 5796 -4384 5830 -4350
rect 5796 -4452 5830 -4418
rect 6054 -4316 6088 -4282
rect 6054 -4384 6088 -4350
rect 6054 -4452 6088 -4418
rect 6312 -4316 6346 -4282
rect 6312 -4384 6346 -4350
rect 6312 -4452 6346 -4418
rect 6570 -4316 6604 -4282
rect 6570 -4384 6604 -4350
rect 6570 -4452 6604 -4418
rect 6828 -4316 6862 -4282
rect 6828 -4384 6862 -4350
rect 6828 -4452 6862 -4418
rect 7022 -4316 7056 -4282
rect 7022 -4384 7056 -4350
rect 7022 -4452 7056 -4418
rect 7280 -4316 7314 -4282
rect 7280 -4384 7314 -4350
rect 7280 -4452 7314 -4418
rect 7538 -4316 7572 -4282
rect 7538 -4384 7572 -4350
rect 7538 -4452 7572 -4418
rect 7796 -4316 7830 -4282
rect 7796 -4384 7830 -4350
rect 7796 -4452 7830 -4418
rect 7990 -4316 8024 -4282
rect 7990 -4384 8024 -4350
rect 7990 -4452 8024 -4418
rect 8248 -4316 8282 -4282
rect 8248 -4384 8282 -4350
rect 8248 -4452 8282 -4418
rect 8506 -4316 8540 -4282
rect 8506 -4384 8540 -4350
rect 8506 -4452 8540 -4418
rect 8764 -4316 8798 -4282
rect 8764 -4384 8798 -4350
rect 8764 -4452 8798 -4418
rect 9022 -4316 9056 -4282
rect 9022 -4384 9056 -4350
rect 9022 -4452 9056 -4418
rect 9216 -4316 9250 -4282
rect 9216 -4384 9250 -4350
rect 9216 -4452 9250 -4418
rect 9474 -4316 9508 -4282
rect 9474 -4384 9508 -4350
rect 9474 -4452 9508 -4418
rect 987 -5306 1021 -5272
rect 987 -5374 1021 -5340
rect 987 -5442 1021 -5408
rect 1245 -5306 1279 -5272
rect 1245 -5374 1279 -5340
rect 1245 -5442 1279 -5408
rect 1439 -5306 1473 -5272
rect 1439 -5374 1473 -5340
rect 1439 -5442 1473 -5408
rect 1697 -5306 1731 -5272
rect 1697 -5374 1731 -5340
rect 1697 -5442 1731 -5408
rect 1955 -5306 1989 -5272
rect 1955 -5374 1989 -5340
rect 1955 -5442 1989 -5408
rect 2213 -5306 2247 -5272
rect 2213 -5374 2247 -5340
rect 2213 -5442 2247 -5408
rect 2471 -5306 2505 -5272
rect 2471 -5374 2505 -5340
rect 2471 -5442 2505 -5408
rect 2665 -5306 2699 -5272
rect 2665 -5374 2699 -5340
rect 2665 -5442 2699 -5408
rect 2923 -5306 2957 -5272
rect 2923 -5374 2957 -5340
rect 2923 -5442 2957 -5408
rect 3181 -5306 3215 -5272
rect 3181 -5374 3215 -5340
rect 3181 -5442 3215 -5408
rect 3439 -5306 3473 -5272
rect 3439 -5374 3473 -5340
rect 3439 -5442 3473 -5408
rect 3633 -5306 3667 -5272
rect 3633 -5374 3667 -5340
rect 3633 -5442 3667 -5408
rect 3891 -5306 3925 -5272
rect 3891 -5374 3925 -5340
rect 3891 -5442 3925 -5408
rect 4149 -5306 4183 -5272
rect 4149 -5374 4183 -5340
rect 4149 -5442 4183 -5408
rect 4407 -5306 4441 -5272
rect 4407 -5374 4441 -5340
rect 4407 -5442 4441 -5408
rect 4665 -5306 4699 -5272
rect 4665 -5374 4699 -5340
rect 4665 -5442 4699 -5408
rect 4859 -5306 4893 -5272
rect 4859 -5374 4893 -5340
rect 4859 -5442 4893 -5408
rect 5117 -5306 5151 -5272
rect 5117 -5374 5151 -5340
rect 5117 -5442 5151 -5408
rect 5345 -5306 5379 -5272
rect 5345 -5374 5379 -5340
rect 5345 -5442 5379 -5408
rect 5603 -5306 5637 -5272
rect 5603 -5374 5637 -5340
rect 5603 -5442 5637 -5408
rect 5796 -5306 5830 -5272
rect 5796 -5374 5830 -5340
rect 5796 -5442 5830 -5408
rect 6054 -5306 6088 -5272
rect 6054 -5374 6088 -5340
rect 6054 -5442 6088 -5408
rect 6312 -5306 6346 -5272
rect 6312 -5374 6346 -5340
rect 6312 -5442 6346 -5408
rect 6570 -5306 6604 -5272
rect 6570 -5374 6604 -5340
rect 6570 -5442 6604 -5408
rect 6828 -5306 6862 -5272
rect 6828 -5374 6862 -5340
rect 6828 -5442 6862 -5408
rect 7022 -5306 7056 -5272
rect 7022 -5374 7056 -5340
rect 7022 -5442 7056 -5408
rect 7280 -5306 7314 -5272
rect 7280 -5374 7314 -5340
rect 7280 -5442 7314 -5408
rect 7538 -5306 7572 -5272
rect 7538 -5374 7572 -5340
rect 7538 -5442 7572 -5408
rect 7796 -5306 7830 -5272
rect 7796 -5374 7830 -5340
rect 7796 -5442 7830 -5408
rect 7990 -5306 8024 -5272
rect 7990 -5374 8024 -5340
rect 7990 -5442 8024 -5408
rect 8248 -5306 8282 -5272
rect 8248 -5374 8282 -5340
rect 8248 -5442 8282 -5408
rect 8506 -5306 8540 -5272
rect 8506 -5374 8540 -5340
rect 8506 -5442 8540 -5408
rect 8764 -5306 8798 -5272
rect 8764 -5374 8798 -5340
rect 8764 -5442 8798 -5408
rect 9022 -5306 9056 -5272
rect 9022 -5374 9056 -5340
rect 9022 -5442 9056 -5408
rect 9216 -5306 9250 -5272
rect 9216 -5374 9250 -5340
rect 9216 -5442 9250 -5408
rect 9474 -5306 9508 -5272
rect 9474 -5374 9508 -5340
rect 9474 -5442 9508 -5408
rect 987 -5996 1021 -5962
rect 987 -6064 1021 -6030
rect 987 -6132 1021 -6098
rect 1245 -5996 1279 -5962
rect 1245 -6064 1279 -6030
rect 1245 -6132 1279 -6098
rect 1439 -5996 1473 -5962
rect 1439 -6064 1473 -6030
rect 1439 -6132 1473 -6098
rect 1697 -5996 1731 -5962
rect 1697 -6064 1731 -6030
rect 1697 -6132 1731 -6098
rect 1955 -5996 1989 -5962
rect 1955 -6064 1989 -6030
rect 1955 -6132 1989 -6098
rect 2213 -5996 2247 -5962
rect 2213 -6064 2247 -6030
rect 2213 -6132 2247 -6098
rect 2471 -5996 2505 -5962
rect 2471 -6064 2505 -6030
rect 2471 -6132 2505 -6098
rect 2665 -5996 2699 -5962
rect 2665 -6064 2699 -6030
rect 2665 -6132 2699 -6098
rect 2923 -5996 2957 -5962
rect 2923 -6064 2957 -6030
rect 2923 -6132 2957 -6098
rect 3181 -5996 3215 -5962
rect 3181 -6064 3215 -6030
rect 3181 -6132 3215 -6098
rect 3439 -5996 3473 -5962
rect 3439 -6064 3473 -6030
rect 3439 -6132 3473 -6098
rect 3633 -5996 3667 -5962
rect 3633 -6064 3667 -6030
rect 3633 -6132 3667 -6098
rect 3891 -5996 3925 -5962
rect 3891 -6064 3925 -6030
rect 3891 -6132 3925 -6098
rect 4149 -5996 4183 -5962
rect 4149 -6064 4183 -6030
rect 4149 -6132 4183 -6098
rect 4407 -5996 4441 -5962
rect 4407 -6064 4441 -6030
rect 4407 -6132 4441 -6098
rect 4665 -5996 4699 -5962
rect 4665 -6064 4699 -6030
rect 4665 -6132 4699 -6098
rect 4859 -5996 4893 -5962
rect 4859 -6064 4893 -6030
rect 4859 -6132 4893 -6098
rect 5117 -5996 5151 -5962
rect 5117 -6064 5151 -6030
rect 5117 -6132 5151 -6098
rect 5345 -5996 5379 -5962
rect 5345 -6064 5379 -6030
rect 5345 -6132 5379 -6098
rect 5603 -5996 5637 -5962
rect 5603 -6064 5637 -6030
rect 5603 -6132 5637 -6098
rect 5796 -5996 5830 -5962
rect 5796 -6064 5830 -6030
rect 5796 -6132 5830 -6098
rect 6054 -5996 6088 -5962
rect 6054 -6064 6088 -6030
rect 6054 -6132 6088 -6098
rect 6312 -5996 6346 -5962
rect 6312 -6064 6346 -6030
rect 6312 -6132 6346 -6098
rect 6570 -5996 6604 -5962
rect 6570 -6064 6604 -6030
rect 6570 -6132 6604 -6098
rect 6828 -5996 6862 -5962
rect 6828 -6064 6862 -6030
rect 6828 -6132 6862 -6098
rect 7022 -5996 7056 -5962
rect 7022 -6064 7056 -6030
rect 7022 -6132 7056 -6098
rect 7280 -5996 7314 -5962
rect 7280 -6064 7314 -6030
rect 7280 -6132 7314 -6098
rect 7538 -5996 7572 -5962
rect 7538 -6064 7572 -6030
rect 7538 -6132 7572 -6098
rect 7796 -5996 7830 -5962
rect 7796 -6064 7830 -6030
rect 7796 -6132 7830 -6098
rect 7990 -5996 8024 -5962
rect 7990 -6064 8024 -6030
rect 7990 -6132 8024 -6098
rect 8248 -5996 8282 -5962
rect 8248 -6064 8282 -6030
rect 8248 -6132 8282 -6098
rect 8506 -5996 8540 -5962
rect 8506 -6064 8540 -6030
rect 8506 -6132 8540 -6098
rect 8764 -5996 8798 -5962
rect 8764 -6064 8798 -6030
rect 8764 -6132 8798 -6098
rect 9022 -5996 9056 -5962
rect 9022 -6064 9056 -6030
rect 9022 -6132 9056 -6098
rect 9216 -5996 9250 -5962
rect 9216 -6064 9250 -6030
rect 9216 -6132 9250 -6098
rect 9474 -5996 9508 -5962
rect 9474 -6064 9508 -6030
rect 9474 -6132 9508 -6098
rect 987 -6953 1021 -6919
rect 987 -7021 1021 -6987
rect 987 -7089 1021 -7055
rect 1245 -6953 1279 -6919
rect 1245 -7021 1279 -6987
rect 1245 -7089 1279 -7055
rect 1439 -6953 1473 -6919
rect 1439 -7021 1473 -6987
rect 1439 -7089 1473 -7055
rect 1697 -6953 1731 -6919
rect 1697 -7021 1731 -6987
rect 1697 -7089 1731 -7055
rect 1955 -6953 1989 -6919
rect 1955 -7021 1989 -6987
rect 1955 -7089 1989 -7055
rect 2213 -6953 2247 -6919
rect 2213 -7021 2247 -6987
rect 2213 -7089 2247 -7055
rect 2471 -6953 2505 -6919
rect 2471 -7021 2505 -6987
rect 2471 -7089 2505 -7055
rect 2665 -6953 2699 -6919
rect 2665 -7021 2699 -6987
rect 2665 -7089 2699 -7055
rect 2923 -6953 2957 -6919
rect 2923 -7021 2957 -6987
rect 2923 -7089 2957 -7055
rect 3181 -6953 3215 -6919
rect 3181 -7021 3215 -6987
rect 3181 -7089 3215 -7055
rect 3439 -6953 3473 -6919
rect 3439 -7021 3473 -6987
rect 3439 -7089 3473 -7055
rect 3633 -6953 3667 -6919
rect 3633 -7021 3667 -6987
rect 3633 -7089 3667 -7055
rect 3891 -6953 3925 -6919
rect 3891 -7021 3925 -6987
rect 3891 -7089 3925 -7055
rect 4149 -6953 4183 -6919
rect 4149 -7021 4183 -6987
rect 4149 -7089 4183 -7055
rect 4407 -6953 4441 -6919
rect 4407 -7021 4441 -6987
rect 4407 -7089 4441 -7055
rect 4665 -6953 4699 -6919
rect 4665 -7021 4699 -6987
rect 4665 -7089 4699 -7055
rect 4859 -6953 4893 -6919
rect 4859 -7021 4893 -6987
rect 4859 -7089 4893 -7055
rect 5117 -6953 5151 -6919
rect 5117 -7021 5151 -6987
rect 5117 -7089 5151 -7055
rect 5345 -6953 5379 -6919
rect 5345 -7021 5379 -6987
rect 5345 -7089 5379 -7055
rect 5603 -6953 5637 -6919
rect 5603 -7021 5637 -6987
rect 5603 -7089 5637 -7055
rect 5796 -6953 5830 -6919
rect 5796 -7021 5830 -6987
rect 5796 -7089 5830 -7055
rect 6054 -6953 6088 -6919
rect 6054 -7021 6088 -6987
rect 6054 -7089 6088 -7055
rect 6312 -6953 6346 -6919
rect 6312 -7021 6346 -6987
rect 6312 -7089 6346 -7055
rect 6570 -6953 6604 -6919
rect 6570 -7021 6604 -6987
rect 6570 -7089 6604 -7055
rect 6828 -6953 6862 -6919
rect 6828 -7021 6862 -6987
rect 6828 -7089 6862 -7055
rect 7022 -6953 7056 -6919
rect 7022 -7021 7056 -6987
rect 7022 -7089 7056 -7055
rect 7280 -6953 7314 -6919
rect 7280 -7021 7314 -6987
rect 7280 -7089 7314 -7055
rect 7538 -6953 7572 -6919
rect 7538 -7021 7572 -6987
rect 7538 -7089 7572 -7055
rect 7796 -6953 7830 -6919
rect 7796 -7021 7830 -6987
rect 7796 -7089 7830 -7055
rect 7990 -6953 8024 -6919
rect 7990 -7021 8024 -6987
rect 7990 -7089 8024 -7055
rect 8248 -6953 8282 -6919
rect 8248 -7021 8282 -6987
rect 8248 -7089 8282 -7055
rect 8506 -6953 8540 -6919
rect 8506 -7021 8540 -6987
rect 8506 -7089 8540 -7055
rect 8764 -6953 8798 -6919
rect 8764 -7021 8798 -6987
rect 8764 -7089 8798 -7055
rect 9022 -6953 9056 -6919
rect 9022 -7021 9056 -6987
rect 9022 -7089 9056 -7055
rect 9216 -6953 9250 -6919
rect 9216 -7021 9250 -6987
rect 9216 -7089 9250 -7055
rect 9474 -6953 9508 -6919
rect 9474 -7021 9508 -6987
rect 9474 -7089 9508 -7055
rect 987 -7643 1021 -7609
rect 987 -7711 1021 -7677
rect 987 -7779 1021 -7745
rect 1245 -7643 1279 -7609
rect 1245 -7711 1279 -7677
rect 1245 -7779 1279 -7745
rect 1439 -7643 1473 -7609
rect 1439 -7711 1473 -7677
rect 1439 -7779 1473 -7745
rect 1697 -7643 1731 -7609
rect 1697 -7711 1731 -7677
rect 1697 -7779 1731 -7745
rect 1955 -7643 1989 -7609
rect 1955 -7711 1989 -7677
rect 1955 -7779 1989 -7745
rect 2213 -7643 2247 -7609
rect 2213 -7711 2247 -7677
rect 2213 -7779 2247 -7745
rect 2471 -7643 2505 -7609
rect 2471 -7711 2505 -7677
rect 2471 -7779 2505 -7745
rect 2665 -7643 2699 -7609
rect 2665 -7711 2699 -7677
rect 2665 -7779 2699 -7745
rect 2923 -7643 2957 -7609
rect 2923 -7711 2957 -7677
rect 2923 -7779 2957 -7745
rect 3181 -7643 3215 -7609
rect 3181 -7711 3215 -7677
rect 3181 -7779 3215 -7745
rect 3439 -7643 3473 -7609
rect 3439 -7711 3473 -7677
rect 3439 -7779 3473 -7745
rect 3633 -7643 3667 -7609
rect 3633 -7711 3667 -7677
rect 3633 -7779 3667 -7745
rect 3891 -7643 3925 -7609
rect 3891 -7711 3925 -7677
rect 3891 -7779 3925 -7745
rect 4149 -7643 4183 -7609
rect 4149 -7711 4183 -7677
rect 4149 -7779 4183 -7745
rect 4407 -7643 4441 -7609
rect 4407 -7711 4441 -7677
rect 4407 -7779 4441 -7745
rect 4665 -7643 4699 -7609
rect 4665 -7711 4699 -7677
rect 4665 -7779 4699 -7745
rect 4859 -7643 4893 -7609
rect 4859 -7711 4893 -7677
rect 4859 -7779 4893 -7745
rect 5117 -7643 5151 -7609
rect 5117 -7711 5151 -7677
rect 5117 -7779 5151 -7745
rect 5345 -7643 5379 -7609
rect 5345 -7711 5379 -7677
rect 5345 -7779 5379 -7745
rect 5603 -7643 5637 -7609
rect 5603 -7711 5637 -7677
rect 5603 -7779 5637 -7745
rect 5796 -7643 5830 -7609
rect 5796 -7711 5830 -7677
rect 5796 -7779 5830 -7745
rect 6054 -7643 6088 -7609
rect 6054 -7711 6088 -7677
rect 6054 -7779 6088 -7745
rect 6312 -7643 6346 -7609
rect 6312 -7711 6346 -7677
rect 6312 -7779 6346 -7745
rect 6570 -7643 6604 -7609
rect 6570 -7711 6604 -7677
rect 6570 -7779 6604 -7745
rect 6828 -7643 6862 -7609
rect 6828 -7711 6862 -7677
rect 6828 -7779 6862 -7745
rect 7022 -7643 7056 -7609
rect 7022 -7711 7056 -7677
rect 7022 -7779 7056 -7745
rect 7280 -7643 7314 -7609
rect 7280 -7711 7314 -7677
rect 7280 -7779 7314 -7745
rect 7538 -7643 7572 -7609
rect 7538 -7711 7572 -7677
rect 7538 -7779 7572 -7745
rect 7796 -7643 7830 -7609
rect 7796 -7711 7830 -7677
rect 7796 -7779 7830 -7745
rect 7990 -7643 8024 -7609
rect 7990 -7711 8024 -7677
rect 7990 -7779 8024 -7745
rect 8248 -7643 8282 -7609
rect 8248 -7711 8282 -7677
rect 8248 -7779 8282 -7745
rect 8506 -7643 8540 -7609
rect 8506 -7711 8540 -7677
rect 8506 -7779 8540 -7745
rect 8764 -7643 8798 -7609
rect 8764 -7711 8798 -7677
rect 8764 -7779 8798 -7745
rect 9022 -7643 9056 -7609
rect 9022 -7711 9056 -7677
rect 9022 -7779 9056 -7745
rect 9216 -7643 9250 -7609
rect 9216 -7711 9250 -7677
rect 9216 -7779 9250 -7745
rect 9474 -7643 9508 -7609
rect 9474 -7711 9508 -7677
rect 9474 -7779 9508 -7745
rect 987 -8587 1021 -8553
rect 987 -8655 1021 -8621
rect 987 -8723 1021 -8689
rect 1245 -8587 1279 -8553
rect 1245 -8655 1279 -8621
rect 1245 -8723 1279 -8689
rect 1439 -8587 1473 -8553
rect 1439 -8655 1473 -8621
rect 1439 -8723 1473 -8689
rect 1697 -8587 1731 -8553
rect 1697 -8655 1731 -8621
rect 1697 -8723 1731 -8689
rect 1955 -8587 1989 -8553
rect 1955 -8655 1989 -8621
rect 1955 -8723 1989 -8689
rect 2213 -8587 2247 -8553
rect 2213 -8655 2247 -8621
rect 2213 -8723 2247 -8689
rect 2471 -8587 2505 -8553
rect 2471 -8655 2505 -8621
rect 2471 -8723 2505 -8689
rect 2665 -8587 2699 -8553
rect 2665 -8655 2699 -8621
rect 2665 -8723 2699 -8689
rect 2923 -8587 2957 -8553
rect 2923 -8655 2957 -8621
rect 2923 -8723 2957 -8689
rect 3181 -8587 3215 -8553
rect 3181 -8655 3215 -8621
rect 3181 -8723 3215 -8689
rect 3439 -8587 3473 -8553
rect 3439 -8655 3473 -8621
rect 3439 -8723 3473 -8689
rect 3633 -8587 3667 -8553
rect 3633 -8655 3667 -8621
rect 3633 -8723 3667 -8689
rect 3891 -8587 3925 -8553
rect 3891 -8655 3925 -8621
rect 3891 -8723 3925 -8689
rect 4149 -8587 4183 -8553
rect 4149 -8655 4183 -8621
rect 4149 -8723 4183 -8689
rect 4407 -8587 4441 -8553
rect 4407 -8655 4441 -8621
rect 4407 -8723 4441 -8689
rect 4665 -8587 4699 -8553
rect 4665 -8655 4699 -8621
rect 4665 -8723 4699 -8689
rect 4859 -8587 4893 -8553
rect 4859 -8655 4893 -8621
rect 4859 -8723 4893 -8689
rect 5117 -8587 5151 -8553
rect 5117 -8655 5151 -8621
rect 5117 -8723 5151 -8689
rect 5345 -8587 5379 -8553
rect 5345 -8655 5379 -8621
rect 5345 -8723 5379 -8689
rect 5603 -8587 5637 -8553
rect 5603 -8655 5637 -8621
rect 5603 -8723 5637 -8689
rect 5796 -8587 5830 -8553
rect 5796 -8655 5830 -8621
rect 5796 -8723 5830 -8689
rect 6054 -8587 6088 -8553
rect 6054 -8655 6088 -8621
rect 6054 -8723 6088 -8689
rect 6312 -8587 6346 -8553
rect 6312 -8655 6346 -8621
rect 6312 -8723 6346 -8689
rect 6570 -8587 6604 -8553
rect 6570 -8655 6604 -8621
rect 6570 -8723 6604 -8689
rect 6828 -8587 6862 -8553
rect 6828 -8655 6862 -8621
rect 6828 -8723 6862 -8689
rect 7022 -8587 7056 -8553
rect 7022 -8655 7056 -8621
rect 7022 -8723 7056 -8689
rect 7280 -8587 7314 -8553
rect 7280 -8655 7314 -8621
rect 7280 -8723 7314 -8689
rect 7538 -8587 7572 -8553
rect 7538 -8655 7572 -8621
rect 7538 -8723 7572 -8689
rect 7796 -8587 7830 -8553
rect 7796 -8655 7830 -8621
rect 7796 -8723 7830 -8689
rect 7990 -8587 8024 -8553
rect 7990 -8655 8024 -8621
rect 7990 -8723 8024 -8689
rect 8248 -8587 8282 -8553
rect 8248 -8655 8282 -8621
rect 8248 -8723 8282 -8689
rect 8506 -8587 8540 -8553
rect 8506 -8655 8540 -8621
rect 8506 -8723 8540 -8689
rect 8764 -8587 8798 -8553
rect 8764 -8655 8798 -8621
rect 8764 -8723 8798 -8689
rect 9022 -8587 9056 -8553
rect 9022 -8655 9056 -8621
rect 9022 -8723 9056 -8689
rect 9216 -8587 9250 -8553
rect 9216 -8655 9250 -8621
rect 9216 -8723 9250 -8689
rect 9474 -8587 9508 -8553
rect 9474 -8655 9508 -8621
rect 9474 -8723 9508 -8689
<< nsubdiff >>
rect 872 722 993 756
rect 1027 722 1061 756
rect 1095 722 1129 756
rect 1163 722 1197 756
rect 1231 722 1265 756
rect 1299 722 1333 756
rect 1367 722 1401 756
rect 1435 722 1469 756
rect 1503 722 1537 756
rect 1571 722 1605 756
rect 1639 722 1673 756
rect 1707 722 1741 756
rect 1775 722 1809 756
rect 1843 722 1877 756
rect 1911 722 1945 756
rect 1979 722 2013 756
rect 2047 722 2081 756
rect 2115 722 2149 756
rect 2183 722 2217 756
rect 2251 722 2285 756
rect 2319 722 2353 756
rect 2387 722 2421 756
rect 2455 722 2489 756
rect 2523 722 2557 756
rect 2591 722 2625 756
rect 2659 722 2693 756
rect 2727 722 2761 756
rect 2795 722 2829 756
rect 2863 722 2897 756
rect 2931 722 2965 756
rect 2999 722 3033 756
rect 3067 722 3101 756
rect 3135 722 3169 756
rect 3203 722 3237 756
rect 3271 722 3305 756
rect 3339 722 3373 756
rect 3407 722 3441 756
rect 3475 722 3509 756
rect 3543 722 3577 756
rect 3611 722 3645 756
rect 3679 722 3713 756
rect 3747 722 3781 756
rect 3815 722 3849 756
rect 3883 722 3917 756
rect 3951 722 3985 756
rect 4019 722 4053 756
rect 4087 722 4121 756
rect 4155 722 4189 756
rect 4223 722 4257 756
rect 4291 722 4325 756
rect 4359 722 4393 756
rect 4427 722 4461 756
rect 4495 722 4529 756
rect 4563 722 4597 756
rect 4631 722 4665 756
rect 4699 722 4733 756
rect 4767 722 4801 756
rect 4835 722 4869 756
rect 4903 722 4937 756
rect 4971 722 5005 756
rect 5039 722 5073 756
rect 5107 722 5388 756
rect 5422 722 5456 756
rect 5490 722 5524 756
rect 5558 722 5592 756
rect 5626 722 5660 756
rect 5694 722 5728 756
rect 5762 722 5796 756
rect 5830 722 5864 756
rect 5898 722 5932 756
rect 5966 722 6000 756
rect 6034 722 6068 756
rect 6102 722 6136 756
rect 6170 722 6204 756
rect 6238 722 6272 756
rect 6306 722 6340 756
rect 6374 722 6408 756
rect 6442 722 6476 756
rect 6510 722 6544 756
rect 6578 722 6612 756
rect 6646 722 6680 756
rect 6714 722 6748 756
rect 6782 722 6816 756
rect 6850 722 6884 756
rect 6918 722 6952 756
rect 6986 722 7020 756
rect 7054 722 7088 756
rect 7122 722 7156 756
rect 7190 722 7224 756
rect 7258 722 7292 756
rect 7326 722 7360 756
rect 7394 722 7428 756
rect 7462 722 7496 756
rect 7530 722 7564 756
rect 7598 722 7632 756
rect 7666 722 7700 756
rect 7734 722 7768 756
rect 7802 722 7836 756
rect 7870 722 7904 756
rect 7938 722 7972 756
rect 8006 722 8040 756
rect 8074 722 8108 756
rect 8142 722 8176 756
rect 8210 722 8244 756
rect 8278 722 8312 756
rect 8346 722 8380 756
rect 8414 722 8448 756
rect 8482 722 8516 756
rect 8550 722 8584 756
rect 8618 722 8652 756
rect 8686 722 8720 756
rect 8754 722 8788 756
rect 8822 722 8856 756
rect 8890 722 8924 756
rect 8958 722 8992 756
rect 9026 722 9060 756
rect 9094 722 9128 756
rect 9162 722 9196 756
rect 9230 722 9264 756
rect 9298 722 9332 756
rect 9366 722 9400 756
rect 9434 722 9468 756
rect 9502 722 9623 756
rect 872 543 906 722
rect 872 475 906 509
rect 872 407 906 441
rect 872 339 906 373
rect 5231 543 5265 722
rect 5231 475 5265 509
rect 5231 407 5265 441
rect 5231 339 5265 373
rect 9589 543 9623 722
rect 9589 475 9623 509
rect 9589 407 9623 441
rect 872 271 906 305
rect 872 203 906 237
rect 872 135 906 169
rect 872 67 906 101
rect 872 -1 906 33
rect 9589 339 9623 373
rect 5231 271 5265 305
rect 5231 203 5265 237
rect 5231 135 5265 169
rect 5231 67 5265 101
rect 5231 -1 5265 33
rect 9589 271 9623 305
rect 9589 203 9623 237
rect 9589 135 9623 169
rect 9589 67 9623 101
rect 9589 -1 9623 33
rect 872 -69 993 -35
rect 1027 -69 1061 -35
rect 1095 -69 1129 -35
rect 1163 -69 1197 -35
rect 1231 -69 1265 -35
rect 1299 -69 1333 -35
rect 1367 -69 1401 -35
rect 1435 -69 1469 -35
rect 1503 -69 1537 -35
rect 1571 -69 1605 -35
rect 1639 -69 1673 -35
rect 1707 -69 1741 -35
rect 1775 -69 1809 -35
rect 1843 -69 1877 -35
rect 1911 -69 1945 -35
rect 1979 -69 2013 -35
rect 2047 -69 2081 -35
rect 2115 -69 2149 -35
rect 2183 -69 2217 -35
rect 2251 -69 2285 -35
rect 2319 -69 2353 -35
rect 2387 -69 2421 -35
rect 2455 -69 2489 -35
rect 2523 -69 2557 -35
rect 2591 -69 2625 -35
rect 2659 -69 2693 -35
rect 2727 -69 2761 -35
rect 2795 -69 2829 -35
rect 2863 -69 2897 -35
rect 2931 -69 2965 -35
rect 2999 -69 3033 -35
rect 3067 -69 3101 -35
rect 3135 -69 3169 -35
rect 3203 -69 3237 -35
rect 3271 -69 3305 -35
rect 3339 -69 3373 -35
rect 3407 -69 3441 -35
rect 3475 -69 3509 -35
rect 3543 -69 3577 -35
rect 3611 -69 3645 -35
rect 3679 -69 3713 -35
rect 3747 -69 3781 -35
rect 3815 -69 3849 -35
rect 3883 -69 3917 -35
rect 3951 -69 3985 -35
rect 4019 -69 4053 -35
rect 4087 -69 4121 -35
rect 4155 -69 4189 -35
rect 4223 -69 4257 -35
rect 4291 -69 4325 -35
rect 4359 -69 4393 -35
rect 4427 -69 4461 -35
rect 4495 -69 4529 -35
rect 4563 -69 4597 -35
rect 4631 -69 4665 -35
rect 4699 -69 4733 -35
rect 4767 -69 4801 -35
rect 4835 -69 4869 -35
rect 4903 -69 4937 -35
rect 4971 -69 5005 -35
rect 5039 -69 5073 -35
rect 5107 -69 5388 -35
rect 5422 -69 5456 -35
rect 5490 -69 5524 -35
rect 5558 -69 5592 -35
rect 5626 -69 5660 -35
rect 5694 -69 5728 -35
rect 5762 -69 5796 -35
rect 5830 -69 5864 -35
rect 5898 -69 5932 -35
rect 5966 -69 6000 -35
rect 6034 -69 6068 -35
rect 6102 -69 6136 -35
rect 6170 -69 6204 -35
rect 6238 -69 6272 -35
rect 6306 -69 6340 -35
rect 6374 -69 6408 -35
rect 6442 -69 6476 -35
rect 6510 -69 6544 -35
rect 6578 -69 6612 -35
rect 6646 -69 6680 -35
rect 6714 -69 6748 -35
rect 6782 -69 6816 -35
rect 6850 -69 6884 -35
rect 6918 -69 6952 -35
rect 6986 -69 7020 -35
rect 7054 -69 7088 -35
rect 7122 -69 7156 -35
rect 7190 -69 7224 -35
rect 7258 -69 7292 -35
rect 7326 -69 7360 -35
rect 7394 -69 7428 -35
rect 7462 -69 7496 -35
rect 7530 -69 7564 -35
rect 7598 -69 7632 -35
rect 7666 -69 7700 -35
rect 7734 -69 7768 -35
rect 7802 -69 7836 -35
rect 7870 -69 7904 -35
rect 7938 -69 7972 -35
rect 8006 -69 8040 -35
rect 8074 -69 8108 -35
rect 8142 -69 8176 -35
rect 8210 -69 8244 -35
rect 8278 -69 8312 -35
rect 8346 -69 8380 -35
rect 8414 -69 8448 -35
rect 8482 -69 8516 -35
rect 8550 -69 8584 -35
rect 8618 -69 8652 -35
rect 8686 -69 8720 -35
rect 8754 -69 8788 -35
rect 8822 -69 8856 -35
rect 8890 -69 8924 -35
rect 8958 -69 8992 -35
rect 9026 -69 9060 -35
rect 9094 -69 9128 -35
rect 9162 -69 9196 -35
rect 9230 -69 9264 -35
rect 9298 -69 9332 -35
rect 9366 -69 9400 -35
rect 9434 -69 9468 -35
rect 9502 -69 9623 -35
rect 872 -137 906 -103
rect 872 -205 906 -171
rect 872 -273 906 -239
rect 872 -341 906 -307
rect 5231 -137 5265 -103
rect 5231 -205 5265 -171
rect 5231 -273 5265 -239
rect 5231 -341 5265 -307
rect 872 -409 906 -375
rect 9589 -137 9623 -103
rect 9589 -205 9623 -171
rect 9589 -273 9623 -239
rect 9589 -341 9623 -307
rect 872 -477 906 -443
rect 872 -545 906 -511
rect 872 -613 906 -579
rect 5231 -409 5265 -375
rect 5231 -477 5265 -443
rect 5231 -545 5265 -511
rect 872 -681 906 -647
rect 5231 -613 5265 -579
rect 9589 -409 9623 -375
rect 9589 -477 9623 -443
rect 9589 -545 9623 -511
rect 872 -749 906 -715
rect 872 -817 906 -783
rect 872 -885 906 -851
rect 872 -953 906 -919
rect 5231 -681 5265 -647
rect 9589 -613 9623 -579
rect 5231 -749 5265 -715
rect 5231 -817 5265 -783
rect 5231 -885 5265 -851
rect 5231 -953 5265 -919
rect 872 -1021 906 -987
rect 872 -1089 906 -1055
rect 9589 -681 9623 -647
rect 9589 -749 9623 -715
rect 9589 -817 9623 -783
rect 9589 -885 9623 -851
rect 9589 -953 9623 -919
rect 5231 -1021 5265 -987
rect 872 -1157 906 -1123
rect 872 -1225 906 -1191
rect 872 -1293 906 -1259
rect 5231 -1089 5265 -1055
rect 9589 -1021 9623 -987
rect 5231 -1157 5265 -1123
rect 5231 -1225 5265 -1191
rect 5231 -1293 5265 -1259
rect 9589 -1089 9623 -1055
rect 9589 -1157 9623 -1123
rect 9589 -1225 9623 -1191
rect 872 -1361 906 -1327
rect 872 -1429 906 -1395
rect 872 -1497 906 -1463
rect 872 -1633 906 -1531
rect 9589 -1293 9623 -1259
rect 5231 -1361 5265 -1327
rect 5231 -1429 5265 -1395
rect 5231 -1497 5265 -1463
rect 5231 -1633 5265 -1531
rect 9589 -1361 9623 -1327
rect 9589 -1429 9623 -1395
rect 9589 -1497 9623 -1463
rect 9589 -1633 9623 -1531
rect 872 -1667 993 -1633
rect 1027 -1667 1061 -1633
rect 1095 -1667 1129 -1633
rect 1163 -1667 1197 -1633
rect 1231 -1667 1265 -1633
rect 1299 -1667 1333 -1633
rect 1367 -1667 1401 -1633
rect 1435 -1667 1469 -1633
rect 1503 -1667 1537 -1633
rect 1571 -1667 1605 -1633
rect 1639 -1667 1673 -1633
rect 1707 -1667 1741 -1633
rect 1775 -1667 1809 -1633
rect 1843 -1667 1877 -1633
rect 1911 -1667 1945 -1633
rect 1979 -1667 2013 -1633
rect 2047 -1667 2081 -1633
rect 2115 -1667 2149 -1633
rect 2183 -1667 2217 -1633
rect 2251 -1667 2285 -1633
rect 2319 -1667 2353 -1633
rect 2387 -1667 2421 -1633
rect 2455 -1667 2489 -1633
rect 2523 -1667 2557 -1633
rect 2591 -1667 2625 -1633
rect 2659 -1667 2693 -1633
rect 2727 -1667 2761 -1633
rect 2795 -1667 2829 -1633
rect 2863 -1667 2897 -1633
rect 2931 -1667 2965 -1633
rect 2999 -1667 3033 -1633
rect 3067 -1667 3101 -1633
rect 3135 -1667 3169 -1633
rect 3203 -1667 3237 -1633
rect 3271 -1667 3305 -1633
rect 3339 -1667 3373 -1633
rect 3407 -1667 3441 -1633
rect 3475 -1667 3509 -1633
rect 3543 -1667 3577 -1633
rect 3611 -1667 3645 -1633
rect 3679 -1667 3713 -1633
rect 3747 -1667 3781 -1633
rect 3815 -1667 3849 -1633
rect 3883 -1667 3917 -1633
rect 3951 -1667 3985 -1633
rect 4019 -1667 4053 -1633
rect 4087 -1667 4121 -1633
rect 4155 -1667 4189 -1633
rect 4223 -1667 4257 -1633
rect 4291 -1667 4325 -1633
rect 4359 -1667 4393 -1633
rect 4427 -1667 4461 -1633
rect 4495 -1667 4529 -1633
rect 4563 -1667 4597 -1633
rect 4631 -1667 4665 -1633
rect 4699 -1667 4733 -1633
rect 4767 -1667 4801 -1633
rect 4835 -1667 4869 -1633
rect 4903 -1667 4937 -1633
rect 4971 -1667 5005 -1633
rect 5039 -1667 5073 -1633
rect 5107 -1667 5388 -1633
rect 5422 -1667 5456 -1633
rect 5490 -1667 5524 -1633
rect 5558 -1667 5592 -1633
rect 5626 -1667 5660 -1633
rect 5694 -1667 5728 -1633
rect 5762 -1667 5796 -1633
rect 5830 -1667 5864 -1633
rect 5898 -1667 5932 -1633
rect 5966 -1667 6000 -1633
rect 6034 -1667 6068 -1633
rect 6102 -1667 6136 -1633
rect 6170 -1667 6204 -1633
rect 6238 -1667 6272 -1633
rect 6306 -1667 6340 -1633
rect 6374 -1667 6408 -1633
rect 6442 -1667 6476 -1633
rect 6510 -1667 6544 -1633
rect 6578 -1667 6612 -1633
rect 6646 -1667 6680 -1633
rect 6714 -1667 6748 -1633
rect 6782 -1667 6816 -1633
rect 6850 -1667 6884 -1633
rect 6918 -1667 6952 -1633
rect 6986 -1667 7020 -1633
rect 7054 -1667 7088 -1633
rect 7122 -1667 7156 -1633
rect 7190 -1667 7224 -1633
rect 7258 -1667 7292 -1633
rect 7326 -1667 7360 -1633
rect 7394 -1667 7428 -1633
rect 7462 -1667 7496 -1633
rect 7530 -1667 7564 -1633
rect 7598 -1667 7632 -1633
rect 7666 -1667 7700 -1633
rect 7734 -1667 7768 -1633
rect 7802 -1667 7836 -1633
rect 7870 -1667 7904 -1633
rect 7938 -1667 7972 -1633
rect 8006 -1667 8040 -1633
rect 8074 -1667 8108 -1633
rect 8142 -1667 8176 -1633
rect 8210 -1667 8244 -1633
rect 8278 -1667 8312 -1633
rect 8346 -1667 8380 -1633
rect 8414 -1667 8448 -1633
rect 8482 -1667 8516 -1633
rect 8550 -1667 8584 -1633
rect 8618 -1667 8652 -1633
rect 8686 -1667 8720 -1633
rect 8754 -1667 8788 -1633
rect 8822 -1667 8856 -1633
rect 8890 -1667 8924 -1633
rect 8958 -1667 8992 -1633
rect 9026 -1667 9060 -1633
rect 9094 -1667 9128 -1633
rect 9162 -1667 9196 -1633
rect 9230 -1667 9264 -1633
rect 9298 -1667 9332 -1633
rect 9366 -1667 9400 -1633
rect 9434 -1667 9468 -1633
rect 9502 -1667 9623 -1633
rect 872 -1769 906 -1667
rect 872 -1837 906 -1803
rect 872 -1905 906 -1871
rect 872 -1973 906 -1939
rect 5231 -1769 5265 -1667
rect 5231 -1837 5265 -1803
rect 5231 -1905 5265 -1871
rect 5231 -1973 5265 -1939
rect 872 -2041 906 -2007
rect 9589 -1769 9623 -1667
rect 9589 -1837 9623 -1803
rect 9589 -1905 9623 -1871
rect 9589 -1973 9623 -1939
rect 872 -2109 906 -2075
rect 872 -2177 906 -2143
rect 872 -2245 906 -2211
rect 5231 -2041 5265 -2007
rect 5231 -2109 5265 -2075
rect 5231 -2177 5265 -2143
rect 872 -2313 906 -2279
rect 5231 -2245 5265 -2211
rect 9589 -2041 9623 -2007
rect 9589 -2109 9623 -2075
rect 9589 -2177 9623 -2143
rect 5231 -2313 5265 -2279
rect 872 -2381 906 -2347
rect 872 -2449 906 -2415
rect 872 -2517 906 -2483
rect 872 -2585 906 -2551
rect 872 -2653 906 -2619
rect 9589 -2245 9623 -2211
rect 9589 -2313 9623 -2279
rect 5231 -2381 5265 -2347
rect 5231 -2449 5265 -2415
rect 5231 -2517 5265 -2483
rect 5231 -2585 5265 -2551
rect 872 -2721 906 -2687
rect 5231 -2653 5265 -2619
rect 9589 -2381 9623 -2347
rect 9589 -2449 9623 -2415
rect 9589 -2517 9623 -2483
rect 9589 -2585 9623 -2551
rect 5231 -2721 5265 -2687
rect 9589 -2653 9623 -2619
rect 9589 -2721 9623 -2687
rect 872 -2789 906 -2755
rect 872 -2857 906 -2823
rect 872 -2925 906 -2891
rect 5231 -2789 5265 -2755
rect 5231 -2857 5265 -2823
rect 5231 -2925 5265 -2891
rect 9589 -2789 9623 -2755
rect 9589 -2857 9623 -2823
rect 872 -2993 906 -2959
rect 872 -3061 906 -3027
rect 872 -3129 906 -3095
rect 872 -3197 906 -3163
rect 872 -3265 906 -3231
rect 9589 -2925 9623 -2891
rect 5231 -2993 5265 -2959
rect 5231 -3061 5265 -3027
rect 5231 -3129 5265 -3095
rect 5231 -3197 5265 -3163
rect 5231 -3265 5265 -3231
rect 9589 -2993 9623 -2959
rect 9589 -3061 9623 -3027
rect 9589 -3129 9623 -3095
rect 9589 -3197 9623 -3163
rect 9589 -3265 9623 -3231
rect 872 -3333 993 -3299
rect 1027 -3333 1061 -3299
rect 1095 -3333 1129 -3299
rect 1163 -3333 1197 -3299
rect 1231 -3333 1265 -3299
rect 1299 -3333 1333 -3299
rect 1367 -3333 1401 -3299
rect 1435 -3333 1469 -3299
rect 1503 -3333 1537 -3299
rect 1571 -3333 1605 -3299
rect 1639 -3333 1673 -3299
rect 1707 -3333 1741 -3299
rect 1775 -3333 1809 -3299
rect 1843 -3333 1877 -3299
rect 1911 -3333 1945 -3299
rect 1979 -3333 2013 -3299
rect 2047 -3333 2081 -3299
rect 2115 -3333 2149 -3299
rect 2183 -3333 2217 -3299
rect 2251 -3333 2285 -3299
rect 2319 -3333 2353 -3299
rect 2387 -3333 2421 -3299
rect 2455 -3333 2489 -3299
rect 2523 -3333 2557 -3299
rect 2591 -3333 2625 -3299
rect 2659 -3333 2693 -3299
rect 2727 -3333 2761 -3299
rect 2795 -3333 2829 -3299
rect 2863 -3333 2897 -3299
rect 2931 -3333 2965 -3299
rect 2999 -3333 3033 -3299
rect 3067 -3333 3101 -3299
rect 3135 -3333 3169 -3299
rect 3203 -3333 3237 -3299
rect 3271 -3333 3305 -3299
rect 3339 -3333 3373 -3299
rect 3407 -3333 3441 -3299
rect 3475 -3333 3509 -3299
rect 3543 -3333 3577 -3299
rect 3611 -3333 3645 -3299
rect 3679 -3333 3713 -3299
rect 3747 -3333 3781 -3299
rect 3815 -3333 3849 -3299
rect 3883 -3333 3917 -3299
rect 3951 -3333 3985 -3299
rect 4019 -3333 4053 -3299
rect 4087 -3333 4121 -3299
rect 4155 -3333 4189 -3299
rect 4223 -3333 4257 -3299
rect 4291 -3333 4325 -3299
rect 4359 -3333 4393 -3299
rect 4427 -3333 4461 -3299
rect 4495 -3333 4529 -3299
rect 4563 -3333 4597 -3299
rect 4631 -3333 4665 -3299
rect 4699 -3333 4733 -3299
rect 4767 -3333 4801 -3299
rect 4835 -3333 4869 -3299
rect 4903 -3333 4937 -3299
rect 4971 -3333 5005 -3299
rect 5039 -3333 5073 -3299
rect 5107 -3333 5388 -3299
rect 5422 -3333 5456 -3299
rect 5490 -3333 5524 -3299
rect 5558 -3333 5592 -3299
rect 5626 -3333 5660 -3299
rect 5694 -3333 5728 -3299
rect 5762 -3333 5796 -3299
rect 5830 -3333 5864 -3299
rect 5898 -3333 5932 -3299
rect 5966 -3333 6000 -3299
rect 6034 -3333 6068 -3299
rect 6102 -3333 6136 -3299
rect 6170 -3333 6204 -3299
rect 6238 -3333 6272 -3299
rect 6306 -3333 6340 -3299
rect 6374 -3333 6408 -3299
rect 6442 -3333 6476 -3299
rect 6510 -3333 6544 -3299
rect 6578 -3333 6612 -3299
rect 6646 -3333 6680 -3299
rect 6714 -3333 6748 -3299
rect 6782 -3333 6816 -3299
rect 6850 -3333 6884 -3299
rect 6918 -3333 6952 -3299
rect 6986 -3333 7020 -3299
rect 7054 -3333 7088 -3299
rect 7122 -3333 7156 -3299
rect 7190 -3333 7224 -3299
rect 7258 -3333 7292 -3299
rect 7326 -3333 7360 -3299
rect 7394 -3333 7428 -3299
rect 7462 -3333 7496 -3299
rect 7530 -3333 7564 -3299
rect 7598 -3333 7632 -3299
rect 7666 -3333 7700 -3299
rect 7734 -3333 7768 -3299
rect 7802 -3333 7836 -3299
rect 7870 -3333 7904 -3299
rect 7938 -3333 7972 -3299
rect 8006 -3333 8040 -3299
rect 8074 -3333 8108 -3299
rect 8142 -3333 8176 -3299
rect 8210 -3333 8244 -3299
rect 8278 -3333 8312 -3299
rect 8346 -3333 8380 -3299
rect 8414 -3333 8448 -3299
rect 8482 -3333 8516 -3299
rect 8550 -3333 8584 -3299
rect 8618 -3333 8652 -3299
rect 8686 -3333 8720 -3299
rect 8754 -3333 8788 -3299
rect 8822 -3333 8856 -3299
rect 8890 -3333 8924 -3299
rect 8958 -3333 8992 -3299
rect 9026 -3333 9060 -3299
rect 9094 -3333 9128 -3299
rect 9162 -3333 9196 -3299
rect 9230 -3333 9264 -3299
rect 9298 -3333 9332 -3299
rect 9366 -3333 9400 -3299
rect 9434 -3333 9468 -3299
rect 9502 -3333 9623 -3299
rect 872 -3401 906 -3367
rect 872 -3469 906 -3435
rect 872 -3537 906 -3503
rect 872 -3605 906 -3571
rect 872 -3673 906 -3639
rect 5231 -3401 5265 -3367
rect 5231 -3469 5265 -3435
rect 5231 -3537 5265 -3503
rect 5231 -3605 5265 -3571
rect 5231 -3673 5265 -3639
rect 872 -3741 906 -3707
rect 9589 -3401 9623 -3367
rect 9589 -3469 9623 -3435
rect 9589 -3537 9623 -3503
rect 9589 -3605 9623 -3571
rect 9589 -3673 9623 -3639
rect 872 -3809 906 -3775
rect 872 -4072 906 -3843
rect 5231 -3741 5265 -3707
rect 5231 -3809 5265 -3775
rect 5231 -4072 5265 -3843
rect 9589 -3741 9623 -3707
rect 9589 -3809 9623 -3775
rect 9589 -4072 9623 -3843
rect 872 -4106 993 -4072
rect 1027 -4106 1061 -4072
rect 1095 -4106 1129 -4072
rect 1163 -4106 1197 -4072
rect 1231 -4106 1265 -4072
rect 1299 -4106 1333 -4072
rect 1367 -4106 1401 -4072
rect 1435 -4106 1469 -4072
rect 1503 -4106 1537 -4072
rect 1571 -4106 1605 -4072
rect 1639 -4106 1673 -4072
rect 1707 -4106 1741 -4072
rect 1775 -4106 1809 -4072
rect 1843 -4106 1877 -4072
rect 1911 -4106 1945 -4072
rect 1979 -4106 2013 -4072
rect 2047 -4106 2081 -4072
rect 2115 -4106 2149 -4072
rect 2183 -4106 2217 -4072
rect 2251 -4106 2285 -4072
rect 2319 -4106 2353 -4072
rect 2387 -4106 2421 -4072
rect 2455 -4106 2489 -4072
rect 2523 -4106 2557 -4072
rect 2591 -4106 2625 -4072
rect 2659 -4106 2693 -4072
rect 2727 -4106 2761 -4072
rect 2795 -4106 2829 -4072
rect 2863 -4106 2897 -4072
rect 2931 -4106 2965 -4072
rect 2999 -4106 3033 -4072
rect 3067 -4106 3101 -4072
rect 3135 -4106 3169 -4072
rect 3203 -4106 3237 -4072
rect 3271 -4106 3305 -4072
rect 3339 -4106 3373 -4072
rect 3407 -4106 3441 -4072
rect 3475 -4106 3509 -4072
rect 3543 -4106 3577 -4072
rect 3611 -4106 3645 -4072
rect 3679 -4106 3713 -4072
rect 3747 -4106 3781 -4072
rect 3815 -4106 3849 -4072
rect 3883 -4106 3917 -4072
rect 3951 -4106 3985 -4072
rect 4019 -4106 4053 -4072
rect 4087 -4106 4121 -4072
rect 4155 -4106 4189 -4072
rect 4223 -4106 4257 -4072
rect 4291 -4106 4325 -4072
rect 4359 -4106 4393 -4072
rect 4427 -4106 4461 -4072
rect 4495 -4106 4529 -4072
rect 4563 -4106 4597 -4072
rect 4631 -4106 4665 -4072
rect 4699 -4106 4733 -4072
rect 4767 -4106 4801 -4072
rect 4835 -4106 4869 -4072
rect 4903 -4106 4937 -4072
rect 4971 -4106 5005 -4072
rect 5039 -4106 5073 -4072
rect 5107 -4106 5388 -4072
rect 5422 -4106 5456 -4072
rect 5490 -4106 5524 -4072
rect 5558 -4106 5592 -4072
rect 5626 -4106 5660 -4072
rect 5694 -4106 5728 -4072
rect 5762 -4106 5796 -4072
rect 5830 -4106 5864 -4072
rect 5898 -4106 5932 -4072
rect 5966 -4106 6000 -4072
rect 6034 -4106 6068 -4072
rect 6102 -4106 6136 -4072
rect 6170 -4106 6204 -4072
rect 6238 -4106 6272 -4072
rect 6306 -4106 6340 -4072
rect 6374 -4106 6408 -4072
rect 6442 -4106 6476 -4072
rect 6510 -4106 6544 -4072
rect 6578 -4106 6612 -4072
rect 6646 -4106 6680 -4072
rect 6714 -4106 6748 -4072
rect 6782 -4106 6816 -4072
rect 6850 -4106 6884 -4072
rect 6918 -4106 6952 -4072
rect 6986 -4106 7020 -4072
rect 7054 -4106 7088 -4072
rect 7122 -4106 7156 -4072
rect 7190 -4106 7224 -4072
rect 7258 -4106 7292 -4072
rect 7326 -4106 7360 -4072
rect 7394 -4106 7428 -4072
rect 7462 -4106 7496 -4072
rect 7530 -4106 7564 -4072
rect 7598 -4106 7632 -4072
rect 7666 -4106 7700 -4072
rect 7734 -4106 7768 -4072
rect 7802 -4106 7836 -4072
rect 7870 -4106 7904 -4072
rect 7938 -4106 7972 -4072
rect 8006 -4106 8040 -4072
rect 8074 -4106 8108 -4072
rect 8142 -4106 8176 -4072
rect 8210 -4106 8244 -4072
rect 8278 -4106 8312 -4072
rect 8346 -4106 8380 -4072
rect 8414 -4106 8448 -4072
rect 8482 -4106 8516 -4072
rect 8550 -4106 8584 -4072
rect 8618 -4106 8652 -4072
rect 8686 -4106 8720 -4072
rect 8754 -4106 8788 -4072
rect 8822 -4106 8856 -4072
rect 8890 -4106 8924 -4072
rect 8958 -4106 8992 -4072
rect 9026 -4106 9060 -4072
rect 9094 -4106 9128 -4072
rect 9162 -4106 9196 -4072
rect 9230 -4106 9264 -4072
rect 9298 -4106 9332 -4072
rect 9366 -4106 9400 -4072
rect 9434 -4106 9468 -4072
rect 9502 -4106 9623 -4072
rect 872 -4335 906 -4106
rect 872 -4403 906 -4369
rect 872 -4471 906 -4437
rect 5231 -4335 5265 -4106
rect 5231 -4403 5265 -4369
rect 5231 -4471 5265 -4437
rect 9589 -4335 9623 -4106
rect 9589 -4403 9623 -4369
rect 872 -4539 906 -4505
rect 872 -4607 906 -4573
rect 872 -4675 906 -4641
rect 872 -4743 906 -4709
rect 872 -4811 906 -4777
rect 9589 -4471 9623 -4437
rect 5231 -4539 5265 -4505
rect 5231 -4607 5265 -4573
rect 5231 -4675 5265 -4641
rect 5231 -4743 5265 -4709
rect 5231 -4811 5265 -4777
rect 9589 -4539 9623 -4505
rect 9589 -4607 9623 -4573
rect 9589 -4675 9623 -4641
rect 9589 -4743 9623 -4709
rect 9589 -4811 9623 -4777
rect 872 -4879 993 -4845
rect 1027 -4879 1061 -4845
rect 1095 -4879 1129 -4845
rect 1163 -4879 1197 -4845
rect 1231 -4879 1265 -4845
rect 1299 -4879 1333 -4845
rect 1367 -4879 1401 -4845
rect 1435 -4879 1469 -4845
rect 1503 -4879 1537 -4845
rect 1571 -4879 1605 -4845
rect 1639 -4879 1673 -4845
rect 1707 -4879 1741 -4845
rect 1775 -4879 1809 -4845
rect 1843 -4879 1877 -4845
rect 1911 -4879 1945 -4845
rect 1979 -4879 2013 -4845
rect 2047 -4879 2081 -4845
rect 2115 -4879 2149 -4845
rect 2183 -4879 2217 -4845
rect 2251 -4879 2285 -4845
rect 2319 -4879 2353 -4845
rect 2387 -4879 2421 -4845
rect 2455 -4879 2489 -4845
rect 2523 -4879 2557 -4845
rect 2591 -4879 2625 -4845
rect 2659 -4879 2693 -4845
rect 2727 -4879 2761 -4845
rect 2795 -4879 2829 -4845
rect 2863 -4879 2897 -4845
rect 2931 -4879 2965 -4845
rect 2999 -4879 3033 -4845
rect 3067 -4879 3101 -4845
rect 3135 -4879 3169 -4845
rect 3203 -4879 3237 -4845
rect 3271 -4879 3305 -4845
rect 3339 -4879 3373 -4845
rect 3407 -4879 3441 -4845
rect 3475 -4879 3509 -4845
rect 3543 -4879 3577 -4845
rect 3611 -4879 3645 -4845
rect 3679 -4879 3713 -4845
rect 3747 -4879 3781 -4845
rect 3815 -4879 3849 -4845
rect 3883 -4879 3917 -4845
rect 3951 -4879 3985 -4845
rect 4019 -4879 4053 -4845
rect 4087 -4879 4121 -4845
rect 4155 -4879 4189 -4845
rect 4223 -4879 4257 -4845
rect 4291 -4879 4325 -4845
rect 4359 -4879 4393 -4845
rect 4427 -4879 4461 -4845
rect 4495 -4879 4529 -4845
rect 4563 -4879 4597 -4845
rect 4631 -4879 4665 -4845
rect 4699 -4879 4733 -4845
rect 4767 -4879 4801 -4845
rect 4835 -4879 4869 -4845
rect 4903 -4879 4937 -4845
rect 4971 -4879 5005 -4845
rect 5039 -4879 5073 -4845
rect 5107 -4879 5388 -4845
rect 5422 -4879 5456 -4845
rect 5490 -4879 5524 -4845
rect 5558 -4879 5592 -4845
rect 5626 -4879 5660 -4845
rect 5694 -4879 5728 -4845
rect 5762 -4879 5796 -4845
rect 5830 -4879 5864 -4845
rect 5898 -4879 5932 -4845
rect 5966 -4879 6000 -4845
rect 6034 -4879 6068 -4845
rect 6102 -4879 6136 -4845
rect 6170 -4879 6204 -4845
rect 6238 -4879 6272 -4845
rect 6306 -4879 6340 -4845
rect 6374 -4879 6408 -4845
rect 6442 -4879 6476 -4845
rect 6510 -4879 6544 -4845
rect 6578 -4879 6612 -4845
rect 6646 -4879 6680 -4845
rect 6714 -4879 6748 -4845
rect 6782 -4879 6816 -4845
rect 6850 -4879 6884 -4845
rect 6918 -4879 6952 -4845
rect 6986 -4879 7020 -4845
rect 7054 -4879 7088 -4845
rect 7122 -4879 7156 -4845
rect 7190 -4879 7224 -4845
rect 7258 -4879 7292 -4845
rect 7326 -4879 7360 -4845
rect 7394 -4879 7428 -4845
rect 7462 -4879 7496 -4845
rect 7530 -4879 7564 -4845
rect 7598 -4879 7632 -4845
rect 7666 -4879 7700 -4845
rect 7734 -4879 7768 -4845
rect 7802 -4879 7836 -4845
rect 7870 -4879 7904 -4845
rect 7938 -4879 7972 -4845
rect 8006 -4879 8040 -4845
rect 8074 -4879 8108 -4845
rect 8142 -4879 8176 -4845
rect 8210 -4879 8244 -4845
rect 8278 -4879 8312 -4845
rect 8346 -4879 8380 -4845
rect 8414 -4879 8448 -4845
rect 8482 -4879 8516 -4845
rect 8550 -4879 8584 -4845
rect 8618 -4879 8652 -4845
rect 8686 -4879 8720 -4845
rect 8754 -4879 8788 -4845
rect 8822 -4879 8856 -4845
rect 8890 -4879 8924 -4845
rect 8958 -4879 8992 -4845
rect 9026 -4879 9060 -4845
rect 9094 -4879 9128 -4845
rect 9162 -4879 9196 -4845
rect 9230 -4879 9264 -4845
rect 9298 -4879 9332 -4845
rect 9366 -4879 9400 -4845
rect 9434 -4879 9468 -4845
rect 9502 -4879 9623 -4845
rect 872 -4947 906 -4913
rect 872 -5015 906 -4981
rect 872 -5083 906 -5049
rect 872 -5151 906 -5117
rect 872 -5219 906 -5185
rect 5231 -4947 5265 -4913
rect 5231 -5015 5265 -4981
rect 5231 -5083 5265 -5049
rect 5231 -5151 5265 -5117
rect 5231 -5219 5265 -5185
rect 872 -5287 906 -5253
rect 9589 -4947 9623 -4913
rect 9589 -5015 9623 -4981
rect 9589 -5083 9623 -5049
rect 9589 -5151 9623 -5117
rect 9589 -5219 9623 -5185
rect 872 -5355 906 -5321
rect 872 -5423 906 -5389
rect 5231 -5287 5265 -5253
rect 5231 -5355 5265 -5321
rect 5231 -5423 5265 -5389
rect 9589 -5287 9623 -5253
rect 9589 -5355 9623 -5321
rect 9589 -5423 9623 -5389
rect 872 -5491 906 -5457
rect 872 -5559 906 -5525
rect 5231 -5491 5265 -5457
rect 872 -5627 906 -5593
rect 872 -5695 906 -5661
rect 872 -5763 906 -5729
rect 872 -5831 906 -5797
rect 5231 -5559 5265 -5525
rect 9589 -5491 9623 -5457
rect 5231 -5627 5265 -5593
rect 5231 -5695 5265 -5661
rect 5231 -5763 5265 -5729
rect 5231 -5831 5265 -5797
rect 872 -5899 906 -5865
rect 872 -5967 906 -5933
rect 9589 -5559 9623 -5525
rect 9589 -5627 9623 -5593
rect 9589 -5695 9623 -5661
rect 9589 -5763 9623 -5729
rect 9589 -5831 9623 -5797
rect 5231 -5899 5265 -5865
rect 872 -6035 906 -6001
rect 872 -6103 906 -6069
rect 872 -6171 906 -6137
rect 5231 -5967 5265 -5933
rect 9589 -5899 9623 -5865
rect 5231 -6035 5265 -6001
rect 5231 -6103 5265 -6069
rect 5231 -6171 5265 -6137
rect 9589 -5967 9623 -5933
rect 9589 -6035 9623 -6001
rect 9589 -6103 9623 -6069
rect 872 -6239 906 -6205
rect 872 -6307 906 -6273
rect 872 -6375 906 -6341
rect 872 -6511 906 -6409
rect 9589 -6171 9623 -6137
rect 5231 -6239 5265 -6205
rect 5231 -6307 5265 -6273
rect 5231 -6375 5265 -6341
rect 5231 -6511 5265 -6409
rect 9589 -6239 9623 -6205
rect 9589 -6307 9623 -6273
rect 9589 -6375 9623 -6341
rect 9589 -6511 9623 -6409
rect 872 -6545 993 -6511
rect 1027 -6545 1061 -6511
rect 1095 -6545 1129 -6511
rect 1163 -6545 1197 -6511
rect 1231 -6545 1265 -6511
rect 1299 -6545 1333 -6511
rect 1367 -6545 1401 -6511
rect 1435 -6545 1469 -6511
rect 1503 -6545 1537 -6511
rect 1571 -6545 1605 -6511
rect 1639 -6545 1673 -6511
rect 1707 -6545 1741 -6511
rect 1775 -6545 1809 -6511
rect 1843 -6545 1877 -6511
rect 1911 -6545 1945 -6511
rect 1979 -6545 2013 -6511
rect 2047 -6545 2081 -6511
rect 2115 -6545 2149 -6511
rect 2183 -6545 2217 -6511
rect 2251 -6545 2285 -6511
rect 2319 -6545 2353 -6511
rect 2387 -6545 2421 -6511
rect 2455 -6545 2489 -6511
rect 2523 -6545 2557 -6511
rect 2591 -6545 2625 -6511
rect 2659 -6545 2693 -6511
rect 2727 -6545 2761 -6511
rect 2795 -6545 2829 -6511
rect 2863 -6545 2897 -6511
rect 2931 -6545 2965 -6511
rect 2999 -6545 3033 -6511
rect 3067 -6545 3101 -6511
rect 3135 -6545 3169 -6511
rect 3203 -6545 3237 -6511
rect 3271 -6545 3305 -6511
rect 3339 -6545 3373 -6511
rect 3407 -6545 3441 -6511
rect 3475 -6545 3509 -6511
rect 3543 -6545 3577 -6511
rect 3611 -6545 3645 -6511
rect 3679 -6545 3713 -6511
rect 3747 -6545 3781 -6511
rect 3815 -6545 3849 -6511
rect 3883 -6545 3917 -6511
rect 3951 -6545 3985 -6511
rect 4019 -6545 4053 -6511
rect 4087 -6545 4121 -6511
rect 4155 -6545 4189 -6511
rect 4223 -6545 4257 -6511
rect 4291 -6545 4325 -6511
rect 4359 -6545 4393 -6511
rect 4427 -6545 4461 -6511
rect 4495 -6545 4529 -6511
rect 4563 -6545 4597 -6511
rect 4631 -6545 4665 -6511
rect 4699 -6545 4733 -6511
rect 4767 -6545 4801 -6511
rect 4835 -6545 4869 -6511
rect 4903 -6545 4937 -6511
rect 4971 -6545 5005 -6511
rect 5039 -6545 5073 -6511
rect 5107 -6545 5388 -6511
rect 5422 -6545 5456 -6511
rect 5490 -6545 5524 -6511
rect 5558 -6545 5592 -6511
rect 5626 -6545 5660 -6511
rect 5694 -6545 5728 -6511
rect 5762 -6545 5796 -6511
rect 5830 -6545 5864 -6511
rect 5898 -6545 5932 -6511
rect 5966 -6545 6000 -6511
rect 6034 -6545 6068 -6511
rect 6102 -6545 6136 -6511
rect 6170 -6545 6204 -6511
rect 6238 -6545 6272 -6511
rect 6306 -6545 6340 -6511
rect 6374 -6545 6408 -6511
rect 6442 -6545 6476 -6511
rect 6510 -6545 6544 -6511
rect 6578 -6545 6612 -6511
rect 6646 -6545 6680 -6511
rect 6714 -6545 6748 -6511
rect 6782 -6545 6816 -6511
rect 6850 -6545 6884 -6511
rect 6918 -6545 6952 -6511
rect 6986 -6545 7020 -6511
rect 7054 -6545 7088 -6511
rect 7122 -6545 7156 -6511
rect 7190 -6545 7224 -6511
rect 7258 -6545 7292 -6511
rect 7326 -6545 7360 -6511
rect 7394 -6545 7428 -6511
rect 7462 -6545 7496 -6511
rect 7530 -6545 7564 -6511
rect 7598 -6545 7632 -6511
rect 7666 -6545 7700 -6511
rect 7734 -6545 7768 -6511
rect 7802 -6545 7836 -6511
rect 7870 -6545 7904 -6511
rect 7938 -6545 7972 -6511
rect 8006 -6545 8040 -6511
rect 8074 -6545 8108 -6511
rect 8142 -6545 8176 -6511
rect 8210 -6545 8244 -6511
rect 8278 -6545 8312 -6511
rect 8346 -6545 8380 -6511
rect 8414 -6545 8448 -6511
rect 8482 -6545 8516 -6511
rect 8550 -6545 8584 -6511
rect 8618 -6545 8652 -6511
rect 8686 -6545 8720 -6511
rect 8754 -6545 8788 -6511
rect 8822 -6545 8856 -6511
rect 8890 -6545 8924 -6511
rect 8958 -6545 8992 -6511
rect 9026 -6545 9060 -6511
rect 9094 -6545 9128 -6511
rect 9162 -6545 9196 -6511
rect 9230 -6545 9264 -6511
rect 9298 -6545 9332 -6511
rect 9366 -6545 9400 -6511
rect 9434 -6545 9468 -6511
rect 9502 -6545 9623 -6511
rect 872 -6647 906 -6545
rect 872 -6715 906 -6681
rect 872 -6783 906 -6749
rect 872 -6851 906 -6817
rect 5231 -6647 5265 -6545
rect 5231 -6715 5265 -6681
rect 5231 -6783 5265 -6749
rect 5231 -6851 5265 -6817
rect 872 -6919 906 -6885
rect 9589 -6647 9623 -6545
rect 9589 -6715 9623 -6681
rect 9589 -6783 9623 -6749
rect 9589 -6851 9623 -6817
rect 872 -6987 906 -6953
rect 872 -7055 906 -7021
rect 872 -7123 906 -7089
rect 5231 -6919 5265 -6885
rect 5231 -6987 5265 -6953
rect 5231 -7055 5265 -7021
rect 872 -7191 906 -7157
rect 5231 -7123 5265 -7089
rect 9589 -6919 9623 -6885
rect 9589 -6987 9623 -6953
rect 9589 -7055 9623 -7021
rect 5231 -7191 5265 -7157
rect 872 -7259 906 -7225
rect 872 -7327 906 -7293
rect 872 -7395 906 -7361
rect 872 -7463 906 -7429
rect 9589 -7123 9623 -7089
rect 9589 -7191 9623 -7157
rect 5231 -7259 5265 -7225
rect 5231 -7327 5265 -7293
rect 5231 -7395 5265 -7361
rect 5231 -7463 5265 -7429
rect 9589 -7259 9623 -7225
rect 9589 -7327 9623 -7293
rect 9589 -7395 9623 -7361
rect 9589 -7463 9623 -7429
rect 872 -7531 906 -7497
rect 872 -7599 906 -7565
rect 5231 -7531 5265 -7497
rect 872 -7667 906 -7633
rect 872 -7735 906 -7701
rect 872 -7803 906 -7769
rect 5231 -7599 5265 -7565
rect 9589 -7531 9623 -7497
rect 5231 -7667 5265 -7633
rect 5231 -7735 5265 -7701
rect 5231 -7803 5265 -7769
rect 9589 -7599 9623 -7565
rect 9589 -7667 9623 -7633
rect 9589 -7735 9623 -7701
rect 872 -7871 906 -7837
rect 872 -7939 906 -7905
rect 872 -8007 906 -7973
rect 872 -8075 906 -8041
rect 9589 -7803 9623 -7769
rect 5231 -7871 5265 -7837
rect 5231 -7939 5265 -7905
rect 5231 -8007 5265 -7973
rect 5231 -8075 5265 -8041
rect 9589 -7871 9623 -7837
rect 9589 -7939 9623 -7905
rect 9589 -8007 9623 -7973
rect 9589 -8075 9623 -8041
rect 872 -8143 993 -8109
rect 1027 -8143 1061 -8109
rect 1095 -8143 1129 -8109
rect 1163 -8143 1197 -8109
rect 1231 -8143 1265 -8109
rect 1299 -8143 1333 -8109
rect 1367 -8143 1401 -8109
rect 1435 -8143 1469 -8109
rect 1503 -8143 1537 -8109
rect 1571 -8143 1605 -8109
rect 1639 -8143 1673 -8109
rect 1707 -8143 1741 -8109
rect 1775 -8143 1809 -8109
rect 1843 -8143 1877 -8109
rect 1911 -8143 1945 -8109
rect 1979 -8143 2013 -8109
rect 2047 -8143 2081 -8109
rect 2115 -8143 2149 -8109
rect 2183 -8143 2217 -8109
rect 2251 -8143 2285 -8109
rect 2319 -8143 2353 -8109
rect 2387 -8143 2421 -8109
rect 2455 -8143 2489 -8109
rect 2523 -8143 2557 -8109
rect 2591 -8143 2625 -8109
rect 2659 -8143 2693 -8109
rect 2727 -8143 2761 -8109
rect 2795 -8143 2829 -8109
rect 2863 -8143 2897 -8109
rect 2931 -8143 2965 -8109
rect 2999 -8143 3033 -8109
rect 3067 -8143 3101 -8109
rect 3135 -8143 3169 -8109
rect 3203 -8143 3237 -8109
rect 3271 -8143 3305 -8109
rect 3339 -8143 3373 -8109
rect 3407 -8143 3441 -8109
rect 3475 -8143 3509 -8109
rect 3543 -8143 3577 -8109
rect 3611 -8143 3645 -8109
rect 3679 -8143 3713 -8109
rect 3747 -8143 3781 -8109
rect 3815 -8143 3849 -8109
rect 3883 -8143 3917 -8109
rect 3951 -8143 3985 -8109
rect 4019 -8143 4053 -8109
rect 4087 -8143 4121 -8109
rect 4155 -8143 4189 -8109
rect 4223 -8143 4257 -8109
rect 4291 -8143 4325 -8109
rect 4359 -8143 4393 -8109
rect 4427 -8143 4461 -8109
rect 4495 -8143 4529 -8109
rect 4563 -8143 4597 -8109
rect 4631 -8143 4665 -8109
rect 4699 -8143 4733 -8109
rect 4767 -8143 4801 -8109
rect 4835 -8143 4869 -8109
rect 4903 -8143 4937 -8109
rect 4971 -8143 5005 -8109
rect 5039 -8143 5073 -8109
rect 5107 -8143 5388 -8109
rect 5422 -8143 5456 -8109
rect 5490 -8143 5524 -8109
rect 5558 -8143 5592 -8109
rect 5626 -8143 5660 -8109
rect 5694 -8143 5728 -8109
rect 5762 -8143 5796 -8109
rect 5830 -8143 5864 -8109
rect 5898 -8143 5932 -8109
rect 5966 -8143 6000 -8109
rect 6034 -8143 6068 -8109
rect 6102 -8143 6136 -8109
rect 6170 -8143 6204 -8109
rect 6238 -8143 6272 -8109
rect 6306 -8143 6340 -8109
rect 6374 -8143 6408 -8109
rect 6442 -8143 6476 -8109
rect 6510 -8143 6544 -8109
rect 6578 -8143 6612 -8109
rect 6646 -8143 6680 -8109
rect 6714 -8143 6748 -8109
rect 6782 -8143 6816 -8109
rect 6850 -8143 6884 -8109
rect 6918 -8143 6952 -8109
rect 6986 -8143 7020 -8109
rect 7054 -8143 7088 -8109
rect 7122 -8143 7156 -8109
rect 7190 -8143 7224 -8109
rect 7258 -8143 7292 -8109
rect 7326 -8143 7360 -8109
rect 7394 -8143 7428 -8109
rect 7462 -8143 7496 -8109
rect 7530 -8143 7564 -8109
rect 7598 -8143 7632 -8109
rect 7666 -8143 7700 -8109
rect 7734 -8143 7768 -8109
rect 7802 -8143 7836 -8109
rect 7870 -8143 7904 -8109
rect 7938 -8143 7972 -8109
rect 8006 -8143 8040 -8109
rect 8074 -8143 8108 -8109
rect 8142 -8143 8176 -8109
rect 8210 -8143 8244 -8109
rect 8278 -8143 8312 -8109
rect 8346 -8143 8380 -8109
rect 8414 -8143 8448 -8109
rect 8482 -8143 8516 -8109
rect 8550 -8143 8584 -8109
rect 8618 -8143 8652 -8109
rect 8686 -8143 8720 -8109
rect 8754 -8143 8788 -8109
rect 8822 -8143 8856 -8109
rect 8890 -8143 8924 -8109
rect 8958 -8143 8992 -8109
rect 9026 -8143 9060 -8109
rect 9094 -8143 9128 -8109
rect 9162 -8143 9196 -8109
rect 9230 -8143 9264 -8109
rect 9298 -8143 9332 -8109
rect 9366 -8143 9400 -8109
rect 9434 -8143 9468 -8109
rect 9502 -8143 9623 -8109
rect 872 -8211 906 -8177
rect 872 -8279 906 -8245
rect 872 -8347 906 -8313
rect 872 -8415 906 -8381
rect 872 -8483 906 -8449
rect 5231 -8211 5265 -8177
rect 5231 -8279 5265 -8245
rect 5231 -8347 5265 -8313
rect 5231 -8415 5265 -8381
rect 5231 -8483 5265 -8449
rect 872 -8551 906 -8517
rect 9589 -8211 9623 -8177
rect 9589 -8279 9623 -8245
rect 9589 -8347 9623 -8313
rect 9589 -8415 9623 -8381
rect 9589 -8483 9623 -8449
rect 872 -8619 906 -8585
rect 872 -8687 906 -8653
rect 872 -8899 906 -8721
rect 5231 -8551 5265 -8517
rect 5231 -8619 5265 -8585
rect 5231 -8687 5265 -8653
rect 5231 -8899 5265 -8721
rect 9589 -8551 9623 -8517
rect 9589 -8619 9623 -8585
rect 9589 -8687 9623 -8653
rect 9589 -8899 9623 -8721
rect 872 -8933 993 -8899
rect 1027 -8933 1061 -8899
rect 1095 -8933 1129 -8899
rect 1163 -8933 1197 -8899
rect 1231 -8933 1265 -8899
rect 1299 -8933 1333 -8899
rect 1367 -8933 1401 -8899
rect 1435 -8933 1469 -8899
rect 1503 -8933 1537 -8899
rect 1571 -8933 1605 -8899
rect 1639 -8933 1673 -8899
rect 1707 -8933 1741 -8899
rect 1775 -8933 1809 -8899
rect 1843 -8933 1877 -8899
rect 1911 -8933 1945 -8899
rect 1979 -8933 2013 -8899
rect 2047 -8933 2081 -8899
rect 2115 -8933 2149 -8899
rect 2183 -8933 2217 -8899
rect 2251 -8933 2285 -8899
rect 2319 -8933 2353 -8899
rect 2387 -8933 2421 -8899
rect 2455 -8933 2489 -8899
rect 2523 -8933 2557 -8899
rect 2591 -8933 2625 -8899
rect 2659 -8933 2693 -8899
rect 2727 -8933 2761 -8899
rect 2795 -8933 2829 -8899
rect 2863 -8933 2897 -8899
rect 2931 -8933 2965 -8899
rect 2999 -8933 3033 -8899
rect 3067 -8933 3101 -8899
rect 3135 -8933 3169 -8899
rect 3203 -8933 3237 -8899
rect 3271 -8933 3305 -8899
rect 3339 -8933 3373 -8899
rect 3407 -8933 3441 -8899
rect 3475 -8933 3509 -8899
rect 3543 -8933 3577 -8899
rect 3611 -8933 3645 -8899
rect 3679 -8933 3713 -8899
rect 3747 -8933 3781 -8899
rect 3815 -8933 3849 -8899
rect 3883 -8933 3917 -8899
rect 3951 -8933 3985 -8899
rect 4019 -8933 4053 -8899
rect 4087 -8933 4121 -8899
rect 4155 -8933 4189 -8899
rect 4223 -8933 4257 -8899
rect 4291 -8933 4325 -8899
rect 4359 -8933 4393 -8899
rect 4427 -8933 4461 -8899
rect 4495 -8933 4529 -8899
rect 4563 -8933 4597 -8899
rect 4631 -8933 4665 -8899
rect 4699 -8933 4733 -8899
rect 4767 -8933 4801 -8899
rect 4835 -8933 4869 -8899
rect 4903 -8933 4937 -8899
rect 4971 -8933 5005 -8899
rect 5039 -8933 5073 -8899
rect 5107 -8933 5388 -8899
rect 5422 -8933 5456 -8899
rect 5490 -8933 5524 -8899
rect 5558 -8933 5592 -8899
rect 5626 -8933 5660 -8899
rect 5694 -8933 5728 -8899
rect 5762 -8933 5796 -8899
rect 5830 -8933 5864 -8899
rect 5898 -8933 5932 -8899
rect 5966 -8933 6000 -8899
rect 6034 -8933 6068 -8899
rect 6102 -8933 6136 -8899
rect 6170 -8933 6204 -8899
rect 6238 -8933 6272 -8899
rect 6306 -8933 6340 -8899
rect 6374 -8933 6408 -8899
rect 6442 -8933 6476 -8899
rect 6510 -8933 6544 -8899
rect 6578 -8933 6612 -8899
rect 6646 -8933 6680 -8899
rect 6714 -8933 6748 -8899
rect 6782 -8933 6816 -8899
rect 6850 -8933 6884 -8899
rect 6918 -8933 6952 -8899
rect 6986 -8933 7020 -8899
rect 7054 -8933 7088 -8899
rect 7122 -8933 7156 -8899
rect 7190 -8933 7224 -8899
rect 7258 -8933 7292 -8899
rect 7326 -8933 7360 -8899
rect 7394 -8933 7428 -8899
rect 7462 -8933 7496 -8899
rect 7530 -8933 7564 -8899
rect 7598 -8933 7632 -8899
rect 7666 -8933 7700 -8899
rect 7734 -8933 7768 -8899
rect 7802 -8933 7836 -8899
rect 7870 -8933 7904 -8899
rect 7938 -8933 7972 -8899
rect 8006 -8933 8040 -8899
rect 8074 -8933 8108 -8899
rect 8142 -8933 8176 -8899
rect 8210 -8933 8244 -8899
rect 8278 -8933 8312 -8899
rect 8346 -8933 8380 -8899
rect 8414 -8933 8448 -8899
rect 8482 -8933 8516 -8899
rect 8550 -8933 8584 -8899
rect 8618 -8933 8652 -8899
rect 8686 -8933 8720 -8899
rect 8754 -8933 8788 -8899
rect 8822 -8933 8856 -8899
rect 8890 -8933 8924 -8899
rect 8958 -8933 8992 -8899
rect 9026 -8933 9060 -8899
rect 9094 -8933 9128 -8899
rect 9162 -8933 9196 -8899
rect 9230 -8933 9264 -8899
rect 9298 -8933 9332 -8899
rect 9366 -8933 9400 -8899
rect 9434 -8933 9468 -8899
rect 9502 -8933 9623 -8899
<< nsubdiffcont >>
rect 993 722 1027 756
rect 1061 722 1095 756
rect 1129 722 1163 756
rect 1197 722 1231 756
rect 1265 722 1299 756
rect 1333 722 1367 756
rect 1401 722 1435 756
rect 1469 722 1503 756
rect 1537 722 1571 756
rect 1605 722 1639 756
rect 1673 722 1707 756
rect 1741 722 1775 756
rect 1809 722 1843 756
rect 1877 722 1911 756
rect 1945 722 1979 756
rect 2013 722 2047 756
rect 2081 722 2115 756
rect 2149 722 2183 756
rect 2217 722 2251 756
rect 2285 722 2319 756
rect 2353 722 2387 756
rect 2421 722 2455 756
rect 2489 722 2523 756
rect 2557 722 2591 756
rect 2625 722 2659 756
rect 2693 722 2727 756
rect 2761 722 2795 756
rect 2829 722 2863 756
rect 2897 722 2931 756
rect 2965 722 2999 756
rect 3033 722 3067 756
rect 3101 722 3135 756
rect 3169 722 3203 756
rect 3237 722 3271 756
rect 3305 722 3339 756
rect 3373 722 3407 756
rect 3441 722 3475 756
rect 3509 722 3543 756
rect 3577 722 3611 756
rect 3645 722 3679 756
rect 3713 722 3747 756
rect 3781 722 3815 756
rect 3849 722 3883 756
rect 3917 722 3951 756
rect 3985 722 4019 756
rect 4053 722 4087 756
rect 4121 722 4155 756
rect 4189 722 4223 756
rect 4257 722 4291 756
rect 4325 722 4359 756
rect 4393 722 4427 756
rect 4461 722 4495 756
rect 4529 722 4563 756
rect 4597 722 4631 756
rect 4665 722 4699 756
rect 4733 722 4767 756
rect 4801 722 4835 756
rect 4869 722 4903 756
rect 4937 722 4971 756
rect 5005 722 5039 756
rect 5073 722 5107 756
rect 5388 722 5422 756
rect 5456 722 5490 756
rect 5524 722 5558 756
rect 5592 722 5626 756
rect 5660 722 5694 756
rect 5728 722 5762 756
rect 5796 722 5830 756
rect 5864 722 5898 756
rect 5932 722 5966 756
rect 6000 722 6034 756
rect 6068 722 6102 756
rect 6136 722 6170 756
rect 6204 722 6238 756
rect 6272 722 6306 756
rect 6340 722 6374 756
rect 6408 722 6442 756
rect 6476 722 6510 756
rect 6544 722 6578 756
rect 6612 722 6646 756
rect 6680 722 6714 756
rect 6748 722 6782 756
rect 6816 722 6850 756
rect 6884 722 6918 756
rect 6952 722 6986 756
rect 7020 722 7054 756
rect 7088 722 7122 756
rect 7156 722 7190 756
rect 7224 722 7258 756
rect 7292 722 7326 756
rect 7360 722 7394 756
rect 7428 722 7462 756
rect 7496 722 7530 756
rect 7564 722 7598 756
rect 7632 722 7666 756
rect 7700 722 7734 756
rect 7768 722 7802 756
rect 7836 722 7870 756
rect 7904 722 7938 756
rect 7972 722 8006 756
rect 8040 722 8074 756
rect 8108 722 8142 756
rect 8176 722 8210 756
rect 8244 722 8278 756
rect 8312 722 8346 756
rect 8380 722 8414 756
rect 8448 722 8482 756
rect 8516 722 8550 756
rect 8584 722 8618 756
rect 8652 722 8686 756
rect 8720 722 8754 756
rect 8788 722 8822 756
rect 8856 722 8890 756
rect 8924 722 8958 756
rect 8992 722 9026 756
rect 9060 722 9094 756
rect 9128 722 9162 756
rect 9196 722 9230 756
rect 9264 722 9298 756
rect 9332 722 9366 756
rect 9400 722 9434 756
rect 9468 722 9502 756
rect 872 509 906 543
rect 872 441 906 475
rect 872 373 906 407
rect 5231 509 5265 543
rect 5231 441 5265 475
rect 5231 373 5265 407
rect 872 305 906 339
rect 9589 509 9623 543
rect 9589 441 9623 475
rect 9589 373 9623 407
rect 872 237 906 271
rect 872 169 906 203
rect 872 101 906 135
rect 872 33 906 67
rect 872 -35 906 -1
rect 5231 305 5265 339
rect 5231 237 5265 271
rect 5231 169 5265 203
rect 5231 101 5265 135
rect 5231 33 5265 67
rect 5231 -35 5265 -1
rect 9589 305 9623 339
rect 9589 237 9623 271
rect 9589 169 9623 203
rect 9589 101 9623 135
rect 9589 33 9623 67
rect 9589 -35 9623 -1
rect 993 -69 1027 -35
rect 1061 -69 1095 -35
rect 1129 -69 1163 -35
rect 1197 -69 1231 -35
rect 1265 -69 1299 -35
rect 1333 -69 1367 -35
rect 1401 -69 1435 -35
rect 1469 -69 1503 -35
rect 1537 -69 1571 -35
rect 1605 -69 1639 -35
rect 1673 -69 1707 -35
rect 1741 -69 1775 -35
rect 1809 -69 1843 -35
rect 1877 -69 1911 -35
rect 1945 -69 1979 -35
rect 2013 -69 2047 -35
rect 2081 -69 2115 -35
rect 2149 -69 2183 -35
rect 2217 -69 2251 -35
rect 2285 -69 2319 -35
rect 2353 -69 2387 -35
rect 2421 -69 2455 -35
rect 2489 -69 2523 -35
rect 2557 -69 2591 -35
rect 2625 -69 2659 -35
rect 2693 -69 2727 -35
rect 2761 -69 2795 -35
rect 2829 -69 2863 -35
rect 2897 -69 2931 -35
rect 2965 -69 2999 -35
rect 3033 -69 3067 -35
rect 3101 -69 3135 -35
rect 3169 -69 3203 -35
rect 3237 -69 3271 -35
rect 3305 -69 3339 -35
rect 3373 -69 3407 -35
rect 3441 -69 3475 -35
rect 3509 -69 3543 -35
rect 3577 -69 3611 -35
rect 3645 -69 3679 -35
rect 3713 -69 3747 -35
rect 3781 -69 3815 -35
rect 3849 -69 3883 -35
rect 3917 -69 3951 -35
rect 3985 -69 4019 -35
rect 4053 -69 4087 -35
rect 4121 -69 4155 -35
rect 4189 -69 4223 -35
rect 4257 -69 4291 -35
rect 4325 -69 4359 -35
rect 4393 -69 4427 -35
rect 4461 -69 4495 -35
rect 4529 -69 4563 -35
rect 4597 -69 4631 -35
rect 4665 -69 4699 -35
rect 4733 -69 4767 -35
rect 4801 -69 4835 -35
rect 4869 -69 4903 -35
rect 4937 -69 4971 -35
rect 5005 -69 5039 -35
rect 5073 -69 5107 -35
rect 5388 -69 5422 -35
rect 5456 -69 5490 -35
rect 5524 -69 5558 -35
rect 5592 -69 5626 -35
rect 5660 -69 5694 -35
rect 5728 -69 5762 -35
rect 5796 -69 5830 -35
rect 5864 -69 5898 -35
rect 5932 -69 5966 -35
rect 6000 -69 6034 -35
rect 6068 -69 6102 -35
rect 6136 -69 6170 -35
rect 6204 -69 6238 -35
rect 6272 -69 6306 -35
rect 6340 -69 6374 -35
rect 6408 -69 6442 -35
rect 6476 -69 6510 -35
rect 6544 -69 6578 -35
rect 6612 -69 6646 -35
rect 6680 -69 6714 -35
rect 6748 -69 6782 -35
rect 6816 -69 6850 -35
rect 6884 -69 6918 -35
rect 6952 -69 6986 -35
rect 7020 -69 7054 -35
rect 7088 -69 7122 -35
rect 7156 -69 7190 -35
rect 7224 -69 7258 -35
rect 7292 -69 7326 -35
rect 7360 -69 7394 -35
rect 7428 -69 7462 -35
rect 7496 -69 7530 -35
rect 7564 -69 7598 -35
rect 7632 -69 7666 -35
rect 7700 -69 7734 -35
rect 7768 -69 7802 -35
rect 7836 -69 7870 -35
rect 7904 -69 7938 -35
rect 7972 -69 8006 -35
rect 8040 -69 8074 -35
rect 8108 -69 8142 -35
rect 8176 -69 8210 -35
rect 8244 -69 8278 -35
rect 8312 -69 8346 -35
rect 8380 -69 8414 -35
rect 8448 -69 8482 -35
rect 8516 -69 8550 -35
rect 8584 -69 8618 -35
rect 8652 -69 8686 -35
rect 8720 -69 8754 -35
rect 8788 -69 8822 -35
rect 8856 -69 8890 -35
rect 8924 -69 8958 -35
rect 8992 -69 9026 -35
rect 9060 -69 9094 -35
rect 9128 -69 9162 -35
rect 9196 -69 9230 -35
rect 9264 -69 9298 -35
rect 9332 -69 9366 -35
rect 9400 -69 9434 -35
rect 9468 -69 9502 -35
rect 872 -103 906 -69
rect 872 -171 906 -137
rect 872 -239 906 -205
rect 872 -307 906 -273
rect 872 -375 906 -341
rect 5231 -103 5265 -69
rect 5231 -171 5265 -137
rect 5231 -239 5265 -205
rect 5231 -307 5265 -273
rect 5231 -375 5265 -341
rect 9589 -103 9623 -69
rect 9589 -171 9623 -137
rect 9589 -239 9623 -205
rect 9589 -307 9623 -273
rect 872 -443 906 -409
rect 872 -511 906 -477
rect 872 -579 906 -545
rect 9589 -375 9623 -341
rect 5231 -443 5265 -409
rect 5231 -511 5265 -477
rect 5231 -579 5265 -545
rect 872 -647 906 -613
rect 9589 -443 9623 -409
rect 9589 -511 9623 -477
rect 9589 -579 9623 -545
rect 5231 -647 5265 -613
rect 872 -715 906 -681
rect 872 -783 906 -749
rect 872 -851 906 -817
rect 872 -919 906 -885
rect 872 -987 906 -953
rect 9589 -647 9623 -613
rect 5231 -715 5265 -681
rect 5231 -783 5265 -749
rect 5231 -851 5265 -817
rect 5231 -919 5265 -885
rect 872 -1055 906 -1021
rect 5231 -987 5265 -953
rect 9589 -715 9623 -681
rect 9589 -783 9623 -749
rect 9589 -851 9623 -817
rect 9589 -919 9623 -885
rect 5231 -1055 5265 -1021
rect 872 -1123 906 -1089
rect 872 -1191 906 -1157
rect 872 -1259 906 -1225
rect 9589 -987 9623 -953
rect 9589 -1055 9623 -1021
rect 5231 -1123 5265 -1089
rect 5231 -1191 5265 -1157
rect 5231 -1259 5265 -1225
rect 872 -1327 906 -1293
rect 9589 -1123 9623 -1089
rect 9589 -1191 9623 -1157
rect 9589 -1259 9623 -1225
rect 872 -1395 906 -1361
rect 872 -1463 906 -1429
rect 872 -1531 906 -1497
rect 5231 -1327 5265 -1293
rect 5231 -1395 5265 -1361
rect 5231 -1463 5265 -1429
rect 5231 -1531 5265 -1497
rect 9589 -1327 9623 -1293
rect 9589 -1395 9623 -1361
rect 9589 -1463 9623 -1429
rect 9589 -1531 9623 -1497
rect 993 -1667 1027 -1633
rect 1061 -1667 1095 -1633
rect 1129 -1667 1163 -1633
rect 1197 -1667 1231 -1633
rect 1265 -1667 1299 -1633
rect 1333 -1667 1367 -1633
rect 1401 -1667 1435 -1633
rect 1469 -1667 1503 -1633
rect 1537 -1667 1571 -1633
rect 1605 -1667 1639 -1633
rect 1673 -1667 1707 -1633
rect 1741 -1667 1775 -1633
rect 1809 -1667 1843 -1633
rect 1877 -1667 1911 -1633
rect 1945 -1667 1979 -1633
rect 2013 -1667 2047 -1633
rect 2081 -1667 2115 -1633
rect 2149 -1667 2183 -1633
rect 2217 -1667 2251 -1633
rect 2285 -1667 2319 -1633
rect 2353 -1667 2387 -1633
rect 2421 -1667 2455 -1633
rect 2489 -1667 2523 -1633
rect 2557 -1667 2591 -1633
rect 2625 -1667 2659 -1633
rect 2693 -1667 2727 -1633
rect 2761 -1667 2795 -1633
rect 2829 -1667 2863 -1633
rect 2897 -1667 2931 -1633
rect 2965 -1667 2999 -1633
rect 3033 -1667 3067 -1633
rect 3101 -1667 3135 -1633
rect 3169 -1667 3203 -1633
rect 3237 -1667 3271 -1633
rect 3305 -1667 3339 -1633
rect 3373 -1667 3407 -1633
rect 3441 -1667 3475 -1633
rect 3509 -1667 3543 -1633
rect 3577 -1667 3611 -1633
rect 3645 -1667 3679 -1633
rect 3713 -1667 3747 -1633
rect 3781 -1667 3815 -1633
rect 3849 -1667 3883 -1633
rect 3917 -1667 3951 -1633
rect 3985 -1667 4019 -1633
rect 4053 -1667 4087 -1633
rect 4121 -1667 4155 -1633
rect 4189 -1667 4223 -1633
rect 4257 -1667 4291 -1633
rect 4325 -1667 4359 -1633
rect 4393 -1667 4427 -1633
rect 4461 -1667 4495 -1633
rect 4529 -1667 4563 -1633
rect 4597 -1667 4631 -1633
rect 4665 -1667 4699 -1633
rect 4733 -1667 4767 -1633
rect 4801 -1667 4835 -1633
rect 4869 -1667 4903 -1633
rect 4937 -1667 4971 -1633
rect 5005 -1667 5039 -1633
rect 5073 -1667 5107 -1633
rect 5388 -1667 5422 -1633
rect 5456 -1667 5490 -1633
rect 5524 -1667 5558 -1633
rect 5592 -1667 5626 -1633
rect 5660 -1667 5694 -1633
rect 5728 -1667 5762 -1633
rect 5796 -1667 5830 -1633
rect 5864 -1667 5898 -1633
rect 5932 -1667 5966 -1633
rect 6000 -1667 6034 -1633
rect 6068 -1667 6102 -1633
rect 6136 -1667 6170 -1633
rect 6204 -1667 6238 -1633
rect 6272 -1667 6306 -1633
rect 6340 -1667 6374 -1633
rect 6408 -1667 6442 -1633
rect 6476 -1667 6510 -1633
rect 6544 -1667 6578 -1633
rect 6612 -1667 6646 -1633
rect 6680 -1667 6714 -1633
rect 6748 -1667 6782 -1633
rect 6816 -1667 6850 -1633
rect 6884 -1667 6918 -1633
rect 6952 -1667 6986 -1633
rect 7020 -1667 7054 -1633
rect 7088 -1667 7122 -1633
rect 7156 -1667 7190 -1633
rect 7224 -1667 7258 -1633
rect 7292 -1667 7326 -1633
rect 7360 -1667 7394 -1633
rect 7428 -1667 7462 -1633
rect 7496 -1667 7530 -1633
rect 7564 -1667 7598 -1633
rect 7632 -1667 7666 -1633
rect 7700 -1667 7734 -1633
rect 7768 -1667 7802 -1633
rect 7836 -1667 7870 -1633
rect 7904 -1667 7938 -1633
rect 7972 -1667 8006 -1633
rect 8040 -1667 8074 -1633
rect 8108 -1667 8142 -1633
rect 8176 -1667 8210 -1633
rect 8244 -1667 8278 -1633
rect 8312 -1667 8346 -1633
rect 8380 -1667 8414 -1633
rect 8448 -1667 8482 -1633
rect 8516 -1667 8550 -1633
rect 8584 -1667 8618 -1633
rect 8652 -1667 8686 -1633
rect 8720 -1667 8754 -1633
rect 8788 -1667 8822 -1633
rect 8856 -1667 8890 -1633
rect 8924 -1667 8958 -1633
rect 8992 -1667 9026 -1633
rect 9060 -1667 9094 -1633
rect 9128 -1667 9162 -1633
rect 9196 -1667 9230 -1633
rect 9264 -1667 9298 -1633
rect 9332 -1667 9366 -1633
rect 9400 -1667 9434 -1633
rect 9468 -1667 9502 -1633
rect 872 -1803 906 -1769
rect 872 -1871 906 -1837
rect 872 -1939 906 -1905
rect 872 -2007 906 -1973
rect 5231 -1803 5265 -1769
rect 5231 -1871 5265 -1837
rect 5231 -1939 5265 -1905
rect 5231 -2007 5265 -1973
rect 9589 -1803 9623 -1769
rect 9589 -1871 9623 -1837
rect 9589 -1939 9623 -1905
rect 872 -2075 906 -2041
rect 872 -2143 906 -2109
rect 872 -2211 906 -2177
rect 9589 -2007 9623 -1973
rect 5231 -2075 5265 -2041
rect 5231 -2143 5265 -2109
rect 5231 -2211 5265 -2177
rect 872 -2279 906 -2245
rect 872 -2347 906 -2313
rect 9589 -2075 9623 -2041
rect 9589 -2143 9623 -2109
rect 9589 -2211 9623 -2177
rect 5231 -2279 5265 -2245
rect 872 -2415 906 -2381
rect 872 -2483 906 -2449
rect 872 -2551 906 -2517
rect 872 -2619 906 -2585
rect 5231 -2347 5265 -2313
rect 9589 -2279 9623 -2245
rect 5231 -2415 5265 -2381
rect 5231 -2483 5265 -2449
rect 5231 -2551 5265 -2517
rect 5231 -2619 5265 -2585
rect 872 -2687 906 -2653
rect 9589 -2347 9623 -2313
rect 9589 -2415 9623 -2381
rect 9589 -2483 9623 -2449
rect 9589 -2551 9623 -2517
rect 9589 -2619 9623 -2585
rect 5231 -2687 5265 -2653
rect 9589 -2687 9623 -2653
rect 872 -2755 906 -2721
rect 872 -2823 906 -2789
rect 872 -2891 906 -2857
rect 5231 -2755 5265 -2721
rect 5231 -2823 5265 -2789
rect 5231 -2891 5265 -2857
rect 872 -2959 906 -2925
rect 9589 -2755 9623 -2721
rect 9589 -2823 9623 -2789
rect 9589 -2891 9623 -2857
rect 872 -3027 906 -2993
rect 872 -3095 906 -3061
rect 872 -3163 906 -3129
rect 872 -3231 906 -3197
rect 872 -3299 906 -3265
rect 5231 -2959 5265 -2925
rect 5231 -3027 5265 -2993
rect 5231 -3095 5265 -3061
rect 5231 -3163 5265 -3129
rect 5231 -3231 5265 -3197
rect 5231 -3299 5265 -3265
rect 9589 -2959 9623 -2925
rect 9589 -3027 9623 -2993
rect 9589 -3095 9623 -3061
rect 9589 -3163 9623 -3129
rect 9589 -3231 9623 -3197
rect 9589 -3299 9623 -3265
rect 993 -3333 1027 -3299
rect 1061 -3333 1095 -3299
rect 1129 -3333 1163 -3299
rect 1197 -3333 1231 -3299
rect 1265 -3333 1299 -3299
rect 1333 -3333 1367 -3299
rect 1401 -3333 1435 -3299
rect 1469 -3333 1503 -3299
rect 1537 -3333 1571 -3299
rect 1605 -3333 1639 -3299
rect 1673 -3333 1707 -3299
rect 1741 -3333 1775 -3299
rect 1809 -3333 1843 -3299
rect 1877 -3333 1911 -3299
rect 1945 -3333 1979 -3299
rect 2013 -3333 2047 -3299
rect 2081 -3333 2115 -3299
rect 2149 -3333 2183 -3299
rect 2217 -3333 2251 -3299
rect 2285 -3333 2319 -3299
rect 2353 -3333 2387 -3299
rect 2421 -3333 2455 -3299
rect 2489 -3333 2523 -3299
rect 2557 -3333 2591 -3299
rect 2625 -3333 2659 -3299
rect 2693 -3333 2727 -3299
rect 2761 -3333 2795 -3299
rect 2829 -3333 2863 -3299
rect 2897 -3333 2931 -3299
rect 2965 -3333 2999 -3299
rect 3033 -3333 3067 -3299
rect 3101 -3333 3135 -3299
rect 3169 -3333 3203 -3299
rect 3237 -3333 3271 -3299
rect 3305 -3333 3339 -3299
rect 3373 -3333 3407 -3299
rect 3441 -3333 3475 -3299
rect 3509 -3333 3543 -3299
rect 3577 -3333 3611 -3299
rect 3645 -3333 3679 -3299
rect 3713 -3333 3747 -3299
rect 3781 -3333 3815 -3299
rect 3849 -3333 3883 -3299
rect 3917 -3333 3951 -3299
rect 3985 -3333 4019 -3299
rect 4053 -3333 4087 -3299
rect 4121 -3333 4155 -3299
rect 4189 -3333 4223 -3299
rect 4257 -3333 4291 -3299
rect 4325 -3333 4359 -3299
rect 4393 -3333 4427 -3299
rect 4461 -3333 4495 -3299
rect 4529 -3333 4563 -3299
rect 4597 -3333 4631 -3299
rect 4665 -3333 4699 -3299
rect 4733 -3333 4767 -3299
rect 4801 -3333 4835 -3299
rect 4869 -3333 4903 -3299
rect 4937 -3333 4971 -3299
rect 5005 -3333 5039 -3299
rect 5073 -3333 5107 -3299
rect 5388 -3333 5422 -3299
rect 5456 -3333 5490 -3299
rect 5524 -3333 5558 -3299
rect 5592 -3333 5626 -3299
rect 5660 -3333 5694 -3299
rect 5728 -3333 5762 -3299
rect 5796 -3333 5830 -3299
rect 5864 -3333 5898 -3299
rect 5932 -3333 5966 -3299
rect 6000 -3333 6034 -3299
rect 6068 -3333 6102 -3299
rect 6136 -3333 6170 -3299
rect 6204 -3333 6238 -3299
rect 6272 -3333 6306 -3299
rect 6340 -3333 6374 -3299
rect 6408 -3333 6442 -3299
rect 6476 -3333 6510 -3299
rect 6544 -3333 6578 -3299
rect 6612 -3333 6646 -3299
rect 6680 -3333 6714 -3299
rect 6748 -3333 6782 -3299
rect 6816 -3333 6850 -3299
rect 6884 -3333 6918 -3299
rect 6952 -3333 6986 -3299
rect 7020 -3333 7054 -3299
rect 7088 -3333 7122 -3299
rect 7156 -3333 7190 -3299
rect 7224 -3333 7258 -3299
rect 7292 -3333 7326 -3299
rect 7360 -3333 7394 -3299
rect 7428 -3333 7462 -3299
rect 7496 -3333 7530 -3299
rect 7564 -3333 7598 -3299
rect 7632 -3333 7666 -3299
rect 7700 -3333 7734 -3299
rect 7768 -3333 7802 -3299
rect 7836 -3333 7870 -3299
rect 7904 -3333 7938 -3299
rect 7972 -3333 8006 -3299
rect 8040 -3333 8074 -3299
rect 8108 -3333 8142 -3299
rect 8176 -3333 8210 -3299
rect 8244 -3333 8278 -3299
rect 8312 -3333 8346 -3299
rect 8380 -3333 8414 -3299
rect 8448 -3333 8482 -3299
rect 8516 -3333 8550 -3299
rect 8584 -3333 8618 -3299
rect 8652 -3333 8686 -3299
rect 8720 -3333 8754 -3299
rect 8788 -3333 8822 -3299
rect 8856 -3333 8890 -3299
rect 8924 -3333 8958 -3299
rect 8992 -3333 9026 -3299
rect 9060 -3333 9094 -3299
rect 9128 -3333 9162 -3299
rect 9196 -3333 9230 -3299
rect 9264 -3333 9298 -3299
rect 9332 -3333 9366 -3299
rect 9400 -3333 9434 -3299
rect 9468 -3333 9502 -3299
rect 872 -3367 906 -3333
rect 872 -3435 906 -3401
rect 872 -3503 906 -3469
rect 872 -3571 906 -3537
rect 872 -3639 906 -3605
rect 872 -3707 906 -3673
rect 5231 -3367 5265 -3333
rect 5231 -3435 5265 -3401
rect 5231 -3503 5265 -3469
rect 5231 -3571 5265 -3537
rect 5231 -3639 5265 -3605
rect 5231 -3707 5265 -3673
rect 9589 -3367 9623 -3333
rect 9589 -3435 9623 -3401
rect 9589 -3503 9623 -3469
rect 9589 -3571 9623 -3537
rect 9589 -3639 9623 -3605
rect 872 -3775 906 -3741
rect 872 -3843 906 -3809
rect 9589 -3707 9623 -3673
rect 5231 -3775 5265 -3741
rect 5231 -3843 5265 -3809
rect 9589 -3775 9623 -3741
rect 9589 -3843 9623 -3809
rect 993 -4106 1027 -4072
rect 1061 -4106 1095 -4072
rect 1129 -4106 1163 -4072
rect 1197 -4106 1231 -4072
rect 1265 -4106 1299 -4072
rect 1333 -4106 1367 -4072
rect 1401 -4106 1435 -4072
rect 1469 -4106 1503 -4072
rect 1537 -4106 1571 -4072
rect 1605 -4106 1639 -4072
rect 1673 -4106 1707 -4072
rect 1741 -4106 1775 -4072
rect 1809 -4106 1843 -4072
rect 1877 -4106 1911 -4072
rect 1945 -4106 1979 -4072
rect 2013 -4106 2047 -4072
rect 2081 -4106 2115 -4072
rect 2149 -4106 2183 -4072
rect 2217 -4106 2251 -4072
rect 2285 -4106 2319 -4072
rect 2353 -4106 2387 -4072
rect 2421 -4106 2455 -4072
rect 2489 -4106 2523 -4072
rect 2557 -4106 2591 -4072
rect 2625 -4106 2659 -4072
rect 2693 -4106 2727 -4072
rect 2761 -4106 2795 -4072
rect 2829 -4106 2863 -4072
rect 2897 -4106 2931 -4072
rect 2965 -4106 2999 -4072
rect 3033 -4106 3067 -4072
rect 3101 -4106 3135 -4072
rect 3169 -4106 3203 -4072
rect 3237 -4106 3271 -4072
rect 3305 -4106 3339 -4072
rect 3373 -4106 3407 -4072
rect 3441 -4106 3475 -4072
rect 3509 -4106 3543 -4072
rect 3577 -4106 3611 -4072
rect 3645 -4106 3679 -4072
rect 3713 -4106 3747 -4072
rect 3781 -4106 3815 -4072
rect 3849 -4106 3883 -4072
rect 3917 -4106 3951 -4072
rect 3985 -4106 4019 -4072
rect 4053 -4106 4087 -4072
rect 4121 -4106 4155 -4072
rect 4189 -4106 4223 -4072
rect 4257 -4106 4291 -4072
rect 4325 -4106 4359 -4072
rect 4393 -4106 4427 -4072
rect 4461 -4106 4495 -4072
rect 4529 -4106 4563 -4072
rect 4597 -4106 4631 -4072
rect 4665 -4106 4699 -4072
rect 4733 -4106 4767 -4072
rect 4801 -4106 4835 -4072
rect 4869 -4106 4903 -4072
rect 4937 -4106 4971 -4072
rect 5005 -4106 5039 -4072
rect 5073 -4106 5107 -4072
rect 5388 -4106 5422 -4072
rect 5456 -4106 5490 -4072
rect 5524 -4106 5558 -4072
rect 5592 -4106 5626 -4072
rect 5660 -4106 5694 -4072
rect 5728 -4106 5762 -4072
rect 5796 -4106 5830 -4072
rect 5864 -4106 5898 -4072
rect 5932 -4106 5966 -4072
rect 6000 -4106 6034 -4072
rect 6068 -4106 6102 -4072
rect 6136 -4106 6170 -4072
rect 6204 -4106 6238 -4072
rect 6272 -4106 6306 -4072
rect 6340 -4106 6374 -4072
rect 6408 -4106 6442 -4072
rect 6476 -4106 6510 -4072
rect 6544 -4106 6578 -4072
rect 6612 -4106 6646 -4072
rect 6680 -4106 6714 -4072
rect 6748 -4106 6782 -4072
rect 6816 -4106 6850 -4072
rect 6884 -4106 6918 -4072
rect 6952 -4106 6986 -4072
rect 7020 -4106 7054 -4072
rect 7088 -4106 7122 -4072
rect 7156 -4106 7190 -4072
rect 7224 -4106 7258 -4072
rect 7292 -4106 7326 -4072
rect 7360 -4106 7394 -4072
rect 7428 -4106 7462 -4072
rect 7496 -4106 7530 -4072
rect 7564 -4106 7598 -4072
rect 7632 -4106 7666 -4072
rect 7700 -4106 7734 -4072
rect 7768 -4106 7802 -4072
rect 7836 -4106 7870 -4072
rect 7904 -4106 7938 -4072
rect 7972 -4106 8006 -4072
rect 8040 -4106 8074 -4072
rect 8108 -4106 8142 -4072
rect 8176 -4106 8210 -4072
rect 8244 -4106 8278 -4072
rect 8312 -4106 8346 -4072
rect 8380 -4106 8414 -4072
rect 8448 -4106 8482 -4072
rect 8516 -4106 8550 -4072
rect 8584 -4106 8618 -4072
rect 8652 -4106 8686 -4072
rect 8720 -4106 8754 -4072
rect 8788 -4106 8822 -4072
rect 8856 -4106 8890 -4072
rect 8924 -4106 8958 -4072
rect 8992 -4106 9026 -4072
rect 9060 -4106 9094 -4072
rect 9128 -4106 9162 -4072
rect 9196 -4106 9230 -4072
rect 9264 -4106 9298 -4072
rect 9332 -4106 9366 -4072
rect 9400 -4106 9434 -4072
rect 9468 -4106 9502 -4072
rect 872 -4369 906 -4335
rect 872 -4437 906 -4403
rect 5231 -4369 5265 -4335
rect 5231 -4437 5265 -4403
rect 872 -4505 906 -4471
rect 9589 -4369 9623 -4335
rect 9589 -4437 9623 -4403
rect 872 -4573 906 -4539
rect 872 -4641 906 -4607
rect 872 -4709 906 -4675
rect 872 -4777 906 -4743
rect 872 -4845 906 -4811
rect 5231 -4505 5265 -4471
rect 5231 -4573 5265 -4539
rect 5231 -4641 5265 -4607
rect 5231 -4709 5265 -4675
rect 5231 -4777 5265 -4743
rect 5231 -4845 5265 -4811
rect 9589 -4505 9623 -4471
rect 9589 -4573 9623 -4539
rect 9589 -4641 9623 -4607
rect 9589 -4709 9623 -4675
rect 9589 -4777 9623 -4743
rect 9589 -4845 9623 -4811
rect 993 -4879 1027 -4845
rect 1061 -4879 1095 -4845
rect 1129 -4879 1163 -4845
rect 1197 -4879 1231 -4845
rect 1265 -4879 1299 -4845
rect 1333 -4879 1367 -4845
rect 1401 -4879 1435 -4845
rect 1469 -4879 1503 -4845
rect 1537 -4879 1571 -4845
rect 1605 -4879 1639 -4845
rect 1673 -4879 1707 -4845
rect 1741 -4879 1775 -4845
rect 1809 -4879 1843 -4845
rect 1877 -4879 1911 -4845
rect 1945 -4879 1979 -4845
rect 2013 -4879 2047 -4845
rect 2081 -4879 2115 -4845
rect 2149 -4879 2183 -4845
rect 2217 -4879 2251 -4845
rect 2285 -4879 2319 -4845
rect 2353 -4879 2387 -4845
rect 2421 -4879 2455 -4845
rect 2489 -4879 2523 -4845
rect 2557 -4879 2591 -4845
rect 2625 -4879 2659 -4845
rect 2693 -4879 2727 -4845
rect 2761 -4879 2795 -4845
rect 2829 -4879 2863 -4845
rect 2897 -4879 2931 -4845
rect 2965 -4879 2999 -4845
rect 3033 -4879 3067 -4845
rect 3101 -4879 3135 -4845
rect 3169 -4879 3203 -4845
rect 3237 -4879 3271 -4845
rect 3305 -4879 3339 -4845
rect 3373 -4879 3407 -4845
rect 3441 -4879 3475 -4845
rect 3509 -4879 3543 -4845
rect 3577 -4879 3611 -4845
rect 3645 -4879 3679 -4845
rect 3713 -4879 3747 -4845
rect 3781 -4879 3815 -4845
rect 3849 -4879 3883 -4845
rect 3917 -4879 3951 -4845
rect 3985 -4879 4019 -4845
rect 4053 -4879 4087 -4845
rect 4121 -4879 4155 -4845
rect 4189 -4879 4223 -4845
rect 4257 -4879 4291 -4845
rect 4325 -4879 4359 -4845
rect 4393 -4879 4427 -4845
rect 4461 -4879 4495 -4845
rect 4529 -4879 4563 -4845
rect 4597 -4879 4631 -4845
rect 4665 -4879 4699 -4845
rect 4733 -4879 4767 -4845
rect 4801 -4879 4835 -4845
rect 4869 -4879 4903 -4845
rect 4937 -4879 4971 -4845
rect 5005 -4879 5039 -4845
rect 5073 -4879 5107 -4845
rect 5388 -4879 5422 -4845
rect 5456 -4879 5490 -4845
rect 5524 -4879 5558 -4845
rect 5592 -4879 5626 -4845
rect 5660 -4879 5694 -4845
rect 5728 -4879 5762 -4845
rect 5796 -4879 5830 -4845
rect 5864 -4879 5898 -4845
rect 5932 -4879 5966 -4845
rect 6000 -4879 6034 -4845
rect 6068 -4879 6102 -4845
rect 6136 -4879 6170 -4845
rect 6204 -4879 6238 -4845
rect 6272 -4879 6306 -4845
rect 6340 -4879 6374 -4845
rect 6408 -4879 6442 -4845
rect 6476 -4879 6510 -4845
rect 6544 -4879 6578 -4845
rect 6612 -4879 6646 -4845
rect 6680 -4879 6714 -4845
rect 6748 -4879 6782 -4845
rect 6816 -4879 6850 -4845
rect 6884 -4879 6918 -4845
rect 6952 -4879 6986 -4845
rect 7020 -4879 7054 -4845
rect 7088 -4879 7122 -4845
rect 7156 -4879 7190 -4845
rect 7224 -4879 7258 -4845
rect 7292 -4879 7326 -4845
rect 7360 -4879 7394 -4845
rect 7428 -4879 7462 -4845
rect 7496 -4879 7530 -4845
rect 7564 -4879 7598 -4845
rect 7632 -4879 7666 -4845
rect 7700 -4879 7734 -4845
rect 7768 -4879 7802 -4845
rect 7836 -4879 7870 -4845
rect 7904 -4879 7938 -4845
rect 7972 -4879 8006 -4845
rect 8040 -4879 8074 -4845
rect 8108 -4879 8142 -4845
rect 8176 -4879 8210 -4845
rect 8244 -4879 8278 -4845
rect 8312 -4879 8346 -4845
rect 8380 -4879 8414 -4845
rect 8448 -4879 8482 -4845
rect 8516 -4879 8550 -4845
rect 8584 -4879 8618 -4845
rect 8652 -4879 8686 -4845
rect 8720 -4879 8754 -4845
rect 8788 -4879 8822 -4845
rect 8856 -4879 8890 -4845
rect 8924 -4879 8958 -4845
rect 8992 -4879 9026 -4845
rect 9060 -4879 9094 -4845
rect 9128 -4879 9162 -4845
rect 9196 -4879 9230 -4845
rect 9264 -4879 9298 -4845
rect 9332 -4879 9366 -4845
rect 9400 -4879 9434 -4845
rect 9468 -4879 9502 -4845
rect 872 -4913 906 -4879
rect 872 -4981 906 -4947
rect 872 -5049 906 -5015
rect 872 -5117 906 -5083
rect 872 -5185 906 -5151
rect 872 -5253 906 -5219
rect 5231 -4913 5265 -4879
rect 5231 -4981 5265 -4947
rect 5231 -5049 5265 -5015
rect 5231 -5117 5265 -5083
rect 5231 -5185 5265 -5151
rect 5231 -5253 5265 -5219
rect 9589 -4913 9623 -4879
rect 9589 -4981 9623 -4947
rect 9589 -5049 9623 -5015
rect 9589 -5117 9623 -5083
rect 9589 -5185 9623 -5151
rect 872 -5321 906 -5287
rect 872 -5389 906 -5355
rect 872 -5457 906 -5423
rect 9589 -5253 9623 -5219
rect 5231 -5321 5265 -5287
rect 5231 -5389 5265 -5355
rect 5231 -5457 5265 -5423
rect 9589 -5321 9623 -5287
rect 9589 -5389 9623 -5355
rect 9589 -5457 9623 -5423
rect 872 -5525 906 -5491
rect 5231 -5525 5265 -5491
rect 872 -5593 906 -5559
rect 872 -5661 906 -5627
rect 872 -5729 906 -5695
rect 872 -5797 906 -5763
rect 872 -5865 906 -5831
rect 9589 -5525 9623 -5491
rect 5231 -5593 5265 -5559
rect 5231 -5661 5265 -5627
rect 5231 -5729 5265 -5695
rect 5231 -5797 5265 -5763
rect 872 -5933 906 -5899
rect 5231 -5865 5265 -5831
rect 9589 -5593 9623 -5559
rect 9589 -5661 9623 -5627
rect 9589 -5729 9623 -5695
rect 9589 -5797 9623 -5763
rect 5231 -5933 5265 -5899
rect 872 -6001 906 -5967
rect 872 -6069 906 -6035
rect 872 -6137 906 -6103
rect 9589 -5865 9623 -5831
rect 9589 -5933 9623 -5899
rect 5231 -6001 5265 -5967
rect 5231 -6069 5265 -6035
rect 5231 -6137 5265 -6103
rect 872 -6205 906 -6171
rect 9589 -6001 9623 -5967
rect 9589 -6069 9623 -6035
rect 9589 -6137 9623 -6103
rect 872 -6273 906 -6239
rect 872 -6341 906 -6307
rect 872 -6409 906 -6375
rect 5231 -6205 5265 -6171
rect 5231 -6273 5265 -6239
rect 5231 -6341 5265 -6307
rect 5231 -6409 5265 -6375
rect 9589 -6205 9623 -6171
rect 9589 -6273 9623 -6239
rect 9589 -6341 9623 -6307
rect 9589 -6409 9623 -6375
rect 993 -6545 1027 -6511
rect 1061 -6545 1095 -6511
rect 1129 -6545 1163 -6511
rect 1197 -6545 1231 -6511
rect 1265 -6545 1299 -6511
rect 1333 -6545 1367 -6511
rect 1401 -6545 1435 -6511
rect 1469 -6545 1503 -6511
rect 1537 -6545 1571 -6511
rect 1605 -6545 1639 -6511
rect 1673 -6545 1707 -6511
rect 1741 -6545 1775 -6511
rect 1809 -6545 1843 -6511
rect 1877 -6545 1911 -6511
rect 1945 -6545 1979 -6511
rect 2013 -6545 2047 -6511
rect 2081 -6545 2115 -6511
rect 2149 -6545 2183 -6511
rect 2217 -6545 2251 -6511
rect 2285 -6545 2319 -6511
rect 2353 -6545 2387 -6511
rect 2421 -6545 2455 -6511
rect 2489 -6545 2523 -6511
rect 2557 -6545 2591 -6511
rect 2625 -6545 2659 -6511
rect 2693 -6545 2727 -6511
rect 2761 -6545 2795 -6511
rect 2829 -6545 2863 -6511
rect 2897 -6545 2931 -6511
rect 2965 -6545 2999 -6511
rect 3033 -6545 3067 -6511
rect 3101 -6545 3135 -6511
rect 3169 -6545 3203 -6511
rect 3237 -6545 3271 -6511
rect 3305 -6545 3339 -6511
rect 3373 -6545 3407 -6511
rect 3441 -6545 3475 -6511
rect 3509 -6545 3543 -6511
rect 3577 -6545 3611 -6511
rect 3645 -6545 3679 -6511
rect 3713 -6545 3747 -6511
rect 3781 -6545 3815 -6511
rect 3849 -6545 3883 -6511
rect 3917 -6545 3951 -6511
rect 3985 -6545 4019 -6511
rect 4053 -6545 4087 -6511
rect 4121 -6545 4155 -6511
rect 4189 -6545 4223 -6511
rect 4257 -6545 4291 -6511
rect 4325 -6545 4359 -6511
rect 4393 -6545 4427 -6511
rect 4461 -6545 4495 -6511
rect 4529 -6545 4563 -6511
rect 4597 -6545 4631 -6511
rect 4665 -6545 4699 -6511
rect 4733 -6545 4767 -6511
rect 4801 -6545 4835 -6511
rect 4869 -6545 4903 -6511
rect 4937 -6545 4971 -6511
rect 5005 -6545 5039 -6511
rect 5073 -6545 5107 -6511
rect 5388 -6545 5422 -6511
rect 5456 -6545 5490 -6511
rect 5524 -6545 5558 -6511
rect 5592 -6545 5626 -6511
rect 5660 -6545 5694 -6511
rect 5728 -6545 5762 -6511
rect 5796 -6545 5830 -6511
rect 5864 -6545 5898 -6511
rect 5932 -6545 5966 -6511
rect 6000 -6545 6034 -6511
rect 6068 -6545 6102 -6511
rect 6136 -6545 6170 -6511
rect 6204 -6545 6238 -6511
rect 6272 -6545 6306 -6511
rect 6340 -6545 6374 -6511
rect 6408 -6545 6442 -6511
rect 6476 -6545 6510 -6511
rect 6544 -6545 6578 -6511
rect 6612 -6545 6646 -6511
rect 6680 -6545 6714 -6511
rect 6748 -6545 6782 -6511
rect 6816 -6545 6850 -6511
rect 6884 -6545 6918 -6511
rect 6952 -6545 6986 -6511
rect 7020 -6545 7054 -6511
rect 7088 -6545 7122 -6511
rect 7156 -6545 7190 -6511
rect 7224 -6545 7258 -6511
rect 7292 -6545 7326 -6511
rect 7360 -6545 7394 -6511
rect 7428 -6545 7462 -6511
rect 7496 -6545 7530 -6511
rect 7564 -6545 7598 -6511
rect 7632 -6545 7666 -6511
rect 7700 -6545 7734 -6511
rect 7768 -6545 7802 -6511
rect 7836 -6545 7870 -6511
rect 7904 -6545 7938 -6511
rect 7972 -6545 8006 -6511
rect 8040 -6545 8074 -6511
rect 8108 -6545 8142 -6511
rect 8176 -6545 8210 -6511
rect 8244 -6545 8278 -6511
rect 8312 -6545 8346 -6511
rect 8380 -6545 8414 -6511
rect 8448 -6545 8482 -6511
rect 8516 -6545 8550 -6511
rect 8584 -6545 8618 -6511
rect 8652 -6545 8686 -6511
rect 8720 -6545 8754 -6511
rect 8788 -6545 8822 -6511
rect 8856 -6545 8890 -6511
rect 8924 -6545 8958 -6511
rect 8992 -6545 9026 -6511
rect 9060 -6545 9094 -6511
rect 9128 -6545 9162 -6511
rect 9196 -6545 9230 -6511
rect 9264 -6545 9298 -6511
rect 9332 -6545 9366 -6511
rect 9400 -6545 9434 -6511
rect 9468 -6545 9502 -6511
rect 872 -6681 906 -6647
rect 872 -6749 906 -6715
rect 872 -6817 906 -6783
rect 872 -6885 906 -6851
rect 5231 -6681 5265 -6647
rect 5231 -6749 5265 -6715
rect 5231 -6817 5265 -6783
rect 5231 -6885 5265 -6851
rect 9589 -6681 9623 -6647
rect 9589 -6749 9623 -6715
rect 9589 -6817 9623 -6783
rect 872 -6953 906 -6919
rect 872 -7021 906 -6987
rect 872 -7089 906 -7055
rect 9589 -6885 9623 -6851
rect 5231 -6953 5265 -6919
rect 5231 -7021 5265 -6987
rect 5231 -7089 5265 -7055
rect 872 -7157 906 -7123
rect 872 -7225 906 -7191
rect 9589 -6953 9623 -6919
rect 9589 -7021 9623 -6987
rect 9589 -7089 9623 -7055
rect 5231 -7157 5265 -7123
rect 872 -7293 906 -7259
rect 872 -7361 906 -7327
rect 872 -7429 906 -7395
rect 872 -7497 906 -7463
rect 5231 -7225 5265 -7191
rect 9589 -7157 9623 -7123
rect 5231 -7293 5265 -7259
rect 5231 -7361 5265 -7327
rect 5231 -7429 5265 -7395
rect 5231 -7497 5265 -7463
rect 9589 -7225 9623 -7191
rect 9589 -7293 9623 -7259
rect 9589 -7361 9623 -7327
rect 9589 -7429 9623 -7395
rect 9589 -7497 9623 -7463
rect 872 -7565 906 -7531
rect 5231 -7565 5265 -7531
rect 872 -7633 906 -7599
rect 872 -7701 906 -7667
rect 872 -7769 906 -7735
rect 9589 -7565 9623 -7531
rect 5231 -7633 5265 -7599
rect 5231 -7701 5265 -7667
rect 5231 -7769 5265 -7735
rect 872 -7837 906 -7803
rect 9589 -7633 9623 -7599
rect 9589 -7701 9623 -7667
rect 9589 -7769 9623 -7735
rect 872 -7905 906 -7871
rect 872 -7973 906 -7939
rect 872 -8041 906 -8007
rect 872 -8109 906 -8075
rect 5231 -7837 5265 -7803
rect 5231 -7905 5265 -7871
rect 5231 -7973 5265 -7939
rect 5231 -8041 5265 -8007
rect 5231 -8109 5265 -8075
rect 9589 -7837 9623 -7803
rect 9589 -7905 9623 -7871
rect 9589 -7973 9623 -7939
rect 9589 -8041 9623 -8007
rect 9589 -8109 9623 -8075
rect 993 -8143 1027 -8109
rect 1061 -8143 1095 -8109
rect 1129 -8143 1163 -8109
rect 1197 -8143 1231 -8109
rect 1265 -8143 1299 -8109
rect 1333 -8143 1367 -8109
rect 1401 -8143 1435 -8109
rect 1469 -8143 1503 -8109
rect 1537 -8143 1571 -8109
rect 1605 -8143 1639 -8109
rect 1673 -8143 1707 -8109
rect 1741 -8143 1775 -8109
rect 1809 -8143 1843 -8109
rect 1877 -8143 1911 -8109
rect 1945 -8143 1979 -8109
rect 2013 -8143 2047 -8109
rect 2081 -8143 2115 -8109
rect 2149 -8143 2183 -8109
rect 2217 -8143 2251 -8109
rect 2285 -8143 2319 -8109
rect 2353 -8143 2387 -8109
rect 2421 -8143 2455 -8109
rect 2489 -8143 2523 -8109
rect 2557 -8143 2591 -8109
rect 2625 -8143 2659 -8109
rect 2693 -8143 2727 -8109
rect 2761 -8143 2795 -8109
rect 2829 -8143 2863 -8109
rect 2897 -8143 2931 -8109
rect 2965 -8143 2999 -8109
rect 3033 -8143 3067 -8109
rect 3101 -8143 3135 -8109
rect 3169 -8143 3203 -8109
rect 3237 -8143 3271 -8109
rect 3305 -8143 3339 -8109
rect 3373 -8143 3407 -8109
rect 3441 -8143 3475 -8109
rect 3509 -8143 3543 -8109
rect 3577 -8143 3611 -8109
rect 3645 -8143 3679 -8109
rect 3713 -8143 3747 -8109
rect 3781 -8143 3815 -8109
rect 3849 -8143 3883 -8109
rect 3917 -8143 3951 -8109
rect 3985 -8143 4019 -8109
rect 4053 -8143 4087 -8109
rect 4121 -8143 4155 -8109
rect 4189 -8143 4223 -8109
rect 4257 -8143 4291 -8109
rect 4325 -8143 4359 -8109
rect 4393 -8143 4427 -8109
rect 4461 -8143 4495 -8109
rect 4529 -8143 4563 -8109
rect 4597 -8143 4631 -8109
rect 4665 -8143 4699 -8109
rect 4733 -8143 4767 -8109
rect 4801 -8143 4835 -8109
rect 4869 -8143 4903 -8109
rect 4937 -8143 4971 -8109
rect 5005 -8143 5039 -8109
rect 5073 -8143 5107 -8109
rect 5388 -8143 5422 -8109
rect 5456 -8143 5490 -8109
rect 5524 -8143 5558 -8109
rect 5592 -8143 5626 -8109
rect 5660 -8143 5694 -8109
rect 5728 -8143 5762 -8109
rect 5796 -8143 5830 -8109
rect 5864 -8143 5898 -8109
rect 5932 -8143 5966 -8109
rect 6000 -8143 6034 -8109
rect 6068 -8143 6102 -8109
rect 6136 -8143 6170 -8109
rect 6204 -8143 6238 -8109
rect 6272 -8143 6306 -8109
rect 6340 -8143 6374 -8109
rect 6408 -8143 6442 -8109
rect 6476 -8143 6510 -8109
rect 6544 -8143 6578 -8109
rect 6612 -8143 6646 -8109
rect 6680 -8143 6714 -8109
rect 6748 -8143 6782 -8109
rect 6816 -8143 6850 -8109
rect 6884 -8143 6918 -8109
rect 6952 -8143 6986 -8109
rect 7020 -8143 7054 -8109
rect 7088 -8143 7122 -8109
rect 7156 -8143 7190 -8109
rect 7224 -8143 7258 -8109
rect 7292 -8143 7326 -8109
rect 7360 -8143 7394 -8109
rect 7428 -8143 7462 -8109
rect 7496 -8143 7530 -8109
rect 7564 -8143 7598 -8109
rect 7632 -8143 7666 -8109
rect 7700 -8143 7734 -8109
rect 7768 -8143 7802 -8109
rect 7836 -8143 7870 -8109
rect 7904 -8143 7938 -8109
rect 7972 -8143 8006 -8109
rect 8040 -8143 8074 -8109
rect 8108 -8143 8142 -8109
rect 8176 -8143 8210 -8109
rect 8244 -8143 8278 -8109
rect 8312 -8143 8346 -8109
rect 8380 -8143 8414 -8109
rect 8448 -8143 8482 -8109
rect 8516 -8143 8550 -8109
rect 8584 -8143 8618 -8109
rect 8652 -8143 8686 -8109
rect 8720 -8143 8754 -8109
rect 8788 -8143 8822 -8109
rect 8856 -8143 8890 -8109
rect 8924 -8143 8958 -8109
rect 8992 -8143 9026 -8109
rect 9060 -8143 9094 -8109
rect 9128 -8143 9162 -8109
rect 9196 -8143 9230 -8109
rect 9264 -8143 9298 -8109
rect 9332 -8143 9366 -8109
rect 9400 -8143 9434 -8109
rect 9468 -8143 9502 -8109
rect 872 -8177 906 -8143
rect 872 -8245 906 -8211
rect 872 -8313 906 -8279
rect 872 -8381 906 -8347
rect 872 -8449 906 -8415
rect 872 -8517 906 -8483
rect 5231 -8177 5265 -8143
rect 5231 -8245 5265 -8211
rect 5231 -8313 5265 -8279
rect 5231 -8381 5265 -8347
rect 5231 -8449 5265 -8415
rect 5231 -8517 5265 -8483
rect 9589 -8177 9623 -8143
rect 9589 -8245 9623 -8211
rect 9589 -8313 9623 -8279
rect 9589 -8381 9623 -8347
rect 9589 -8449 9623 -8415
rect 872 -8585 906 -8551
rect 872 -8653 906 -8619
rect 872 -8721 906 -8687
rect 9589 -8517 9623 -8483
rect 5231 -8585 5265 -8551
rect 5231 -8653 5265 -8619
rect 5231 -8721 5265 -8687
rect 9589 -8585 9623 -8551
rect 9589 -8653 9623 -8619
rect 9589 -8721 9623 -8687
rect 993 -8933 1027 -8899
rect 1061 -8933 1095 -8899
rect 1129 -8933 1163 -8899
rect 1197 -8933 1231 -8899
rect 1265 -8933 1299 -8899
rect 1333 -8933 1367 -8899
rect 1401 -8933 1435 -8899
rect 1469 -8933 1503 -8899
rect 1537 -8933 1571 -8899
rect 1605 -8933 1639 -8899
rect 1673 -8933 1707 -8899
rect 1741 -8933 1775 -8899
rect 1809 -8933 1843 -8899
rect 1877 -8933 1911 -8899
rect 1945 -8933 1979 -8899
rect 2013 -8933 2047 -8899
rect 2081 -8933 2115 -8899
rect 2149 -8933 2183 -8899
rect 2217 -8933 2251 -8899
rect 2285 -8933 2319 -8899
rect 2353 -8933 2387 -8899
rect 2421 -8933 2455 -8899
rect 2489 -8933 2523 -8899
rect 2557 -8933 2591 -8899
rect 2625 -8933 2659 -8899
rect 2693 -8933 2727 -8899
rect 2761 -8933 2795 -8899
rect 2829 -8933 2863 -8899
rect 2897 -8933 2931 -8899
rect 2965 -8933 2999 -8899
rect 3033 -8933 3067 -8899
rect 3101 -8933 3135 -8899
rect 3169 -8933 3203 -8899
rect 3237 -8933 3271 -8899
rect 3305 -8933 3339 -8899
rect 3373 -8933 3407 -8899
rect 3441 -8933 3475 -8899
rect 3509 -8933 3543 -8899
rect 3577 -8933 3611 -8899
rect 3645 -8933 3679 -8899
rect 3713 -8933 3747 -8899
rect 3781 -8933 3815 -8899
rect 3849 -8933 3883 -8899
rect 3917 -8933 3951 -8899
rect 3985 -8933 4019 -8899
rect 4053 -8933 4087 -8899
rect 4121 -8933 4155 -8899
rect 4189 -8933 4223 -8899
rect 4257 -8933 4291 -8899
rect 4325 -8933 4359 -8899
rect 4393 -8933 4427 -8899
rect 4461 -8933 4495 -8899
rect 4529 -8933 4563 -8899
rect 4597 -8933 4631 -8899
rect 4665 -8933 4699 -8899
rect 4733 -8933 4767 -8899
rect 4801 -8933 4835 -8899
rect 4869 -8933 4903 -8899
rect 4937 -8933 4971 -8899
rect 5005 -8933 5039 -8899
rect 5073 -8933 5107 -8899
rect 5388 -8933 5422 -8899
rect 5456 -8933 5490 -8899
rect 5524 -8933 5558 -8899
rect 5592 -8933 5626 -8899
rect 5660 -8933 5694 -8899
rect 5728 -8933 5762 -8899
rect 5796 -8933 5830 -8899
rect 5864 -8933 5898 -8899
rect 5932 -8933 5966 -8899
rect 6000 -8933 6034 -8899
rect 6068 -8933 6102 -8899
rect 6136 -8933 6170 -8899
rect 6204 -8933 6238 -8899
rect 6272 -8933 6306 -8899
rect 6340 -8933 6374 -8899
rect 6408 -8933 6442 -8899
rect 6476 -8933 6510 -8899
rect 6544 -8933 6578 -8899
rect 6612 -8933 6646 -8899
rect 6680 -8933 6714 -8899
rect 6748 -8933 6782 -8899
rect 6816 -8933 6850 -8899
rect 6884 -8933 6918 -8899
rect 6952 -8933 6986 -8899
rect 7020 -8933 7054 -8899
rect 7088 -8933 7122 -8899
rect 7156 -8933 7190 -8899
rect 7224 -8933 7258 -8899
rect 7292 -8933 7326 -8899
rect 7360 -8933 7394 -8899
rect 7428 -8933 7462 -8899
rect 7496 -8933 7530 -8899
rect 7564 -8933 7598 -8899
rect 7632 -8933 7666 -8899
rect 7700 -8933 7734 -8899
rect 7768 -8933 7802 -8899
rect 7836 -8933 7870 -8899
rect 7904 -8933 7938 -8899
rect 7972 -8933 8006 -8899
rect 8040 -8933 8074 -8899
rect 8108 -8933 8142 -8899
rect 8176 -8933 8210 -8899
rect 8244 -8933 8278 -8899
rect 8312 -8933 8346 -8899
rect 8380 -8933 8414 -8899
rect 8448 -8933 8482 -8899
rect 8516 -8933 8550 -8899
rect 8584 -8933 8618 -8899
rect 8652 -8933 8686 -8899
rect 8720 -8933 8754 -8899
rect 8788 -8933 8822 -8899
rect 8856 -8933 8890 -8899
rect 8924 -8933 8958 -8899
rect 8992 -8933 9026 -8899
rect 9060 -8933 9094 -8899
rect 9128 -8933 9162 -8899
rect 9196 -8933 9230 -8899
rect 9264 -8933 9298 -8899
rect 9332 -8933 9366 -8899
rect 9400 -8933 9434 -8899
rect 9468 -8933 9502 -8899
<< poly >>
rect 1033 642 1233 658
rect 1033 608 1082 642
rect 1116 608 1150 642
rect 1184 608 1233 642
rect 1033 561 1233 608
rect 1485 642 1685 658
rect 1485 608 1534 642
rect 1568 608 1602 642
rect 1636 608 1685 642
rect 1485 561 1685 608
rect 1743 642 1943 658
rect 1743 608 1792 642
rect 1826 608 1860 642
rect 1894 608 1943 642
rect 1743 561 1943 608
rect 2001 642 2201 658
rect 2001 608 2050 642
rect 2084 608 2118 642
rect 2152 608 2201 642
rect 2001 561 2201 608
rect 2259 642 2459 658
rect 2259 608 2308 642
rect 2342 608 2376 642
rect 2410 608 2459 642
rect 2259 561 2459 608
rect 2711 642 2911 658
rect 2711 608 2760 642
rect 2794 608 2828 642
rect 2862 608 2911 642
rect 2711 561 2911 608
rect 2969 642 3169 658
rect 2969 608 3018 642
rect 3052 608 3086 642
rect 3120 608 3169 642
rect 2969 561 3169 608
rect 3227 642 3427 658
rect 3227 608 3276 642
rect 3310 608 3344 642
rect 3378 608 3427 642
rect 3227 561 3427 608
rect 3679 642 3879 658
rect 3679 608 3728 642
rect 3762 608 3796 642
rect 3830 608 3879 642
rect 3679 561 3879 608
rect 3937 642 4137 658
rect 3937 608 3986 642
rect 4020 608 4054 642
rect 4088 608 4137 642
rect 3937 561 4137 608
rect 4195 642 4395 658
rect 4195 608 4244 642
rect 4278 608 4312 642
rect 4346 608 4395 642
rect 4195 561 4395 608
rect 4453 642 4653 658
rect 4453 608 4502 642
rect 4536 608 4570 642
rect 4604 608 4653 642
rect 4453 561 4653 608
rect 4905 642 5105 658
rect 4905 608 4954 642
rect 4988 608 5022 642
rect 5056 608 5105 642
rect 4905 561 5105 608
rect 5391 642 5591 658
rect 5391 608 5440 642
rect 5474 608 5508 642
rect 5542 608 5591 642
rect 5391 561 5591 608
rect 5842 642 6042 658
rect 5842 608 5891 642
rect 5925 608 5959 642
rect 5993 608 6042 642
rect 5842 561 6042 608
rect 6100 642 6300 658
rect 6100 608 6149 642
rect 6183 608 6217 642
rect 6251 608 6300 642
rect 6100 561 6300 608
rect 6358 642 6558 658
rect 6358 608 6407 642
rect 6441 608 6475 642
rect 6509 608 6558 642
rect 6358 561 6558 608
rect 6616 642 6816 658
rect 6616 608 6665 642
rect 6699 608 6733 642
rect 6767 608 6816 642
rect 6616 561 6816 608
rect 7068 642 7268 658
rect 7068 608 7117 642
rect 7151 608 7185 642
rect 7219 608 7268 642
rect 7068 561 7268 608
rect 7326 642 7526 658
rect 7326 608 7375 642
rect 7409 608 7443 642
rect 7477 608 7526 642
rect 7326 561 7526 608
rect 7584 642 7784 658
rect 7584 608 7633 642
rect 7667 608 7701 642
rect 7735 608 7784 642
rect 7584 561 7784 608
rect 8036 642 8236 658
rect 8036 608 8085 642
rect 8119 608 8153 642
rect 8187 608 8236 642
rect 8036 561 8236 608
rect 8294 642 8494 658
rect 8294 608 8343 642
rect 8377 608 8411 642
rect 8445 608 8494 642
rect 8294 561 8494 608
rect 8552 642 8752 658
rect 8552 608 8601 642
rect 8635 608 8669 642
rect 8703 608 8752 642
rect 8552 561 8752 608
rect 8810 642 9010 658
rect 8810 608 8859 642
rect 8893 608 8927 642
rect 8961 608 9010 642
rect 8810 561 9010 608
rect 9262 642 9462 658
rect 9262 608 9311 642
rect 9345 608 9379 642
rect 9413 608 9462 642
rect 9262 561 9462 608
rect 1033 335 1233 361
rect 1485 335 1685 361
rect 1743 335 1943 361
rect 2001 335 2201 361
rect 2259 335 2459 361
rect 2711 335 2911 361
rect 2969 335 3169 361
rect 3227 335 3427 361
rect 3679 335 3879 361
rect 3937 335 4137 361
rect 4195 335 4395 361
rect 4453 335 4653 361
rect 4905 335 5105 361
rect 5391 335 5591 361
rect 5842 335 6042 361
rect 6100 335 6300 361
rect 6358 335 6558 361
rect 6616 335 6816 361
rect 7068 335 7268 361
rect 7326 335 7526 361
rect 7584 335 7784 361
rect 8036 335 8236 361
rect 8294 335 8494 361
rect 8552 335 8752 361
rect 8810 335 9010 361
rect 9262 335 9462 361
rect 1033 -383 1233 -357
rect 1485 -383 1685 -357
rect 1743 -383 1943 -357
rect 2001 -383 2201 -357
rect 2259 -383 2459 -357
rect 2711 -383 2911 -357
rect 2969 -383 3169 -357
rect 3227 -383 3427 -357
rect 3679 -383 3879 -357
rect 3937 -383 4137 -357
rect 4195 -383 4395 -357
rect 4453 -383 4653 -357
rect 4905 -383 5105 -357
rect 5391 -383 5591 -357
rect 5842 -383 6042 -357
rect 6100 -383 6300 -357
rect 6358 -383 6558 -357
rect 6616 -383 6816 -357
rect 7068 -383 7268 -357
rect 7326 -383 7526 -357
rect 7584 -383 7784 -357
rect 8036 -383 8236 -357
rect 8294 -383 8494 -357
rect 8552 -383 8752 -357
rect 8810 -383 9010 -357
rect 9262 -383 9462 -357
rect 1033 -630 1233 -583
rect 1033 -664 1082 -630
rect 1116 -664 1150 -630
rect 1184 -664 1233 -630
rect 1033 -680 1233 -664
rect 1485 -630 1685 -583
rect 1485 -664 1534 -630
rect 1568 -664 1602 -630
rect 1636 -664 1685 -630
rect 1485 -680 1685 -664
rect 1743 -630 1943 -583
rect 1743 -664 1792 -630
rect 1826 -664 1860 -630
rect 1894 -664 1943 -630
rect 1743 -680 1943 -664
rect 2001 -630 2201 -583
rect 2001 -664 2050 -630
rect 2084 -664 2118 -630
rect 2152 -664 2201 -630
rect 2001 -680 2201 -664
rect 2259 -630 2459 -583
rect 2259 -664 2308 -630
rect 2342 -664 2376 -630
rect 2410 -664 2459 -630
rect 2259 -680 2459 -664
rect 2711 -630 2911 -583
rect 2711 -664 2760 -630
rect 2794 -664 2828 -630
rect 2862 -664 2911 -630
rect 2711 -680 2911 -664
rect 2969 -630 3169 -583
rect 2969 -664 3018 -630
rect 3052 -664 3086 -630
rect 3120 -664 3169 -630
rect 2969 -680 3169 -664
rect 3227 -630 3427 -583
rect 3227 -664 3276 -630
rect 3310 -664 3344 -630
rect 3378 -664 3427 -630
rect 3227 -680 3427 -664
rect 3679 -630 3879 -583
rect 3679 -664 3728 -630
rect 3762 -664 3796 -630
rect 3830 -664 3879 -630
rect 3679 -680 3879 -664
rect 3937 -630 4137 -583
rect 3937 -664 3986 -630
rect 4020 -664 4054 -630
rect 4088 -664 4137 -630
rect 3937 -680 4137 -664
rect 4195 -630 4395 -583
rect 4195 -664 4244 -630
rect 4278 -664 4312 -630
rect 4346 -664 4395 -630
rect 4195 -680 4395 -664
rect 4453 -630 4653 -583
rect 4453 -664 4502 -630
rect 4536 -664 4570 -630
rect 4604 -664 4653 -630
rect 4453 -680 4653 -664
rect 4905 -630 5105 -583
rect 4905 -664 4954 -630
rect 4988 -664 5022 -630
rect 5056 -664 5105 -630
rect 4905 -680 5105 -664
rect 5391 -630 5591 -583
rect 5391 -664 5440 -630
rect 5474 -664 5508 -630
rect 5542 -664 5591 -630
rect 5391 -680 5591 -664
rect 5842 -630 6042 -583
rect 5842 -664 5891 -630
rect 5925 -664 5959 -630
rect 5993 -664 6042 -630
rect 5842 -680 6042 -664
rect 6100 -630 6300 -583
rect 6100 -664 6149 -630
rect 6183 -664 6217 -630
rect 6251 -664 6300 -630
rect 6100 -680 6300 -664
rect 6358 -630 6558 -583
rect 6358 -664 6407 -630
rect 6441 -664 6475 -630
rect 6509 -664 6558 -630
rect 6358 -680 6558 -664
rect 6616 -630 6816 -583
rect 6616 -664 6665 -630
rect 6699 -664 6733 -630
rect 6767 -664 6816 -630
rect 6616 -680 6816 -664
rect 7068 -630 7268 -583
rect 7068 -664 7117 -630
rect 7151 -664 7185 -630
rect 7219 -664 7268 -630
rect 7068 -680 7268 -664
rect 7326 -630 7526 -583
rect 7326 -664 7375 -630
rect 7409 -664 7443 -630
rect 7477 -664 7526 -630
rect 7326 -680 7526 -664
rect 7584 -630 7784 -583
rect 7584 -664 7633 -630
rect 7667 -664 7701 -630
rect 7735 -664 7784 -630
rect 7584 -680 7784 -664
rect 8036 -630 8236 -583
rect 8036 -664 8085 -630
rect 8119 -664 8153 -630
rect 8187 -664 8236 -630
rect 8036 -680 8236 -664
rect 8294 -630 8494 -583
rect 8294 -664 8343 -630
rect 8377 -664 8411 -630
rect 8445 -664 8494 -630
rect 8294 -680 8494 -664
rect 8552 -630 8752 -583
rect 8552 -664 8601 -630
rect 8635 -664 8669 -630
rect 8703 -664 8752 -630
rect 8552 -680 8752 -664
rect 8810 -630 9010 -583
rect 8810 -664 8859 -630
rect 8893 -664 8927 -630
rect 8961 -664 9010 -630
rect 8810 -680 9010 -664
rect 9262 -630 9462 -583
rect 9262 -664 9311 -630
rect 9345 -664 9379 -630
rect 9413 -664 9462 -630
rect 9262 -680 9462 -664
rect 1033 -993 1233 -977
rect 1033 -1027 1082 -993
rect 1116 -1027 1150 -993
rect 1184 -1027 1233 -993
rect 1033 -1074 1233 -1027
rect 1485 -993 1685 -977
rect 1485 -1027 1534 -993
rect 1568 -1027 1602 -993
rect 1636 -1027 1685 -993
rect 1485 -1074 1685 -1027
rect 1743 -993 1943 -977
rect 1743 -1027 1792 -993
rect 1826 -1027 1860 -993
rect 1894 -1027 1943 -993
rect 1743 -1074 1943 -1027
rect 2001 -993 2201 -977
rect 2001 -1027 2050 -993
rect 2084 -1027 2118 -993
rect 2152 -1027 2201 -993
rect 2001 -1074 2201 -1027
rect 2259 -993 2459 -977
rect 2259 -1027 2308 -993
rect 2342 -1027 2376 -993
rect 2410 -1027 2459 -993
rect 2259 -1074 2459 -1027
rect 2711 -993 2911 -977
rect 2711 -1027 2760 -993
rect 2794 -1027 2828 -993
rect 2862 -1027 2911 -993
rect 2711 -1074 2911 -1027
rect 2969 -993 3169 -977
rect 2969 -1027 3018 -993
rect 3052 -1027 3086 -993
rect 3120 -1027 3169 -993
rect 2969 -1074 3169 -1027
rect 3227 -993 3427 -977
rect 3227 -1027 3276 -993
rect 3310 -1027 3344 -993
rect 3378 -1027 3427 -993
rect 3227 -1074 3427 -1027
rect 3679 -993 3879 -977
rect 3679 -1027 3728 -993
rect 3762 -1027 3796 -993
rect 3830 -1027 3879 -993
rect 3679 -1074 3879 -1027
rect 3937 -993 4137 -977
rect 3937 -1027 3986 -993
rect 4020 -1027 4054 -993
rect 4088 -1027 4137 -993
rect 3937 -1074 4137 -1027
rect 4195 -993 4395 -977
rect 4195 -1027 4244 -993
rect 4278 -1027 4312 -993
rect 4346 -1027 4395 -993
rect 4195 -1074 4395 -1027
rect 4453 -993 4653 -977
rect 4453 -1027 4502 -993
rect 4536 -1027 4570 -993
rect 4604 -1027 4653 -993
rect 4453 -1074 4653 -1027
rect 4905 -993 5105 -977
rect 4905 -1027 4954 -993
rect 4988 -1027 5022 -993
rect 5056 -1027 5105 -993
rect 4905 -1074 5105 -1027
rect 5391 -993 5591 -977
rect 5391 -1027 5440 -993
rect 5474 -1027 5508 -993
rect 5542 -1027 5591 -993
rect 5391 -1074 5591 -1027
rect 5842 -993 6042 -977
rect 5842 -1027 5891 -993
rect 5925 -1027 5959 -993
rect 5993 -1027 6042 -993
rect 5842 -1074 6042 -1027
rect 6100 -993 6300 -977
rect 6100 -1027 6149 -993
rect 6183 -1027 6217 -993
rect 6251 -1027 6300 -993
rect 6100 -1074 6300 -1027
rect 6358 -993 6558 -977
rect 6358 -1027 6407 -993
rect 6441 -1027 6475 -993
rect 6509 -1027 6558 -993
rect 6358 -1074 6558 -1027
rect 6616 -993 6816 -977
rect 6616 -1027 6665 -993
rect 6699 -1027 6733 -993
rect 6767 -1027 6816 -993
rect 6616 -1074 6816 -1027
rect 7068 -993 7268 -977
rect 7068 -1027 7117 -993
rect 7151 -1027 7185 -993
rect 7219 -1027 7268 -993
rect 7068 -1074 7268 -1027
rect 7326 -993 7526 -977
rect 7326 -1027 7375 -993
rect 7409 -1027 7443 -993
rect 7477 -1027 7526 -993
rect 7326 -1074 7526 -1027
rect 7584 -993 7784 -977
rect 7584 -1027 7633 -993
rect 7667 -1027 7701 -993
rect 7735 -1027 7784 -993
rect 7584 -1074 7784 -1027
rect 8036 -993 8236 -977
rect 8036 -1027 8085 -993
rect 8119 -1027 8153 -993
rect 8187 -1027 8236 -993
rect 8036 -1074 8236 -1027
rect 8294 -993 8494 -977
rect 8294 -1027 8343 -993
rect 8377 -1027 8411 -993
rect 8445 -1027 8494 -993
rect 8294 -1074 8494 -1027
rect 8552 -993 8752 -977
rect 8552 -1027 8601 -993
rect 8635 -1027 8669 -993
rect 8703 -1027 8752 -993
rect 8552 -1074 8752 -1027
rect 8810 -993 9010 -977
rect 8810 -1027 8859 -993
rect 8893 -1027 8927 -993
rect 8961 -1027 9010 -993
rect 8810 -1074 9010 -1027
rect 9262 -993 9462 -977
rect 9262 -1027 9311 -993
rect 9345 -1027 9379 -993
rect 9413 -1027 9462 -993
rect 9262 -1074 9462 -1027
rect 1033 -1300 1233 -1274
rect 1485 -1300 1685 -1274
rect 1743 -1300 1943 -1274
rect 2001 -1300 2201 -1274
rect 2259 -1300 2459 -1274
rect 2711 -1300 2911 -1274
rect 2969 -1300 3169 -1274
rect 3227 -1300 3427 -1274
rect 3679 -1300 3879 -1274
rect 3937 -1300 4137 -1274
rect 4195 -1300 4395 -1274
rect 4453 -1300 4653 -1274
rect 4905 -1300 5105 -1274
rect 5391 -1300 5591 -1274
rect 5842 -1300 6042 -1274
rect 6100 -1300 6300 -1274
rect 6358 -1300 6558 -1274
rect 6616 -1300 6816 -1274
rect 7068 -1300 7268 -1274
rect 7326 -1300 7526 -1274
rect 7584 -1300 7784 -1274
rect 8036 -1300 8236 -1274
rect 8294 -1300 8494 -1274
rect 8552 -1300 8752 -1274
rect 8810 -1300 9010 -1274
rect 9262 -1300 9462 -1274
rect 1033 -2030 1233 -2004
rect 1485 -2030 1685 -2004
rect 1743 -2030 1943 -2004
rect 2001 -2030 2201 -2004
rect 2259 -2030 2459 -2004
rect 2711 -2030 2911 -2004
rect 2969 -2030 3169 -2004
rect 3227 -2030 3427 -2004
rect 3679 -2030 3879 -2004
rect 3937 -2030 4137 -2004
rect 4195 -2030 4395 -2004
rect 4453 -2030 4653 -2004
rect 4905 -2030 5105 -2004
rect 5391 -2030 5591 -2004
rect 5842 -2030 6042 -2004
rect 6100 -2030 6300 -2004
rect 6358 -2030 6558 -2004
rect 6616 -2030 6816 -2004
rect 7068 -2030 7268 -2004
rect 7326 -2030 7526 -2004
rect 7584 -2030 7784 -2004
rect 8036 -2030 8236 -2004
rect 8294 -2030 8494 -2004
rect 8552 -2030 8752 -2004
rect 8810 -2030 9010 -2004
rect 9262 -2030 9462 -2004
rect 1033 -2277 1233 -2230
rect 1033 -2311 1082 -2277
rect 1116 -2311 1150 -2277
rect 1184 -2311 1233 -2277
rect 1033 -2327 1233 -2311
rect 1485 -2277 1685 -2230
rect 1485 -2311 1534 -2277
rect 1568 -2311 1602 -2277
rect 1636 -2311 1685 -2277
rect 1485 -2327 1685 -2311
rect 1743 -2277 1943 -2230
rect 1743 -2311 1792 -2277
rect 1826 -2311 1860 -2277
rect 1894 -2311 1943 -2277
rect 1743 -2327 1943 -2311
rect 2001 -2277 2201 -2230
rect 2001 -2311 2050 -2277
rect 2084 -2311 2118 -2277
rect 2152 -2311 2201 -2277
rect 2001 -2327 2201 -2311
rect 2259 -2277 2459 -2230
rect 2259 -2311 2308 -2277
rect 2342 -2311 2376 -2277
rect 2410 -2311 2459 -2277
rect 2259 -2327 2459 -2311
rect 2711 -2277 2911 -2230
rect 2711 -2311 2760 -2277
rect 2794 -2311 2828 -2277
rect 2862 -2311 2911 -2277
rect 2711 -2327 2911 -2311
rect 2969 -2277 3169 -2230
rect 2969 -2311 3018 -2277
rect 3052 -2311 3086 -2277
rect 3120 -2311 3169 -2277
rect 2969 -2327 3169 -2311
rect 3227 -2277 3427 -2230
rect 3227 -2311 3276 -2277
rect 3310 -2311 3344 -2277
rect 3378 -2311 3427 -2277
rect 3227 -2327 3427 -2311
rect 3679 -2277 3879 -2230
rect 3679 -2311 3728 -2277
rect 3762 -2311 3796 -2277
rect 3830 -2311 3879 -2277
rect 3679 -2327 3879 -2311
rect 3937 -2277 4137 -2230
rect 3937 -2311 3986 -2277
rect 4020 -2311 4054 -2277
rect 4088 -2311 4137 -2277
rect 3937 -2327 4137 -2311
rect 4195 -2277 4395 -2230
rect 4195 -2311 4244 -2277
rect 4278 -2311 4312 -2277
rect 4346 -2311 4395 -2277
rect 4195 -2327 4395 -2311
rect 4453 -2277 4653 -2230
rect 4453 -2311 4502 -2277
rect 4536 -2311 4570 -2277
rect 4604 -2311 4653 -2277
rect 4453 -2327 4653 -2311
rect 4905 -2277 5105 -2230
rect 4905 -2311 4954 -2277
rect 4988 -2311 5022 -2277
rect 5056 -2311 5105 -2277
rect 4905 -2327 5105 -2311
rect 5391 -2277 5591 -2230
rect 5391 -2311 5440 -2277
rect 5474 -2311 5508 -2277
rect 5542 -2311 5591 -2277
rect 5391 -2327 5591 -2311
rect 5842 -2277 6042 -2230
rect 5842 -2311 5891 -2277
rect 5925 -2311 5959 -2277
rect 5993 -2311 6042 -2277
rect 5842 -2327 6042 -2311
rect 6100 -2277 6300 -2230
rect 6100 -2311 6149 -2277
rect 6183 -2311 6217 -2277
rect 6251 -2311 6300 -2277
rect 6100 -2327 6300 -2311
rect 6358 -2277 6558 -2230
rect 6358 -2311 6407 -2277
rect 6441 -2311 6475 -2277
rect 6509 -2311 6558 -2277
rect 6358 -2327 6558 -2311
rect 6616 -2277 6816 -2230
rect 6616 -2311 6665 -2277
rect 6699 -2311 6733 -2277
rect 6767 -2311 6816 -2277
rect 6616 -2327 6816 -2311
rect 7068 -2277 7268 -2230
rect 7068 -2311 7117 -2277
rect 7151 -2311 7185 -2277
rect 7219 -2311 7268 -2277
rect 7068 -2327 7268 -2311
rect 7326 -2277 7526 -2230
rect 7326 -2311 7375 -2277
rect 7409 -2311 7443 -2277
rect 7477 -2311 7526 -2277
rect 7326 -2327 7526 -2311
rect 7584 -2277 7784 -2230
rect 7584 -2311 7633 -2277
rect 7667 -2311 7701 -2277
rect 7735 -2311 7784 -2277
rect 7584 -2327 7784 -2311
rect 8036 -2277 8236 -2230
rect 8036 -2311 8085 -2277
rect 8119 -2311 8153 -2277
rect 8187 -2311 8236 -2277
rect 8036 -2327 8236 -2311
rect 8294 -2277 8494 -2230
rect 8294 -2311 8343 -2277
rect 8377 -2311 8411 -2277
rect 8445 -2311 8494 -2277
rect 8294 -2327 8494 -2311
rect 8552 -2277 8752 -2230
rect 8552 -2311 8601 -2277
rect 8635 -2311 8669 -2277
rect 8703 -2311 8752 -2277
rect 8552 -2327 8752 -2311
rect 8810 -2277 9010 -2230
rect 8810 -2311 8859 -2277
rect 8893 -2311 8927 -2277
rect 8961 -2311 9010 -2277
rect 8810 -2327 9010 -2311
rect 9262 -2277 9462 -2230
rect 9262 -2311 9311 -2277
rect 9345 -2311 9379 -2277
rect 9413 -2311 9462 -2277
rect 9262 -2327 9462 -2311
rect 1033 -2640 1233 -2624
rect 1033 -2674 1082 -2640
rect 1116 -2674 1150 -2640
rect 1184 -2674 1233 -2640
rect 1033 -2721 1233 -2674
rect 1485 -2640 1685 -2624
rect 1485 -2674 1534 -2640
rect 1568 -2674 1602 -2640
rect 1636 -2674 1685 -2640
rect 1485 -2721 1685 -2674
rect 1743 -2640 1943 -2624
rect 1743 -2674 1792 -2640
rect 1826 -2674 1860 -2640
rect 1894 -2674 1943 -2640
rect 1743 -2721 1943 -2674
rect 2001 -2640 2201 -2624
rect 2001 -2674 2050 -2640
rect 2084 -2674 2118 -2640
rect 2152 -2674 2201 -2640
rect 2001 -2721 2201 -2674
rect 2259 -2640 2459 -2624
rect 2259 -2674 2308 -2640
rect 2342 -2674 2376 -2640
rect 2410 -2674 2459 -2640
rect 2259 -2721 2459 -2674
rect 2711 -2640 2911 -2624
rect 2711 -2674 2760 -2640
rect 2794 -2674 2828 -2640
rect 2862 -2674 2911 -2640
rect 2711 -2721 2911 -2674
rect 2969 -2640 3169 -2624
rect 2969 -2674 3018 -2640
rect 3052 -2674 3086 -2640
rect 3120 -2674 3169 -2640
rect 2969 -2721 3169 -2674
rect 3227 -2640 3427 -2624
rect 3227 -2674 3276 -2640
rect 3310 -2674 3344 -2640
rect 3378 -2674 3427 -2640
rect 3227 -2721 3427 -2674
rect 3679 -2640 3879 -2624
rect 3679 -2674 3728 -2640
rect 3762 -2674 3796 -2640
rect 3830 -2674 3879 -2640
rect 3679 -2721 3879 -2674
rect 3937 -2640 4137 -2624
rect 3937 -2674 3986 -2640
rect 4020 -2674 4054 -2640
rect 4088 -2674 4137 -2640
rect 3937 -2721 4137 -2674
rect 4195 -2640 4395 -2624
rect 4195 -2674 4244 -2640
rect 4278 -2674 4312 -2640
rect 4346 -2674 4395 -2640
rect 4195 -2721 4395 -2674
rect 4453 -2640 4653 -2624
rect 4453 -2674 4502 -2640
rect 4536 -2674 4570 -2640
rect 4604 -2674 4653 -2640
rect 4453 -2721 4653 -2674
rect 4905 -2640 5105 -2624
rect 4905 -2674 4954 -2640
rect 4988 -2674 5022 -2640
rect 5056 -2674 5105 -2640
rect 4905 -2721 5105 -2674
rect 5391 -2640 5591 -2624
rect 5391 -2674 5440 -2640
rect 5474 -2674 5508 -2640
rect 5542 -2674 5591 -2640
rect 5391 -2721 5591 -2674
rect 5842 -2640 6042 -2624
rect 5842 -2674 5891 -2640
rect 5925 -2674 5959 -2640
rect 5993 -2674 6042 -2640
rect 5842 -2721 6042 -2674
rect 6100 -2640 6300 -2624
rect 6100 -2674 6149 -2640
rect 6183 -2674 6217 -2640
rect 6251 -2674 6300 -2640
rect 6100 -2721 6300 -2674
rect 6358 -2640 6558 -2624
rect 6358 -2674 6407 -2640
rect 6441 -2674 6475 -2640
rect 6509 -2674 6558 -2640
rect 6358 -2721 6558 -2674
rect 6616 -2640 6816 -2624
rect 6616 -2674 6665 -2640
rect 6699 -2674 6733 -2640
rect 6767 -2674 6816 -2640
rect 6616 -2721 6816 -2674
rect 7068 -2640 7268 -2624
rect 7068 -2674 7117 -2640
rect 7151 -2674 7185 -2640
rect 7219 -2674 7268 -2640
rect 7068 -2721 7268 -2674
rect 7326 -2640 7526 -2624
rect 7326 -2674 7375 -2640
rect 7409 -2674 7443 -2640
rect 7477 -2674 7526 -2640
rect 7326 -2721 7526 -2674
rect 7584 -2640 7784 -2624
rect 7584 -2674 7633 -2640
rect 7667 -2674 7701 -2640
rect 7735 -2674 7784 -2640
rect 7584 -2721 7784 -2674
rect 8036 -2640 8236 -2624
rect 8036 -2674 8085 -2640
rect 8119 -2674 8153 -2640
rect 8187 -2674 8236 -2640
rect 8036 -2721 8236 -2674
rect 8294 -2640 8494 -2624
rect 8294 -2674 8343 -2640
rect 8377 -2674 8411 -2640
rect 8445 -2674 8494 -2640
rect 8294 -2721 8494 -2674
rect 8552 -2640 8752 -2624
rect 8552 -2674 8601 -2640
rect 8635 -2674 8669 -2640
rect 8703 -2674 8752 -2640
rect 8552 -2721 8752 -2674
rect 8810 -2640 9010 -2624
rect 8810 -2674 8859 -2640
rect 8893 -2674 8927 -2640
rect 8961 -2674 9010 -2640
rect 8810 -2721 9010 -2674
rect 9262 -2640 9462 -2624
rect 9262 -2674 9311 -2640
rect 9345 -2674 9379 -2640
rect 9413 -2674 9462 -2640
rect 9262 -2721 9462 -2674
rect 1033 -2947 1233 -2921
rect 1485 -2947 1685 -2921
rect 1743 -2947 1943 -2921
rect 2001 -2947 2201 -2921
rect 2259 -2947 2459 -2921
rect 2711 -2947 2911 -2921
rect 2969 -2947 3169 -2921
rect 3227 -2947 3427 -2921
rect 3679 -2947 3879 -2921
rect 3937 -2947 4137 -2921
rect 4195 -2947 4395 -2921
rect 4453 -2947 4653 -2921
rect 4905 -2947 5105 -2921
rect 5391 -2947 5591 -2921
rect 5842 -2947 6042 -2921
rect 6100 -2947 6300 -2921
rect 6358 -2947 6558 -2921
rect 6616 -2947 6816 -2921
rect 7068 -2947 7268 -2921
rect 7326 -2947 7526 -2921
rect 7584 -2947 7784 -2921
rect 8036 -2947 8236 -2921
rect 8294 -2947 8494 -2921
rect 8552 -2947 8752 -2921
rect 8810 -2947 9010 -2921
rect 9262 -2947 9462 -2921
rect 1033 -3711 1233 -3685
rect 1485 -3711 1685 -3685
rect 1743 -3711 1943 -3685
rect 2001 -3711 2201 -3685
rect 2259 -3711 2459 -3685
rect 2711 -3711 2911 -3685
rect 2969 -3711 3169 -3685
rect 3227 -3711 3427 -3685
rect 3679 -3711 3879 -3685
rect 3937 -3711 4137 -3685
rect 4195 -3711 4395 -3685
rect 4453 -3711 4653 -3685
rect 4905 -3711 5105 -3685
rect 5391 -3711 5591 -3685
rect 5842 -3711 6042 -3685
rect 6100 -3711 6300 -3685
rect 6358 -3711 6558 -3685
rect 6616 -3711 6816 -3685
rect 7068 -3711 7268 -3685
rect 7326 -3711 7526 -3685
rect 7584 -3711 7784 -3685
rect 8036 -3711 8236 -3685
rect 8294 -3711 8494 -3685
rect 8552 -3711 8752 -3685
rect 8810 -3711 9010 -3685
rect 9262 -3711 9462 -3685
rect 1033 -3958 1233 -3911
rect 1033 -3992 1082 -3958
rect 1116 -3992 1150 -3958
rect 1184 -3992 1233 -3958
rect 1033 -4008 1233 -3992
rect 1485 -3958 1685 -3911
rect 1485 -3992 1534 -3958
rect 1568 -3992 1602 -3958
rect 1636 -3992 1685 -3958
rect 1485 -4008 1685 -3992
rect 1743 -3958 1943 -3911
rect 1743 -3992 1792 -3958
rect 1826 -3992 1860 -3958
rect 1894 -3992 1943 -3958
rect 1743 -4008 1943 -3992
rect 2001 -3958 2201 -3911
rect 2001 -3992 2050 -3958
rect 2084 -3992 2118 -3958
rect 2152 -3992 2201 -3958
rect 2001 -4008 2201 -3992
rect 2259 -3958 2459 -3911
rect 2259 -3992 2308 -3958
rect 2342 -3992 2376 -3958
rect 2410 -3992 2459 -3958
rect 2259 -4008 2459 -3992
rect 2711 -3958 2911 -3911
rect 2711 -3992 2760 -3958
rect 2794 -3992 2828 -3958
rect 2862 -3992 2911 -3958
rect 2711 -4008 2911 -3992
rect 2969 -3958 3169 -3911
rect 2969 -3992 3018 -3958
rect 3052 -3992 3086 -3958
rect 3120 -3992 3169 -3958
rect 2969 -4008 3169 -3992
rect 3227 -3958 3427 -3911
rect 3227 -3992 3276 -3958
rect 3310 -3992 3344 -3958
rect 3378 -3992 3427 -3958
rect 3227 -4008 3427 -3992
rect 3679 -3958 3879 -3911
rect 3679 -3992 3728 -3958
rect 3762 -3992 3796 -3958
rect 3830 -3992 3879 -3958
rect 3679 -4008 3879 -3992
rect 3937 -3958 4137 -3911
rect 3937 -3992 3986 -3958
rect 4020 -3992 4054 -3958
rect 4088 -3992 4137 -3958
rect 3937 -4008 4137 -3992
rect 4195 -3958 4395 -3911
rect 4195 -3992 4244 -3958
rect 4278 -3992 4312 -3958
rect 4346 -3992 4395 -3958
rect 4195 -4008 4395 -3992
rect 4453 -3958 4653 -3911
rect 4453 -3992 4502 -3958
rect 4536 -3992 4570 -3958
rect 4604 -3992 4653 -3958
rect 4453 -4008 4653 -3992
rect 4905 -3958 5105 -3911
rect 4905 -3992 4954 -3958
rect 4988 -3992 5022 -3958
rect 5056 -3992 5105 -3958
rect 4905 -4008 5105 -3992
rect 5391 -3958 5591 -3911
rect 5391 -3992 5440 -3958
rect 5474 -3992 5508 -3958
rect 5542 -3992 5591 -3958
rect 5391 -4008 5591 -3992
rect 5842 -3958 6042 -3911
rect 5842 -3992 5891 -3958
rect 5925 -3992 5959 -3958
rect 5993 -3992 6042 -3958
rect 5842 -4008 6042 -3992
rect 6100 -3958 6300 -3911
rect 6100 -3992 6149 -3958
rect 6183 -3992 6217 -3958
rect 6251 -3992 6300 -3958
rect 6100 -4008 6300 -3992
rect 6358 -3958 6558 -3911
rect 6358 -3992 6407 -3958
rect 6441 -3992 6475 -3958
rect 6509 -3992 6558 -3958
rect 6358 -4008 6558 -3992
rect 6616 -3958 6816 -3911
rect 6616 -3992 6665 -3958
rect 6699 -3992 6733 -3958
rect 6767 -3992 6816 -3958
rect 6616 -4008 6816 -3992
rect 7068 -3958 7268 -3911
rect 7068 -3992 7117 -3958
rect 7151 -3992 7185 -3958
rect 7219 -3992 7268 -3958
rect 7068 -4008 7268 -3992
rect 7326 -3958 7526 -3911
rect 7326 -3992 7375 -3958
rect 7409 -3992 7443 -3958
rect 7477 -3992 7526 -3958
rect 7326 -4008 7526 -3992
rect 7584 -3958 7784 -3911
rect 7584 -3992 7633 -3958
rect 7667 -3992 7701 -3958
rect 7735 -3992 7784 -3958
rect 7584 -4008 7784 -3992
rect 8036 -3958 8236 -3911
rect 8036 -3992 8085 -3958
rect 8119 -3992 8153 -3958
rect 8187 -3992 8236 -3958
rect 8036 -4008 8236 -3992
rect 8294 -3958 8494 -3911
rect 8294 -3992 8343 -3958
rect 8377 -3992 8411 -3958
rect 8445 -3992 8494 -3958
rect 8294 -4008 8494 -3992
rect 8552 -3958 8752 -3911
rect 8552 -3992 8601 -3958
rect 8635 -3992 8669 -3958
rect 8703 -3992 8752 -3958
rect 8552 -4008 8752 -3992
rect 8810 -3958 9010 -3911
rect 8810 -3992 8859 -3958
rect 8893 -3992 8927 -3958
rect 8961 -3992 9010 -3958
rect 8810 -4008 9010 -3992
rect 9262 -3958 9462 -3911
rect 9262 -3992 9311 -3958
rect 9345 -3992 9379 -3958
rect 9413 -3992 9462 -3958
rect 9262 -4008 9462 -3992
rect 1033 -4186 1233 -4170
rect 1033 -4220 1082 -4186
rect 1116 -4220 1150 -4186
rect 1184 -4220 1233 -4186
rect 1033 -4267 1233 -4220
rect 1485 -4186 1685 -4170
rect 1485 -4220 1534 -4186
rect 1568 -4220 1602 -4186
rect 1636 -4220 1685 -4186
rect 1485 -4267 1685 -4220
rect 1743 -4186 1943 -4170
rect 1743 -4220 1792 -4186
rect 1826 -4220 1860 -4186
rect 1894 -4220 1943 -4186
rect 1743 -4267 1943 -4220
rect 2001 -4186 2201 -4170
rect 2001 -4220 2050 -4186
rect 2084 -4220 2118 -4186
rect 2152 -4220 2201 -4186
rect 2001 -4267 2201 -4220
rect 2259 -4186 2459 -4170
rect 2259 -4220 2308 -4186
rect 2342 -4220 2376 -4186
rect 2410 -4220 2459 -4186
rect 2259 -4267 2459 -4220
rect 2711 -4186 2911 -4170
rect 2711 -4220 2760 -4186
rect 2794 -4220 2828 -4186
rect 2862 -4220 2911 -4186
rect 2711 -4267 2911 -4220
rect 2969 -4186 3169 -4170
rect 2969 -4220 3018 -4186
rect 3052 -4220 3086 -4186
rect 3120 -4220 3169 -4186
rect 2969 -4267 3169 -4220
rect 3227 -4186 3427 -4170
rect 3227 -4220 3276 -4186
rect 3310 -4220 3344 -4186
rect 3378 -4220 3427 -4186
rect 3227 -4267 3427 -4220
rect 3679 -4186 3879 -4170
rect 3679 -4220 3728 -4186
rect 3762 -4220 3796 -4186
rect 3830 -4220 3879 -4186
rect 3679 -4267 3879 -4220
rect 3937 -4186 4137 -4170
rect 3937 -4220 3986 -4186
rect 4020 -4220 4054 -4186
rect 4088 -4220 4137 -4186
rect 3937 -4267 4137 -4220
rect 4195 -4186 4395 -4170
rect 4195 -4220 4244 -4186
rect 4278 -4220 4312 -4186
rect 4346 -4220 4395 -4186
rect 4195 -4267 4395 -4220
rect 4453 -4186 4653 -4170
rect 4453 -4220 4502 -4186
rect 4536 -4220 4570 -4186
rect 4604 -4220 4653 -4186
rect 4453 -4267 4653 -4220
rect 4905 -4186 5105 -4170
rect 4905 -4220 4954 -4186
rect 4988 -4220 5022 -4186
rect 5056 -4220 5105 -4186
rect 4905 -4267 5105 -4220
rect 5391 -4186 5591 -4170
rect 5391 -4220 5440 -4186
rect 5474 -4220 5508 -4186
rect 5542 -4220 5591 -4186
rect 5391 -4267 5591 -4220
rect 5842 -4186 6042 -4170
rect 5842 -4220 5891 -4186
rect 5925 -4220 5959 -4186
rect 5993 -4220 6042 -4186
rect 5842 -4267 6042 -4220
rect 6100 -4186 6300 -4170
rect 6100 -4220 6149 -4186
rect 6183 -4220 6217 -4186
rect 6251 -4220 6300 -4186
rect 6100 -4267 6300 -4220
rect 6358 -4186 6558 -4170
rect 6358 -4220 6407 -4186
rect 6441 -4220 6475 -4186
rect 6509 -4220 6558 -4186
rect 6358 -4267 6558 -4220
rect 6616 -4186 6816 -4170
rect 6616 -4220 6665 -4186
rect 6699 -4220 6733 -4186
rect 6767 -4220 6816 -4186
rect 6616 -4267 6816 -4220
rect 7068 -4186 7268 -4170
rect 7068 -4220 7117 -4186
rect 7151 -4220 7185 -4186
rect 7219 -4220 7268 -4186
rect 7068 -4267 7268 -4220
rect 7326 -4186 7526 -4170
rect 7326 -4220 7375 -4186
rect 7409 -4220 7443 -4186
rect 7477 -4220 7526 -4186
rect 7326 -4267 7526 -4220
rect 7584 -4186 7784 -4170
rect 7584 -4220 7633 -4186
rect 7667 -4220 7701 -4186
rect 7735 -4220 7784 -4186
rect 7584 -4267 7784 -4220
rect 8036 -4186 8236 -4170
rect 8036 -4220 8085 -4186
rect 8119 -4220 8153 -4186
rect 8187 -4220 8236 -4186
rect 8036 -4267 8236 -4220
rect 8294 -4186 8494 -4170
rect 8294 -4220 8343 -4186
rect 8377 -4220 8411 -4186
rect 8445 -4220 8494 -4186
rect 8294 -4267 8494 -4220
rect 8552 -4186 8752 -4170
rect 8552 -4220 8601 -4186
rect 8635 -4220 8669 -4186
rect 8703 -4220 8752 -4186
rect 8552 -4267 8752 -4220
rect 8810 -4186 9010 -4170
rect 8810 -4220 8859 -4186
rect 8893 -4220 8927 -4186
rect 8961 -4220 9010 -4186
rect 8810 -4267 9010 -4220
rect 9262 -4186 9462 -4170
rect 9262 -4220 9311 -4186
rect 9345 -4220 9379 -4186
rect 9413 -4220 9462 -4186
rect 9262 -4267 9462 -4220
rect 1033 -4493 1233 -4467
rect 1485 -4493 1685 -4467
rect 1743 -4493 1943 -4467
rect 2001 -4493 2201 -4467
rect 2259 -4493 2459 -4467
rect 2711 -4493 2911 -4467
rect 2969 -4493 3169 -4467
rect 3227 -4493 3427 -4467
rect 3679 -4493 3879 -4467
rect 3937 -4493 4137 -4467
rect 4195 -4493 4395 -4467
rect 4453 -4493 4653 -4467
rect 4905 -4493 5105 -4467
rect 5391 -4493 5591 -4467
rect 5842 -4493 6042 -4467
rect 6100 -4493 6300 -4467
rect 6358 -4493 6558 -4467
rect 6616 -4493 6816 -4467
rect 7068 -4493 7268 -4467
rect 7326 -4493 7526 -4467
rect 7584 -4493 7784 -4467
rect 8036 -4493 8236 -4467
rect 8294 -4493 8494 -4467
rect 8552 -4493 8752 -4467
rect 8810 -4493 9010 -4467
rect 9262 -4493 9462 -4467
rect 1033 -5257 1233 -5231
rect 1485 -5257 1685 -5231
rect 1743 -5257 1943 -5231
rect 2001 -5257 2201 -5231
rect 2259 -5257 2459 -5231
rect 2711 -5257 2911 -5231
rect 2969 -5257 3169 -5231
rect 3227 -5257 3427 -5231
rect 3679 -5257 3879 -5231
rect 3937 -5257 4137 -5231
rect 4195 -5257 4395 -5231
rect 4453 -5257 4653 -5231
rect 4905 -5257 5105 -5231
rect 5391 -5257 5591 -5231
rect 5842 -5257 6042 -5231
rect 6100 -5257 6300 -5231
rect 6358 -5257 6558 -5231
rect 6616 -5257 6816 -5231
rect 7068 -5257 7268 -5231
rect 7326 -5257 7526 -5231
rect 7584 -5257 7784 -5231
rect 8036 -5257 8236 -5231
rect 8294 -5257 8494 -5231
rect 8552 -5257 8752 -5231
rect 8810 -5257 9010 -5231
rect 9262 -5257 9462 -5231
rect 1033 -5504 1233 -5457
rect 1033 -5538 1082 -5504
rect 1116 -5538 1150 -5504
rect 1184 -5538 1233 -5504
rect 1033 -5554 1233 -5538
rect 1485 -5504 1685 -5457
rect 1485 -5538 1534 -5504
rect 1568 -5538 1602 -5504
rect 1636 -5538 1685 -5504
rect 1485 -5554 1685 -5538
rect 1743 -5504 1943 -5457
rect 1743 -5538 1792 -5504
rect 1826 -5538 1860 -5504
rect 1894 -5538 1943 -5504
rect 1743 -5554 1943 -5538
rect 2001 -5504 2201 -5457
rect 2001 -5538 2050 -5504
rect 2084 -5538 2118 -5504
rect 2152 -5538 2201 -5504
rect 2001 -5554 2201 -5538
rect 2259 -5504 2459 -5457
rect 2259 -5538 2308 -5504
rect 2342 -5538 2376 -5504
rect 2410 -5538 2459 -5504
rect 2259 -5554 2459 -5538
rect 2711 -5504 2911 -5457
rect 2711 -5538 2760 -5504
rect 2794 -5538 2828 -5504
rect 2862 -5538 2911 -5504
rect 2711 -5554 2911 -5538
rect 2969 -5504 3169 -5457
rect 2969 -5538 3018 -5504
rect 3052 -5538 3086 -5504
rect 3120 -5538 3169 -5504
rect 2969 -5554 3169 -5538
rect 3227 -5504 3427 -5457
rect 3227 -5538 3276 -5504
rect 3310 -5538 3344 -5504
rect 3378 -5538 3427 -5504
rect 3227 -5554 3427 -5538
rect 3679 -5504 3879 -5457
rect 3679 -5538 3728 -5504
rect 3762 -5538 3796 -5504
rect 3830 -5538 3879 -5504
rect 3679 -5554 3879 -5538
rect 3937 -5504 4137 -5457
rect 3937 -5538 3986 -5504
rect 4020 -5538 4054 -5504
rect 4088 -5538 4137 -5504
rect 3937 -5554 4137 -5538
rect 4195 -5504 4395 -5457
rect 4195 -5538 4244 -5504
rect 4278 -5538 4312 -5504
rect 4346 -5538 4395 -5504
rect 4195 -5554 4395 -5538
rect 4453 -5504 4653 -5457
rect 4453 -5538 4502 -5504
rect 4536 -5538 4570 -5504
rect 4604 -5538 4653 -5504
rect 4453 -5554 4653 -5538
rect 4905 -5504 5105 -5457
rect 4905 -5538 4954 -5504
rect 4988 -5538 5022 -5504
rect 5056 -5538 5105 -5504
rect 4905 -5554 5105 -5538
rect 5391 -5504 5591 -5457
rect 5391 -5538 5440 -5504
rect 5474 -5538 5508 -5504
rect 5542 -5538 5591 -5504
rect 5391 -5554 5591 -5538
rect 5842 -5504 6042 -5457
rect 5842 -5538 5891 -5504
rect 5925 -5538 5959 -5504
rect 5993 -5538 6042 -5504
rect 5842 -5554 6042 -5538
rect 6100 -5504 6300 -5457
rect 6100 -5538 6149 -5504
rect 6183 -5538 6217 -5504
rect 6251 -5538 6300 -5504
rect 6100 -5554 6300 -5538
rect 6358 -5504 6558 -5457
rect 6358 -5538 6407 -5504
rect 6441 -5538 6475 -5504
rect 6509 -5538 6558 -5504
rect 6358 -5554 6558 -5538
rect 6616 -5504 6816 -5457
rect 6616 -5538 6665 -5504
rect 6699 -5538 6733 -5504
rect 6767 -5538 6816 -5504
rect 6616 -5554 6816 -5538
rect 7068 -5504 7268 -5457
rect 7068 -5538 7117 -5504
rect 7151 -5538 7185 -5504
rect 7219 -5538 7268 -5504
rect 7068 -5554 7268 -5538
rect 7326 -5504 7526 -5457
rect 7326 -5538 7375 -5504
rect 7409 -5538 7443 -5504
rect 7477 -5538 7526 -5504
rect 7326 -5554 7526 -5538
rect 7584 -5504 7784 -5457
rect 7584 -5538 7633 -5504
rect 7667 -5538 7701 -5504
rect 7735 -5538 7784 -5504
rect 7584 -5554 7784 -5538
rect 8036 -5504 8236 -5457
rect 8036 -5538 8085 -5504
rect 8119 -5538 8153 -5504
rect 8187 -5538 8236 -5504
rect 8036 -5554 8236 -5538
rect 8294 -5504 8494 -5457
rect 8294 -5538 8343 -5504
rect 8377 -5538 8411 -5504
rect 8445 -5538 8494 -5504
rect 8294 -5554 8494 -5538
rect 8552 -5504 8752 -5457
rect 8552 -5538 8601 -5504
rect 8635 -5538 8669 -5504
rect 8703 -5538 8752 -5504
rect 8552 -5554 8752 -5538
rect 8810 -5504 9010 -5457
rect 8810 -5538 8859 -5504
rect 8893 -5538 8927 -5504
rect 8961 -5538 9010 -5504
rect 8810 -5554 9010 -5538
rect 9262 -5504 9462 -5457
rect 9262 -5538 9311 -5504
rect 9345 -5538 9379 -5504
rect 9413 -5538 9462 -5504
rect 9262 -5554 9462 -5538
rect 1033 -5866 1233 -5850
rect 1033 -5900 1082 -5866
rect 1116 -5900 1150 -5866
rect 1184 -5900 1233 -5866
rect 1033 -5947 1233 -5900
rect 1485 -5866 1685 -5850
rect 1485 -5900 1534 -5866
rect 1568 -5900 1602 -5866
rect 1636 -5900 1685 -5866
rect 1485 -5947 1685 -5900
rect 1743 -5866 1943 -5850
rect 1743 -5900 1792 -5866
rect 1826 -5900 1860 -5866
rect 1894 -5900 1943 -5866
rect 1743 -5947 1943 -5900
rect 2001 -5866 2201 -5850
rect 2001 -5900 2050 -5866
rect 2084 -5900 2118 -5866
rect 2152 -5900 2201 -5866
rect 2001 -5947 2201 -5900
rect 2259 -5866 2459 -5850
rect 2259 -5900 2308 -5866
rect 2342 -5900 2376 -5866
rect 2410 -5900 2459 -5866
rect 2259 -5947 2459 -5900
rect 2711 -5866 2911 -5850
rect 2711 -5900 2760 -5866
rect 2794 -5900 2828 -5866
rect 2862 -5900 2911 -5866
rect 2711 -5947 2911 -5900
rect 2969 -5866 3169 -5850
rect 2969 -5900 3018 -5866
rect 3052 -5900 3086 -5866
rect 3120 -5900 3169 -5866
rect 2969 -5947 3169 -5900
rect 3227 -5866 3427 -5850
rect 3227 -5900 3276 -5866
rect 3310 -5900 3344 -5866
rect 3378 -5900 3427 -5866
rect 3227 -5947 3427 -5900
rect 3679 -5866 3879 -5850
rect 3679 -5900 3728 -5866
rect 3762 -5900 3796 -5866
rect 3830 -5900 3879 -5866
rect 3679 -5947 3879 -5900
rect 3937 -5866 4137 -5850
rect 3937 -5900 3986 -5866
rect 4020 -5900 4054 -5866
rect 4088 -5900 4137 -5866
rect 3937 -5947 4137 -5900
rect 4195 -5866 4395 -5850
rect 4195 -5900 4244 -5866
rect 4278 -5900 4312 -5866
rect 4346 -5900 4395 -5866
rect 4195 -5947 4395 -5900
rect 4453 -5866 4653 -5850
rect 4453 -5900 4502 -5866
rect 4536 -5900 4570 -5866
rect 4604 -5900 4653 -5866
rect 4453 -5947 4653 -5900
rect 4905 -5866 5105 -5850
rect 4905 -5900 4954 -5866
rect 4988 -5900 5022 -5866
rect 5056 -5900 5105 -5866
rect 4905 -5947 5105 -5900
rect 5391 -5866 5591 -5850
rect 5391 -5900 5440 -5866
rect 5474 -5900 5508 -5866
rect 5542 -5900 5591 -5866
rect 5391 -5947 5591 -5900
rect 5842 -5866 6042 -5850
rect 5842 -5900 5891 -5866
rect 5925 -5900 5959 -5866
rect 5993 -5900 6042 -5866
rect 5842 -5947 6042 -5900
rect 6100 -5866 6300 -5850
rect 6100 -5900 6149 -5866
rect 6183 -5900 6217 -5866
rect 6251 -5900 6300 -5866
rect 6100 -5947 6300 -5900
rect 6358 -5866 6558 -5850
rect 6358 -5900 6407 -5866
rect 6441 -5900 6475 -5866
rect 6509 -5900 6558 -5866
rect 6358 -5947 6558 -5900
rect 6616 -5866 6816 -5850
rect 6616 -5900 6665 -5866
rect 6699 -5900 6733 -5866
rect 6767 -5900 6816 -5866
rect 6616 -5947 6816 -5900
rect 7068 -5866 7268 -5850
rect 7068 -5900 7117 -5866
rect 7151 -5900 7185 -5866
rect 7219 -5900 7268 -5866
rect 7068 -5947 7268 -5900
rect 7326 -5866 7526 -5850
rect 7326 -5900 7375 -5866
rect 7409 -5900 7443 -5866
rect 7477 -5900 7526 -5866
rect 7326 -5947 7526 -5900
rect 7584 -5866 7784 -5850
rect 7584 -5900 7633 -5866
rect 7667 -5900 7701 -5866
rect 7735 -5900 7784 -5866
rect 7584 -5947 7784 -5900
rect 8036 -5866 8236 -5850
rect 8036 -5900 8085 -5866
rect 8119 -5900 8153 -5866
rect 8187 -5900 8236 -5866
rect 8036 -5947 8236 -5900
rect 8294 -5866 8494 -5850
rect 8294 -5900 8343 -5866
rect 8377 -5900 8411 -5866
rect 8445 -5900 8494 -5866
rect 8294 -5947 8494 -5900
rect 8552 -5866 8752 -5850
rect 8552 -5900 8601 -5866
rect 8635 -5900 8669 -5866
rect 8703 -5900 8752 -5866
rect 8552 -5947 8752 -5900
rect 8810 -5866 9010 -5850
rect 8810 -5900 8859 -5866
rect 8893 -5900 8927 -5866
rect 8961 -5900 9010 -5866
rect 8810 -5947 9010 -5900
rect 9262 -5866 9462 -5850
rect 9262 -5900 9311 -5866
rect 9345 -5900 9379 -5866
rect 9413 -5900 9462 -5866
rect 9262 -5947 9462 -5900
rect 1033 -6173 1233 -6147
rect 1485 -6173 1685 -6147
rect 1743 -6173 1943 -6147
rect 2001 -6173 2201 -6147
rect 2259 -6173 2459 -6147
rect 2711 -6173 2911 -6147
rect 2969 -6173 3169 -6147
rect 3227 -6173 3427 -6147
rect 3679 -6173 3879 -6147
rect 3937 -6173 4137 -6147
rect 4195 -6173 4395 -6147
rect 4453 -6173 4653 -6147
rect 4905 -6173 5105 -6147
rect 5391 -6173 5591 -6147
rect 5842 -6173 6042 -6147
rect 6100 -6173 6300 -6147
rect 6358 -6173 6558 -6147
rect 6616 -6173 6816 -6147
rect 7068 -6173 7268 -6147
rect 7326 -6173 7526 -6147
rect 7584 -6173 7784 -6147
rect 8036 -6173 8236 -6147
rect 8294 -6173 8494 -6147
rect 8552 -6173 8752 -6147
rect 8810 -6173 9010 -6147
rect 9262 -6173 9462 -6147
rect 1033 -6904 1233 -6878
rect 1485 -6904 1685 -6878
rect 1743 -6904 1943 -6878
rect 2001 -6904 2201 -6878
rect 2259 -6904 2459 -6878
rect 2711 -6904 2911 -6878
rect 2969 -6904 3169 -6878
rect 3227 -6904 3427 -6878
rect 3679 -6904 3879 -6878
rect 3937 -6904 4137 -6878
rect 4195 -6904 4395 -6878
rect 4453 -6904 4653 -6878
rect 4905 -6904 5105 -6878
rect 5391 -6904 5591 -6878
rect 5842 -6904 6042 -6878
rect 6100 -6904 6300 -6878
rect 6358 -6904 6558 -6878
rect 6616 -6904 6816 -6878
rect 7068 -6904 7268 -6878
rect 7326 -6904 7526 -6878
rect 7584 -6904 7784 -6878
rect 8036 -6904 8236 -6878
rect 8294 -6904 8494 -6878
rect 8552 -6904 8752 -6878
rect 8810 -6904 9010 -6878
rect 9262 -6904 9462 -6878
rect 1033 -7151 1233 -7104
rect 1033 -7185 1082 -7151
rect 1116 -7185 1150 -7151
rect 1184 -7185 1233 -7151
rect 1033 -7201 1233 -7185
rect 1485 -7151 1685 -7104
rect 1485 -7185 1534 -7151
rect 1568 -7185 1602 -7151
rect 1636 -7185 1685 -7151
rect 1485 -7201 1685 -7185
rect 1743 -7151 1943 -7104
rect 1743 -7185 1792 -7151
rect 1826 -7185 1860 -7151
rect 1894 -7185 1943 -7151
rect 1743 -7201 1943 -7185
rect 2001 -7151 2201 -7104
rect 2001 -7185 2050 -7151
rect 2084 -7185 2118 -7151
rect 2152 -7185 2201 -7151
rect 2001 -7201 2201 -7185
rect 2259 -7151 2459 -7104
rect 2259 -7185 2308 -7151
rect 2342 -7185 2376 -7151
rect 2410 -7185 2459 -7151
rect 2259 -7201 2459 -7185
rect 2711 -7151 2911 -7104
rect 2711 -7185 2760 -7151
rect 2794 -7185 2828 -7151
rect 2862 -7185 2911 -7151
rect 2711 -7201 2911 -7185
rect 2969 -7151 3169 -7104
rect 2969 -7185 3018 -7151
rect 3052 -7185 3086 -7151
rect 3120 -7185 3169 -7151
rect 2969 -7201 3169 -7185
rect 3227 -7151 3427 -7104
rect 3227 -7185 3276 -7151
rect 3310 -7185 3344 -7151
rect 3378 -7185 3427 -7151
rect 3227 -7201 3427 -7185
rect 3679 -7151 3879 -7104
rect 3679 -7185 3728 -7151
rect 3762 -7185 3796 -7151
rect 3830 -7185 3879 -7151
rect 3679 -7201 3879 -7185
rect 3937 -7151 4137 -7104
rect 3937 -7185 3986 -7151
rect 4020 -7185 4054 -7151
rect 4088 -7185 4137 -7151
rect 3937 -7201 4137 -7185
rect 4195 -7151 4395 -7104
rect 4195 -7185 4244 -7151
rect 4278 -7185 4312 -7151
rect 4346 -7185 4395 -7151
rect 4195 -7201 4395 -7185
rect 4453 -7151 4653 -7104
rect 4453 -7185 4502 -7151
rect 4536 -7185 4570 -7151
rect 4604 -7185 4653 -7151
rect 4453 -7201 4653 -7185
rect 4905 -7151 5105 -7104
rect 4905 -7185 4954 -7151
rect 4988 -7185 5022 -7151
rect 5056 -7185 5105 -7151
rect 4905 -7201 5105 -7185
rect 5391 -7151 5591 -7104
rect 5391 -7185 5440 -7151
rect 5474 -7185 5508 -7151
rect 5542 -7185 5591 -7151
rect 5391 -7201 5591 -7185
rect 5842 -7151 6042 -7104
rect 5842 -7185 5891 -7151
rect 5925 -7185 5959 -7151
rect 5993 -7185 6042 -7151
rect 5842 -7201 6042 -7185
rect 6100 -7151 6300 -7104
rect 6100 -7185 6149 -7151
rect 6183 -7185 6217 -7151
rect 6251 -7185 6300 -7151
rect 6100 -7201 6300 -7185
rect 6358 -7151 6558 -7104
rect 6358 -7185 6407 -7151
rect 6441 -7185 6475 -7151
rect 6509 -7185 6558 -7151
rect 6358 -7201 6558 -7185
rect 6616 -7151 6816 -7104
rect 6616 -7185 6665 -7151
rect 6699 -7185 6733 -7151
rect 6767 -7185 6816 -7151
rect 6616 -7201 6816 -7185
rect 7068 -7151 7268 -7104
rect 7068 -7185 7117 -7151
rect 7151 -7185 7185 -7151
rect 7219 -7185 7268 -7151
rect 7068 -7201 7268 -7185
rect 7326 -7151 7526 -7104
rect 7326 -7185 7375 -7151
rect 7409 -7185 7443 -7151
rect 7477 -7185 7526 -7151
rect 7326 -7201 7526 -7185
rect 7584 -7151 7784 -7104
rect 7584 -7185 7633 -7151
rect 7667 -7185 7701 -7151
rect 7735 -7185 7784 -7151
rect 7584 -7201 7784 -7185
rect 8036 -7151 8236 -7104
rect 8036 -7185 8085 -7151
rect 8119 -7185 8153 -7151
rect 8187 -7185 8236 -7151
rect 8036 -7201 8236 -7185
rect 8294 -7151 8494 -7104
rect 8294 -7185 8343 -7151
rect 8377 -7185 8411 -7151
rect 8445 -7185 8494 -7151
rect 8294 -7201 8494 -7185
rect 8552 -7151 8752 -7104
rect 8552 -7185 8601 -7151
rect 8635 -7185 8669 -7151
rect 8703 -7185 8752 -7151
rect 8552 -7201 8752 -7185
rect 8810 -7151 9010 -7104
rect 8810 -7185 8859 -7151
rect 8893 -7185 8927 -7151
rect 8961 -7185 9010 -7151
rect 8810 -7201 9010 -7185
rect 9262 -7151 9462 -7104
rect 9262 -7185 9311 -7151
rect 9345 -7185 9379 -7151
rect 9413 -7185 9462 -7151
rect 9262 -7201 9462 -7185
rect 1033 -7513 1233 -7497
rect 1033 -7547 1082 -7513
rect 1116 -7547 1150 -7513
rect 1184 -7547 1233 -7513
rect 1033 -7594 1233 -7547
rect 1485 -7513 1685 -7497
rect 1485 -7547 1534 -7513
rect 1568 -7547 1602 -7513
rect 1636 -7547 1685 -7513
rect 1485 -7594 1685 -7547
rect 1743 -7513 1943 -7497
rect 1743 -7547 1792 -7513
rect 1826 -7547 1860 -7513
rect 1894 -7547 1943 -7513
rect 1743 -7594 1943 -7547
rect 2001 -7513 2201 -7497
rect 2001 -7547 2050 -7513
rect 2084 -7547 2118 -7513
rect 2152 -7547 2201 -7513
rect 2001 -7594 2201 -7547
rect 2259 -7513 2459 -7497
rect 2259 -7547 2308 -7513
rect 2342 -7547 2376 -7513
rect 2410 -7547 2459 -7513
rect 2259 -7594 2459 -7547
rect 2711 -7513 2911 -7497
rect 2711 -7547 2760 -7513
rect 2794 -7547 2828 -7513
rect 2862 -7547 2911 -7513
rect 2711 -7594 2911 -7547
rect 2969 -7513 3169 -7497
rect 2969 -7547 3018 -7513
rect 3052 -7547 3086 -7513
rect 3120 -7547 3169 -7513
rect 2969 -7594 3169 -7547
rect 3227 -7513 3427 -7497
rect 3227 -7547 3276 -7513
rect 3310 -7547 3344 -7513
rect 3378 -7547 3427 -7513
rect 3227 -7594 3427 -7547
rect 3679 -7513 3879 -7497
rect 3679 -7547 3728 -7513
rect 3762 -7547 3796 -7513
rect 3830 -7547 3879 -7513
rect 3679 -7594 3879 -7547
rect 3937 -7513 4137 -7497
rect 3937 -7547 3986 -7513
rect 4020 -7547 4054 -7513
rect 4088 -7547 4137 -7513
rect 3937 -7594 4137 -7547
rect 4195 -7513 4395 -7497
rect 4195 -7547 4244 -7513
rect 4278 -7547 4312 -7513
rect 4346 -7547 4395 -7513
rect 4195 -7594 4395 -7547
rect 4453 -7513 4653 -7497
rect 4453 -7547 4502 -7513
rect 4536 -7547 4570 -7513
rect 4604 -7547 4653 -7513
rect 4453 -7594 4653 -7547
rect 4905 -7513 5105 -7497
rect 4905 -7547 4954 -7513
rect 4988 -7547 5022 -7513
rect 5056 -7547 5105 -7513
rect 4905 -7594 5105 -7547
rect 5391 -7513 5591 -7497
rect 5391 -7547 5440 -7513
rect 5474 -7547 5508 -7513
rect 5542 -7547 5591 -7513
rect 5391 -7594 5591 -7547
rect 5842 -7513 6042 -7497
rect 5842 -7547 5891 -7513
rect 5925 -7547 5959 -7513
rect 5993 -7547 6042 -7513
rect 5842 -7594 6042 -7547
rect 6100 -7513 6300 -7497
rect 6100 -7547 6149 -7513
rect 6183 -7547 6217 -7513
rect 6251 -7547 6300 -7513
rect 6100 -7594 6300 -7547
rect 6358 -7513 6558 -7497
rect 6358 -7547 6407 -7513
rect 6441 -7547 6475 -7513
rect 6509 -7547 6558 -7513
rect 6358 -7594 6558 -7547
rect 6616 -7513 6816 -7497
rect 6616 -7547 6665 -7513
rect 6699 -7547 6733 -7513
rect 6767 -7547 6816 -7513
rect 6616 -7594 6816 -7547
rect 7068 -7513 7268 -7497
rect 7068 -7547 7117 -7513
rect 7151 -7547 7185 -7513
rect 7219 -7547 7268 -7513
rect 7068 -7594 7268 -7547
rect 7326 -7513 7526 -7497
rect 7326 -7547 7375 -7513
rect 7409 -7547 7443 -7513
rect 7477 -7547 7526 -7513
rect 7326 -7594 7526 -7547
rect 7584 -7513 7784 -7497
rect 7584 -7547 7633 -7513
rect 7667 -7547 7701 -7513
rect 7735 -7547 7784 -7513
rect 7584 -7594 7784 -7547
rect 8036 -7513 8236 -7497
rect 8036 -7547 8085 -7513
rect 8119 -7547 8153 -7513
rect 8187 -7547 8236 -7513
rect 8036 -7594 8236 -7547
rect 8294 -7513 8494 -7497
rect 8294 -7547 8343 -7513
rect 8377 -7547 8411 -7513
rect 8445 -7547 8494 -7513
rect 8294 -7594 8494 -7547
rect 8552 -7513 8752 -7497
rect 8552 -7547 8601 -7513
rect 8635 -7547 8669 -7513
rect 8703 -7547 8752 -7513
rect 8552 -7594 8752 -7547
rect 8810 -7513 9010 -7497
rect 8810 -7547 8859 -7513
rect 8893 -7547 8927 -7513
rect 8961 -7547 9010 -7513
rect 8810 -7594 9010 -7547
rect 9262 -7513 9462 -7497
rect 9262 -7547 9311 -7513
rect 9345 -7547 9379 -7513
rect 9413 -7547 9462 -7513
rect 9262 -7594 9462 -7547
rect 1033 -7820 1233 -7794
rect 1485 -7820 1685 -7794
rect 1743 -7820 1943 -7794
rect 2001 -7820 2201 -7794
rect 2259 -7820 2459 -7794
rect 2711 -7820 2911 -7794
rect 2969 -7820 3169 -7794
rect 3227 -7820 3427 -7794
rect 3679 -7820 3879 -7794
rect 3937 -7820 4137 -7794
rect 4195 -7820 4395 -7794
rect 4453 -7820 4653 -7794
rect 4905 -7820 5105 -7794
rect 5391 -7820 5591 -7794
rect 5842 -7820 6042 -7794
rect 6100 -7820 6300 -7794
rect 6358 -7820 6558 -7794
rect 6616 -7820 6816 -7794
rect 7068 -7820 7268 -7794
rect 7326 -7820 7526 -7794
rect 7584 -7820 7784 -7794
rect 8036 -7820 8236 -7794
rect 8294 -7820 8494 -7794
rect 8552 -7820 8752 -7794
rect 8810 -7820 9010 -7794
rect 9262 -7820 9462 -7794
rect 1033 -8538 1233 -8512
rect 1485 -8538 1685 -8512
rect 1743 -8538 1943 -8512
rect 2001 -8538 2201 -8512
rect 2259 -8538 2459 -8512
rect 2711 -8538 2911 -8512
rect 2969 -8538 3169 -8512
rect 3227 -8538 3427 -8512
rect 3679 -8538 3879 -8512
rect 3937 -8538 4137 -8512
rect 4195 -8538 4395 -8512
rect 4453 -8538 4653 -8512
rect 4905 -8538 5105 -8512
rect 5391 -8538 5591 -8512
rect 5842 -8538 6042 -8512
rect 6100 -8538 6300 -8512
rect 6358 -8538 6558 -8512
rect 6616 -8538 6816 -8512
rect 7068 -8538 7268 -8512
rect 7326 -8538 7526 -8512
rect 7584 -8538 7784 -8512
rect 8036 -8538 8236 -8512
rect 8294 -8538 8494 -8512
rect 8552 -8538 8752 -8512
rect 8810 -8538 9010 -8512
rect 9262 -8538 9462 -8512
rect 1033 -8785 1233 -8738
rect 1033 -8819 1082 -8785
rect 1116 -8819 1150 -8785
rect 1184 -8819 1233 -8785
rect 1033 -8835 1233 -8819
rect 1485 -8785 1685 -8738
rect 1485 -8819 1534 -8785
rect 1568 -8819 1602 -8785
rect 1636 -8819 1685 -8785
rect 1485 -8835 1685 -8819
rect 1743 -8785 1943 -8738
rect 1743 -8819 1792 -8785
rect 1826 -8819 1860 -8785
rect 1894 -8819 1943 -8785
rect 1743 -8835 1943 -8819
rect 2001 -8785 2201 -8738
rect 2001 -8819 2050 -8785
rect 2084 -8819 2118 -8785
rect 2152 -8819 2201 -8785
rect 2001 -8835 2201 -8819
rect 2259 -8785 2459 -8738
rect 2259 -8819 2308 -8785
rect 2342 -8819 2376 -8785
rect 2410 -8819 2459 -8785
rect 2259 -8835 2459 -8819
rect 2711 -8785 2911 -8738
rect 2711 -8819 2760 -8785
rect 2794 -8819 2828 -8785
rect 2862 -8819 2911 -8785
rect 2711 -8835 2911 -8819
rect 2969 -8785 3169 -8738
rect 2969 -8819 3018 -8785
rect 3052 -8819 3086 -8785
rect 3120 -8819 3169 -8785
rect 2969 -8835 3169 -8819
rect 3227 -8785 3427 -8738
rect 3227 -8819 3276 -8785
rect 3310 -8819 3344 -8785
rect 3378 -8819 3427 -8785
rect 3227 -8835 3427 -8819
rect 3679 -8785 3879 -8738
rect 3679 -8819 3728 -8785
rect 3762 -8819 3796 -8785
rect 3830 -8819 3879 -8785
rect 3679 -8835 3879 -8819
rect 3937 -8785 4137 -8738
rect 3937 -8819 3986 -8785
rect 4020 -8819 4054 -8785
rect 4088 -8819 4137 -8785
rect 3937 -8835 4137 -8819
rect 4195 -8785 4395 -8738
rect 4195 -8819 4244 -8785
rect 4278 -8819 4312 -8785
rect 4346 -8819 4395 -8785
rect 4195 -8835 4395 -8819
rect 4453 -8785 4653 -8738
rect 4453 -8819 4502 -8785
rect 4536 -8819 4570 -8785
rect 4604 -8819 4653 -8785
rect 4453 -8835 4653 -8819
rect 4905 -8785 5105 -8738
rect 4905 -8819 4954 -8785
rect 4988 -8819 5022 -8785
rect 5056 -8819 5105 -8785
rect 4905 -8835 5105 -8819
rect 5391 -8785 5591 -8738
rect 5391 -8819 5440 -8785
rect 5474 -8819 5508 -8785
rect 5542 -8819 5591 -8785
rect 5391 -8835 5591 -8819
rect 5842 -8785 6042 -8738
rect 5842 -8819 5891 -8785
rect 5925 -8819 5959 -8785
rect 5993 -8819 6042 -8785
rect 5842 -8835 6042 -8819
rect 6100 -8785 6300 -8738
rect 6100 -8819 6149 -8785
rect 6183 -8819 6217 -8785
rect 6251 -8819 6300 -8785
rect 6100 -8835 6300 -8819
rect 6358 -8785 6558 -8738
rect 6358 -8819 6407 -8785
rect 6441 -8819 6475 -8785
rect 6509 -8819 6558 -8785
rect 6358 -8835 6558 -8819
rect 6616 -8785 6816 -8738
rect 6616 -8819 6665 -8785
rect 6699 -8819 6733 -8785
rect 6767 -8819 6816 -8785
rect 6616 -8835 6816 -8819
rect 7068 -8785 7268 -8738
rect 7068 -8819 7117 -8785
rect 7151 -8819 7185 -8785
rect 7219 -8819 7268 -8785
rect 7068 -8835 7268 -8819
rect 7326 -8785 7526 -8738
rect 7326 -8819 7375 -8785
rect 7409 -8819 7443 -8785
rect 7477 -8819 7526 -8785
rect 7326 -8835 7526 -8819
rect 7584 -8785 7784 -8738
rect 7584 -8819 7633 -8785
rect 7667 -8819 7701 -8785
rect 7735 -8819 7784 -8785
rect 7584 -8835 7784 -8819
rect 8036 -8785 8236 -8738
rect 8036 -8819 8085 -8785
rect 8119 -8819 8153 -8785
rect 8187 -8819 8236 -8785
rect 8036 -8835 8236 -8819
rect 8294 -8785 8494 -8738
rect 8294 -8819 8343 -8785
rect 8377 -8819 8411 -8785
rect 8445 -8819 8494 -8785
rect 8294 -8835 8494 -8819
rect 8552 -8785 8752 -8738
rect 8552 -8819 8601 -8785
rect 8635 -8819 8669 -8785
rect 8703 -8819 8752 -8785
rect 8552 -8835 8752 -8819
rect 8810 -8785 9010 -8738
rect 8810 -8819 8859 -8785
rect 8893 -8819 8927 -8785
rect 8961 -8819 9010 -8785
rect 8810 -8835 9010 -8819
rect 9262 -8785 9462 -8738
rect 9262 -8819 9311 -8785
rect 9345 -8819 9379 -8785
rect 9413 -8819 9462 -8785
rect 9262 -8835 9462 -8819
<< polycont >>
rect 1082 608 1116 642
rect 1150 608 1184 642
rect 1534 608 1568 642
rect 1602 608 1636 642
rect 1792 608 1826 642
rect 1860 608 1894 642
rect 2050 608 2084 642
rect 2118 608 2152 642
rect 2308 608 2342 642
rect 2376 608 2410 642
rect 2760 608 2794 642
rect 2828 608 2862 642
rect 3018 608 3052 642
rect 3086 608 3120 642
rect 3276 608 3310 642
rect 3344 608 3378 642
rect 3728 608 3762 642
rect 3796 608 3830 642
rect 3986 608 4020 642
rect 4054 608 4088 642
rect 4244 608 4278 642
rect 4312 608 4346 642
rect 4502 608 4536 642
rect 4570 608 4604 642
rect 4954 608 4988 642
rect 5022 608 5056 642
rect 5440 608 5474 642
rect 5508 608 5542 642
rect 5891 608 5925 642
rect 5959 608 5993 642
rect 6149 608 6183 642
rect 6217 608 6251 642
rect 6407 608 6441 642
rect 6475 608 6509 642
rect 6665 608 6699 642
rect 6733 608 6767 642
rect 7117 608 7151 642
rect 7185 608 7219 642
rect 7375 608 7409 642
rect 7443 608 7477 642
rect 7633 608 7667 642
rect 7701 608 7735 642
rect 8085 608 8119 642
rect 8153 608 8187 642
rect 8343 608 8377 642
rect 8411 608 8445 642
rect 8601 608 8635 642
rect 8669 608 8703 642
rect 8859 608 8893 642
rect 8927 608 8961 642
rect 9311 608 9345 642
rect 9379 608 9413 642
rect 1082 -664 1116 -630
rect 1150 -664 1184 -630
rect 1534 -664 1568 -630
rect 1602 -664 1636 -630
rect 1792 -664 1826 -630
rect 1860 -664 1894 -630
rect 2050 -664 2084 -630
rect 2118 -664 2152 -630
rect 2308 -664 2342 -630
rect 2376 -664 2410 -630
rect 2760 -664 2794 -630
rect 2828 -664 2862 -630
rect 3018 -664 3052 -630
rect 3086 -664 3120 -630
rect 3276 -664 3310 -630
rect 3344 -664 3378 -630
rect 3728 -664 3762 -630
rect 3796 -664 3830 -630
rect 3986 -664 4020 -630
rect 4054 -664 4088 -630
rect 4244 -664 4278 -630
rect 4312 -664 4346 -630
rect 4502 -664 4536 -630
rect 4570 -664 4604 -630
rect 4954 -664 4988 -630
rect 5022 -664 5056 -630
rect 5440 -664 5474 -630
rect 5508 -664 5542 -630
rect 5891 -664 5925 -630
rect 5959 -664 5993 -630
rect 6149 -664 6183 -630
rect 6217 -664 6251 -630
rect 6407 -664 6441 -630
rect 6475 -664 6509 -630
rect 6665 -664 6699 -630
rect 6733 -664 6767 -630
rect 7117 -664 7151 -630
rect 7185 -664 7219 -630
rect 7375 -664 7409 -630
rect 7443 -664 7477 -630
rect 7633 -664 7667 -630
rect 7701 -664 7735 -630
rect 8085 -664 8119 -630
rect 8153 -664 8187 -630
rect 8343 -664 8377 -630
rect 8411 -664 8445 -630
rect 8601 -664 8635 -630
rect 8669 -664 8703 -630
rect 8859 -664 8893 -630
rect 8927 -664 8961 -630
rect 9311 -664 9345 -630
rect 9379 -664 9413 -630
rect 1082 -1027 1116 -993
rect 1150 -1027 1184 -993
rect 1534 -1027 1568 -993
rect 1602 -1027 1636 -993
rect 1792 -1027 1826 -993
rect 1860 -1027 1894 -993
rect 2050 -1027 2084 -993
rect 2118 -1027 2152 -993
rect 2308 -1027 2342 -993
rect 2376 -1027 2410 -993
rect 2760 -1027 2794 -993
rect 2828 -1027 2862 -993
rect 3018 -1027 3052 -993
rect 3086 -1027 3120 -993
rect 3276 -1027 3310 -993
rect 3344 -1027 3378 -993
rect 3728 -1027 3762 -993
rect 3796 -1027 3830 -993
rect 3986 -1027 4020 -993
rect 4054 -1027 4088 -993
rect 4244 -1027 4278 -993
rect 4312 -1027 4346 -993
rect 4502 -1027 4536 -993
rect 4570 -1027 4604 -993
rect 4954 -1027 4988 -993
rect 5022 -1027 5056 -993
rect 5440 -1027 5474 -993
rect 5508 -1027 5542 -993
rect 5891 -1027 5925 -993
rect 5959 -1027 5993 -993
rect 6149 -1027 6183 -993
rect 6217 -1027 6251 -993
rect 6407 -1027 6441 -993
rect 6475 -1027 6509 -993
rect 6665 -1027 6699 -993
rect 6733 -1027 6767 -993
rect 7117 -1027 7151 -993
rect 7185 -1027 7219 -993
rect 7375 -1027 7409 -993
rect 7443 -1027 7477 -993
rect 7633 -1027 7667 -993
rect 7701 -1027 7735 -993
rect 8085 -1027 8119 -993
rect 8153 -1027 8187 -993
rect 8343 -1027 8377 -993
rect 8411 -1027 8445 -993
rect 8601 -1027 8635 -993
rect 8669 -1027 8703 -993
rect 8859 -1027 8893 -993
rect 8927 -1027 8961 -993
rect 9311 -1027 9345 -993
rect 9379 -1027 9413 -993
rect 1082 -2311 1116 -2277
rect 1150 -2311 1184 -2277
rect 1534 -2311 1568 -2277
rect 1602 -2311 1636 -2277
rect 1792 -2311 1826 -2277
rect 1860 -2311 1894 -2277
rect 2050 -2311 2084 -2277
rect 2118 -2311 2152 -2277
rect 2308 -2311 2342 -2277
rect 2376 -2311 2410 -2277
rect 2760 -2311 2794 -2277
rect 2828 -2311 2862 -2277
rect 3018 -2311 3052 -2277
rect 3086 -2311 3120 -2277
rect 3276 -2311 3310 -2277
rect 3344 -2311 3378 -2277
rect 3728 -2311 3762 -2277
rect 3796 -2311 3830 -2277
rect 3986 -2311 4020 -2277
rect 4054 -2311 4088 -2277
rect 4244 -2311 4278 -2277
rect 4312 -2311 4346 -2277
rect 4502 -2311 4536 -2277
rect 4570 -2311 4604 -2277
rect 4954 -2311 4988 -2277
rect 5022 -2311 5056 -2277
rect 5440 -2311 5474 -2277
rect 5508 -2311 5542 -2277
rect 5891 -2311 5925 -2277
rect 5959 -2311 5993 -2277
rect 6149 -2311 6183 -2277
rect 6217 -2311 6251 -2277
rect 6407 -2311 6441 -2277
rect 6475 -2311 6509 -2277
rect 6665 -2311 6699 -2277
rect 6733 -2311 6767 -2277
rect 7117 -2311 7151 -2277
rect 7185 -2311 7219 -2277
rect 7375 -2311 7409 -2277
rect 7443 -2311 7477 -2277
rect 7633 -2311 7667 -2277
rect 7701 -2311 7735 -2277
rect 8085 -2311 8119 -2277
rect 8153 -2311 8187 -2277
rect 8343 -2311 8377 -2277
rect 8411 -2311 8445 -2277
rect 8601 -2311 8635 -2277
rect 8669 -2311 8703 -2277
rect 8859 -2311 8893 -2277
rect 8927 -2311 8961 -2277
rect 9311 -2311 9345 -2277
rect 9379 -2311 9413 -2277
rect 1082 -2674 1116 -2640
rect 1150 -2674 1184 -2640
rect 1534 -2674 1568 -2640
rect 1602 -2674 1636 -2640
rect 1792 -2674 1826 -2640
rect 1860 -2674 1894 -2640
rect 2050 -2674 2084 -2640
rect 2118 -2674 2152 -2640
rect 2308 -2674 2342 -2640
rect 2376 -2674 2410 -2640
rect 2760 -2674 2794 -2640
rect 2828 -2674 2862 -2640
rect 3018 -2674 3052 -2640
rect 3086 -2674 3120 -2640
rect 3276 -2674 3310 -2640
rect 3344 -2674 3378 -2640
rect 3728 -2674 3762 -2640
rect 3796 -2674 3830 -2640
rect 3986 -2674 4020 -2640
rect 4054 -2674 4088 -2640
rect 4244 -2674 4278 -2640
rect 4312 -2674 4346 -2640
rect 4502 -2674 4536 -2640
rect 4570 -2674 4604 -2640
rect 4954 -2674 4988 -2640
rect 5022 -2674 5056 -2640
rect 5440 -2674 5474 -2640
rect 5508 -2674 5542 -2640
rect 5891 -2674 5925 -2640
rect 5959 -2674 5993 -2640
rect 6149 -2674 6183 -2640
rect 6217 -2674 6251 -2640
rect 6407 -2674 6441 -2640
rect 6475 -2674 6509 -2640
rect 6665 -2674 6699 -2640
rect 6733 -2674 6767 -2640
rect 7117 -2674 7151 -2640
rect 7185 -2674 7219 -2640
rect 7375 -2674 7409 -2640
rect 7443 -2674 7477 -2640
rect 7633 -2674 7667 -2640
rect 7701 -2674 7735 -2640
rect 8085 -2674 8119 -2640
rect 8153 -2674 8187 -2640
rect 8343 -2674 8377 -2640
rect 8411 -2674 8445 -2640
rect 8601 -2674 8635 -2640
rect 8669 -2674 8703 -2640
rect 8859 -2674 8893 -2640
rect 8927 -2674 8961 -2640
rect 9311 -2674 9345 -2640
rect 9379 -2674 9413 -2640
rect 1082 -3992 1116 -3958
rect 1150 -3992 1184 -3958
rect 1534 -3992 1568 -3958
rect 1602 -3992 1636 -3958
rect 1792 -3992 1826 -3958
rect 1860 -3992 1894 -3958
rect 2050 -3992 2084 -3958
rect 2118 -3992 2152 -3958
rect 2308 -3992 2342 -3958
rect 2376 -3992 2410 -3958
rect 2760 -3992 2794 -3958
rect 2828 -3992 2862 -3958
rect 3018 -3992 3052 -3958
rect 3086 -3992 3120 -3958
rect 3276 -3992 3310 -3958
rect 3344 -3992 3378 -3958
rect 3728 -3992 3762 -3958
rect 3796 -3992 3830 -3958
rect 3986 -3992 4020 -3958
rect 4054 -3992 4088 -3958
rect 4244 -3992 4278 -3958
rect 4312 -3992 4346 -3958
rect 4502 -3992 4536 -3958
rect 4570 -3992 4604 -3958
rect 4954 -3992 4988 -3958
rect 5022 -3992 5056 -3958
rect 5440 -3992 5474 -3958
rect 5508 -3992 5542 -3958
rect 5891 -3992 5925 -3958
rect 5959 -3992 5993 -3958
rect 6149 -3992 6183 -3958
rect 6217 -3992 6251 -3958
rect 6407 -3992 6441 -3958
rect 6475 -3992 6509 -3958
rect 6665 -3992 6699 -3958
rect 6733 -3992 6767 -3958
rect 7117 -3992 7151 -3958
rect 7185 -3992 7219 -3958
rect 7375 -3992 7409 -3958
rect 7443 -3992 7477 -3958
rect 7633 -3992 7667 -3958
rect 7701 -3992 7735 -3958
rect 8085 -3992 8119 -3958
rect 8153 -3992 8187 -3958
rect 8343 -3992 8377 -3958
rect 8411 -3992 8445 -3958
rect 8601 -3992 8635 -3958
rect 8669 -3992 8703 -3958
rect 8859 -3992 8893 -3958
rect 8927 -3992 8961 -3958
rect 9311 -3992 9345 -3958
rect 9379 -3992 9413 -3958
rect 1082 -4220 1116 -4186
rect 1150 -4220 1184 -4186
rect 1534 -4220 1568 -4186
rect 1602 -4220 1636 -4186
rect 1792 -4220 1826 -4186
rect 1860 -4220 1894 -4186
rect 2050 -4220 2084 -4186
rect 2118 -4220 2152 -4186
rect 2308 -4220 2342 -4186
rect 2376 -4220 2410 -4186
rect 2760 -4220 2794 -4186
rect 2828 -4220 2862 -4186
rect 3018 -4220 3052 -4186
rect 3086 -4220 3120 -4186
rect 3276 -4220 3310 -4186
rect 3344 -4220 3378 -4186
rect 3728 -4220 3762 -4186
rect 3796 -4220 3830 -4186
rect 3986 -4220 4020 -4186
rect 4054 -4220 4088 -4186
rect 4244 -4220 4278 -4186
rect 4312 -4220 4346 -4186
rect 4502 -4220 4536 -4186
rect 4570 -4220 4604 -4186
rect 4954 -4220 4988 -4186
rect 5022 -4220 5056 -4186
rect 5440 -4220 5474 -4186
rect 5508 -4220 5542 -4186
rect 5891 -4220 5925 -4186
rect 5959 -4220 5993 -4186
rect 6149 -4220 6183 -4186
rect 6217 -4220 6251 -4186
rect 6407 -4220 6441 -4186
rect 6475 -4220 6509 -4186
rect 6665 -4220 6699 -4186
rect 6733 -4220 6767 -4186
rect 7117 -4220 7151 -4186
rect 7185 -4220 7219 -4186
rect 7375 -4220 7409 -4186
rect 7443 -4220 7477 -4186
rect 7633 -4220 7667 -4186
rect 7701 -4220 7735 -4186
rect 8085 -4220 8119 -4186
rect 8153 -4220 8187 -4186
rect 8343 -4220 8377 -4186
rect 8411 -4220 8445 -4186
rect 8601 -4220 8635 -4186
rect 8669 -4220 8703 -4186
rect 8859 -4220 8893 -4186
rect 8927 -4220 8961 -4186
rect 9311 -4220 9345 -4186
rect 9379 -4220 9413 -4186
rect 1082 -5538 1116 -5504
rect 1150 -5538 1184 -5504
rect 1534 -5538 1568 -5504
rect 1602 -5538 1636 -5504
rect 1792 -5538 1826 -5504
rect 1860 -5538 1894 -5504
rect 2050 -5538 2084 -5504
rect 2118 -5538 2152 -5504
rect 2308 -5538 2342 -5504
rect 2376 -5538 2410 -5504
rect 2760 -5538 2794 -5504
rect 2828 -5538 2862 -5504
rect 3018 -5538 3052 -5504
rect 3086 -5538 3120 -5504
rect 3276 -5538 3310 -5504
rect 3344 -5538 3378 -5504
rect 3728 -5538 3762 -5504
rect 3796 -5538 3830 -5504
rect 3986 -5538 4020 -5504
rect 4054 -5538 4088 -5504
rect 4244 -5538 4278 -5504
rect 4312 -5538 4346 -5504
rect 4502 -5538 4536 -5504
rect 4570 -5538 4604 -5504
rect 4954 -5538 4988 -5504
rect 5022 -5538 5056 -5504
rect 5440 -5538 5474 -5504
rect 5508 -5538 5542 -5504
rect 5891 -5538 5925 -5504
rect 5959 -5538 5993 -5504
rect 6149 -5538 6183 -5504
rect 6217 -5538 6251 -5504
rect 6407 -5538 6441 -5504
rect 6475 -5538 6509 -5504
rect 6665 -5538 6699 -5504
rect 6733 -5538 6767 -5504
rect 7117 -5538 7151 -5504
rect 7185 -5538 7219 -5504
rect 7375 -5538 7409 -5504
rect 7443 -5538 7477 -5504
rect 7633 -5538 7667 -5504
rect 7701 -5538 7735 -5504
rect 8085 -5538 8119 -5504
rect 8153 -5538 8187 -5504
rect 8343 -5538 8377 -5504
rect 8411 -5538 8445 -5504
rect 8601 -5538 8635 -5504
rect 8669 -5538 8703 -5504
rect 8859 -5538 8893 -5504
rect 8927 -5538 8961 -5504
rect 9311 -5538 9345 -5504
rect 9379 -5538 9413 -5504
rect 1082 -5900 1116 -5866
rect 1150 -5900 1184 -5866
rect 1534 -5900 1568 -5866
rect 1602 -5900 1636 -5866
rect 1792 -5900 1826 -5866
rect 1860 -5900 1894 -5866
rect 2050 -5900 2084 -5866
rect 2118 -5900 2152 -5866
rect 2308 -5900 2342 -5866
rect 2376 -5900 2410 -5866
rect 2760 -5900 2794 -5866
rect 2828 -5900 2862 -5866
rect 3018 -5900 3052 -5866
rect 3086 -5900 3120 -5866
rect 3276 -5900 3310 -5866
rect 3344 -5900 3378 -5866
rect 3728 -5900 3762 -5866
rect 3796 -5900 3830 -5866
rect 3986 -5900 4020 -5866
rect 4054 -5900 4088 -5866
rect 4244 -5900 4278 -5866
rect 4312 -5900 4346 -5866
rect 4502 -5900 4536 -5866
rect 4570 -5900 4604 -5866
rect 4954 -5900 4988 -5866
rect 5022 -5900 5056 -5866
rect 5440 -5900 5474 -5866
rect 5508 -5900 5542 -5866
rect 5891 -5900 5925 -5866
rect 5959 -5900 5993 -5866
rect 6149 -5900 6183 -5866
rect 6217 -5900 6251 -5866
rect 6407 -5900 6441 -5866
rect 6475 -5900 6509 -5866
rect 6665 -5900 6699 -5866
rect 6733 -5900 6767 -5866
rect 7117 -5900 7151 -5866
rect 7185 -5900 7219 -5866
rect 7375 -5900 7409 -5866
rect 7443 -5900 7477 -5866
rect 7633 -5900 7667 -5866
rect 7701 -5900 7735 -5866
rect 8085 -5900 8119 -5866
rect 8153 -5900 8187 -5866
rect 8343 -5900 8377 -5866
rect 8411 -5900 8445 -5866
rect 8601 -5900 8635 -5866
rect 8669 -5900 8703 -5866
rect 8859 -5900 8893 -5866
rect 8927 -5900 8961 -5866
rect 9311 -5900 9345 -5866
rect 9379 -5900 9413 -5866
rect 1082 -7185 1116 -7151
rect 1150 -7185 1184 -7151
rect 1534 -7185 1568 -7151
rect 1602 -7185 1636 -7151
rect 1792 -7185 1826 -7151
rect 1860 -7185 1894 -7151
rect 2050 -7185 2084 -7151
rect 2118 -7185 2152 -7151
rect 2308 -7185 2342 -7151
rect 2376 -7185 2410 -7151
rect 2760 -7185 2794 -7151
rect 2828 -7185 2862 -7151
rect 3018 -7185 3052 -7151
rect 3086 -7185 3120 -7151
rect 3276 -7185 3310 -7151
rect 3344 -7185 3378 -7151
rect 3728 -7185 3762 -7151
rect 3796 -7185 3830 -7151
rect 3986 -7185 4020 -7151
rect 4054 -7185 4088 -7151
rect 4244 -7185 4278 -7151
rect 4312 -7185 4346 -7151
rect 4502 -7185 4536 -7151
rect 4570 -7185 4604 -7151
rect 4954 -7185 4988 -7151
rect 5022 -7185 5056 -7151
rect 5440 -7185 5474 -7151
rect 5508 -7185 5542 -7151
rect 5891 -7185 5925 -7151
rect 5959 -7185 5993 -7151
rect 6149 -7185 6183 -7151
rect 6217 -7185 6251 -7151
rect 6407 -7185 6441 -7151
rect 6475 -7185 6509 -7151
rect 6665 -7185 6699 -7151
rect 6733 -7185 6767 -7151
rect 7117 -7185 7151 -7151
rect 7185 -7185 7219 -7151
rect 7375 -7185 7409 -7151
rect 7443 -7185 7477 -7151
rect 7633 -7185 7667 -7151
rect 7701 -7185 7735 -7151
rect 8085 -7185 8119 -7151
rect 8153 -7185 8187 -7151
rect 8343 -7185 8377 -7151
rect 8411 -7185 8445 -7151
rect 8601 -7185 8635 -7151
rect 8669 -7185 8703 -7151
rect 8859 -7185 8893 -7151
rect 8927 -7185 8961 -7151
rect 9311 -7185 9345 -7151
rect 9379 -7185 9413 -7151
rect 1082 -7547 1116 -7513
rect 1150 -7547 1184 -7513
rect 1534 -7547 1568 -7513
rect 1602 -7547 1636 -7513
rect 1792 -7547 1826 -7513
rect 1860 -7547 1894 -7513
rect 2050 -7547 2084 -7513
rect 2118 -7547 2152 -7513
rect 2308 -7547 2342 -7513
rect 2376 -7547 2410 -7513
rect 2760 -7547 2794 -7513
rect 2828 -7547 2862 -7513
rect 3018 -7547 3052 -7513
rect 3086 -7547 3120 -7513
rect 3276 -7547 3310 -7513
rect 3344 -7547 3378 -7513
rect 3728 -7547 3762 -7513
rect 3796 -7547 3830 -7513
rect 3986 -7547 4020 -7513
rect 4054 -7547 4088 -7513
rect 4244 -7547 4278 -7513
rect 4312 -7547 4346 -7513
rect 4502 -7547 4536 -7513
rect 4570 -7547 4604 -7513
rect 4954 -7547 4988 -7513
rect 5022 -7547 5056 -7513
rect 5440 -7547 5474 -7513
rect 5508 -7547 5542 -7513
rect 5891 -7547 5925 -7513
rect 5959 -7547 5993 -7513
rect 6149 -7547 6183 -7513
rect 6217 -7547 6251 -7513
rect 6407 -7547 6441 -7513
rect 6475 -7547 6509 -7513
rect 6665 -7547 6699 -7513
rect 6733 -7547 6767 -7513
rect 7117 -7547 7151 -7513
rect 7185 -7547 7219 -7513
rect 7375 -7547 7409 -7513
rect 7443 -7547 7477 -7513
rect 7633 -7547 7667 -7513
rect 7701 -7547 7735 -7513
rect 8085 -7547 8119 -7513
rect 8153 -7547 8187 -7513
rect 8343 -7547 8377 -7513
rect 8411 -7547 8445 -7513
rect 8601 -7547 8635 -7513
rect 8669 -7547 8703 -7513
rect 8859 -7547 8893 -7513
rect 8927 -7547 8961 -7513
rect 9311 -7547 9345 -7513
rect 9379 -7547 9413 -7513
rect 1082 -8819 1116 -8785
rect 1150 -8819 1184 -8785
rect 1534 -8819 1568 -8785
rect 1602 -8819 1636 -8785
rect 1792 -8819 1826 -8785
rect 1860 -8819 1894 -8785
rect 2050 -8819 2084 -8785
rect 2118 -8819 2152 -8785
rect 2308 -8819 2342 -8785
rect 2376 -8819 2410 -8785
rect 2760 -8819 2794 -8785
rect 2828 -8819 2862 -8785
rect 3018 -8819 3052 -8785
rect 3086 -8819 3120 -8785
rect 3276 -8819 3310 -8785
rect 3344 -8819 3378 -8785
rect 3728 -8819 3762 -8785
rect 3796 -8819 3830 -8785
rect 3986 -8819 4020 -8785
rect 4054 -8819 4088 -8785
rect 4244 -8819 4278 -8785
rect 4312 -8819 4346 -8785
rect 4502 -8819 4536 -8785
rect 4570 -8819 4604 -8785
rect 4954 -8819 4988 -8785
rect 5022 -8819 5056 -8785
rect 5440 -8819 5474 -8785
rect 5508 -8819 5542 -8785
rect 5891 -8819 5925 -8785
rect 5959 -8819 5993 -8785
rect 6149 -8819 6183 -8785
rect 6217 -8819 6251 -8785
rect 6407 -8819 6441 -8785
rect 6475 -8819 6509 -8785
rect 6665 -8819 6699 -8785
rect 6733 -8819 6767 -8785
rect 7117 -8819 7151 -8785
rect 7185 -8819 7219 -8785
rect 7375 -8819 7409 -8785
rect 7443 -8819 7477 -8785
rect 7633 -8819 7667 -8785
rect 7701 -8819 7735 -8785
rect 8085 -8819 8119 -8785
rect 8153 -8819 8187 -8785
rect 8343 -8819 8377 -8785
rect 8411 -8819 8445 -8785
rect 8601 -8819 8635 -8785
rect 8669 -8819 8703 -8785
rect 8859 -8819 8893 -8785
rect 8927 -8819 8961 -8785
rect 9311 -8819 9345 -8785
rect 9379 -8819 9413 -8785
<< locali >>
rect 872 722 946 756
rect 980 722 993 756
rect 1052 722 1061 756
rect 1124 722 1129 756
rect 1196 722 1197 756
rect 1231 722 1234 756
rect 1299 722 1306 756
rect 1367 722 1378 756
rect 1435 722 1450 756
rect 1503 722 1522 756
rect 1571 722 1594 756
rect 1639 722 1666 756
rect 1707 722 1738 756
rect 1775 722 1809 756
rect 1844 722 1877 756
rect 1916 722 1945 756
rect 1988 722 2013 756
rect 2060 722 2081 756
rect 2132 722 2149 756
rect 2204 722 2217 756
rect 2276 722 2285 756
rect 2348 722 2353 756
rect 2420 722 2421 756
rect 2455 722 2458 756
rect 2523 722 2530 756
rect 2591 722 2602 756
rect 2659 722 2674 756
rect 2727 722 2746 756
rect 2795 722 2818 756
rect 2863 722 2890 756
rect 2931 722 2962 756
rect 2999 722 3033 756
rect 3068 722 3101 756
rect 3140 722 3169 756
rect 3212 722 3237 756
rect 3284 722 3305 756
rect 3356 722 3373 756
rect 3428 722 3441 756
rect 3500 722 3509 756
rect 3572 722 3577 756
rect 3644 722 3645 756
rect 3679 722 3682 756
rect 3747 722 3754 756
rect 3815 722 3826 756
rect 3883 722 3898 756
rect 3951 722 3970 756
rect 4019 722 4042 756
rect 4087 722 4114 756
rect 4155 722 4186 756
rect 4223 722 4257 756
rect 4292 722 4325 756
rect 4364 722 4393 756
rect 4436 722 4461 756
rect 4508 722 4529 756
rect 4580 722 4597 756
rect 4652 722 4665 756
rect 4724 722 4733 756
rect 4796 722 4801 756
rect 4868 722 4869 756
rect 4903 722 4906 756
rect 4971 722 4978 756
rect 5039 722 5050 756
rect 5107 722 5122 756
rect 5156 722 5339 756
rect 5373 722 5388 756
rect 5445 722 5456 756
rect 5517 722 5524 756
rect 5589 722 5592 756
rect 5626 722 5627 756
rect 5694 722 5699 756
rect 5762 722 5771 756
rect 5830 722 5843 756
rect 5898 722 5915 756
rect 5966 722 5987 756
rect 6034 722 6059 756
rect 6102 722 6131 756
rect 6170 722 6203 756
rect 6238 722 6272 756
rect 6309 722 6340 756
rect 6381 722 6408 756
rect 6453 722 6476 756
rect 6525 722 6544 756
rect 6597 722 6612 756
rect 6669 722 6680 756
rect 6741 722 6748 756
rect 6813 722 6816 756
rect 6850 722 6851 756
rect 6918 722 6923 756
rect 6986 722 6995 756
rect 7054 722 7067 756
rect 7122 722 7139 756
rect 7190 722 7211 756
rect 7258 722 7283 756
rect 7326 722 7355 756
rect 7394 722 7427 756
rect 7462 722 7496 756
rect 7533 722 7564 756
rect 7605 722 7632 756
rect 7677 722 7700 756
rect 7749 722 7768 756
rect 7821 722 7836 756
rect 7893 722 7904 756
rect 7965 722 7972 756
rect 8037 722 8040 756
rect 8074 722 8075 756
rect 8142 722 8147 756
rect 8210 722 8219 756
rect 8278 722 8291 756
rect 8346 722 8363 756
rect 8414 722 8435 756
rect 8482 722 8507 756
rect 8550 722 8579 756
rect 8618 722 8651 756
rect 8686 722 8720 756
rect 8757 722 8788 756
rect 8829 722 8856 756
rect 8901 722 8924 756
rect 8973 722 8992 756
rect 9045 722 9060 756
rect 9117 722 9128 756
rect 9189 722 9196 756
rect 9261 722 9264 756
rect 9298 722 9299 756
rect 9366 722 9371 756
rect 9434 722 9443 756
rect 9502 722 9515 756
rect 9549 722 9623 756
rect 872 599 906 722
rect 1033 608 1080 642
rect 1116 608 1150 642
rect 1186 608 1233 642
rect 1485 608 1532 642
rect 1568 608 1602 642
rect 1638 608 1685 642
rect 1743 608 1790 642
rect 1826 608 1860 642
rect 1896 608 1943 642
rect 2001 608 2048 642
rect 2084 608 2118 642
rect 2154 608 2201 642
rect 2259 608 2306 642
rect 2342 608 2376 642
rect 2412 608 2459 642
rect 2711 608 2758 642
rect 2794 608 2828 642
rect 2864 608 2911 642
rect 2969 608 3016 642
rect 3052 608 3086 642
rect 3122 608 3169 642
rect 3227 608 3274 642
rect 3310 608 3344 642
rect 3380 608 3427 642
rect 3679 608 3726 642
rect 3762 608 3796 642
rect 3832 608 3879 642
rect 3937 608 3984 642
rect 4020 608 4054 642
rect 4090 608 4137 642
rect 4195 608 4242 642
rect 4278 608 4312 642
rect 4348 608 4395 642
rect 4453 608 4500 642
rect 4536 608 4570 642
rect 4606 608 4653 642
rect 4905 608 4952 642
rect 4988 608 5022 642
rect 5058 608 5105 642
rect 5230 599 5265 722
rect 5391 608 5438 642
rect 5474 608 5508 642
rect 5544 608 5591 642
rect 5842 608 5889 642
rect 5925 608 5959 642
rect 5995 608 6042 642
rect 6100 608 6147 642
rect 6183 608 6217 642
rect 6253 608 6300 642
rect 6358 608 6405 642
rect 6441 608 6475 642
rect 6511 608 6558 642
rect 6616 608 6663 642
rect 6699 608 6733 642
rect 6769 608 6816 642
rect 7068 608 7115 642
rect 7151 608 7185 642
rect 7221 608 7268 642
rect 7326 608 7373 642
rect 7409 608 7443 642
rect 7479 608 7526 642
rect 7584 608 7631 642
rect 7667 608 7701 642
rect 7737 608 7784 642
rect 8036 608 8083 642
rect 8119 608 8153 642
rect 8189 608 8236 642
rect 8294 608 8341 642
rect 8377 608 8411 642
rect 8447 608 8494 642
rect 8552 608 8599 642
rect 8635 608 8669 642
rect 8705 608 8752 642
rect 8810 608 8857 642
rect 8893 608 8927 642
rect 8963 608 9010 642
rect 9262 608 9309 642
rect 9345 608 9379 642
rect 9415 608 9462 642
rect 5230 565 5231 599
rect 9589 599 9623 722
rect 872 543 906 565
rect 872 475 906 493
rect 872 407 906 421
rect 987 546 1021 565
rect 987 478 1021 480
rect 987 442 1021 444
rect 987 357 1021 376
rect 1245 546 1279 565
rect 1245 478 1279 480
rect 1245 442 1279 444
rect 1245 357 1279 376
rect 1439 546 1473 565
rect 1439 478 1473 480
rect 1439 442 1473 444
rect 1439 357 1473 376
rect 1697 546 1731 565
rect 1697 478 1731 480
rect 1697 442 1731 444
rect 1697 357 1731 376
rect 1955 546 1989 565
rect 1955 478 1989 480
rect 1955 442 1989 444
rect 1955 357 1989 376
rect 2213 546 2247 565
rect 2213 478 2247 480
rect 2213 442 2247 444
rect 2213 357 2247 376
rect 2471 546 2505 565
rect 2471 478 2505 480
rect 2471 442 2505 444
rect 2471 357 2505 376
rect 2665 546 2699 565
rect 2665 478 2699 480
rect 2665 442 2699 444
rect 2665 357 2699 376
rect 2923 546 2957 565
rect 2923 478 2957 480
rect 2923 442 2957 444
rect 2923 357 2957 376
rect 3181 546 3215 565
rect 3181 478 3215 480
rect 3181 442 3215 444
rect 3181 357 3215 376
rect 3439 546 3473 565
rect 3439 478 3473 480
rect 3439 442 3473 444
rect 3439 357 3473 376
rect 3633 546 3667 565
rect 3633 478 3667 480
rect 3633 442 3667 444
rect 3633 357 3667 376
rect 3891 546 3925 565
rect 3891 478 3925 480
rect 3891 442 3925 444
rect 3891 357 3925 376
rect 4149 546 4183 565
rect 4149 478 4183 480
rect 4149 442 4183 444
rect 4149 357 4183 376
rect 4407 546 4441 565
rect 4407 478 4441 480
rect 4407 442 4441 444
rect 4407 357 4441 376
rect 4665 546 4699 565
rect 4665 478 4699 480
rect 4665 442 4699 444
rect 4665 357 4699 376
rect 4859 546 4893 565
rect 4859 478 4893 480
rect 4859 442 4893 444
rect 4859 357 4893 376
rect 5117 546 5151 565
rect 5117 478 5151 480
rect 5117 442 5151 444
rect 5117 357 5151 376
rect 5230 543 5265 565
rect 5230 493 5231 543
rect 5230 475 5265 493
rect 5230 421 5231 475
rect 5230 407 5265 421
rect 872 339 906 349
rect 872 271 906 277
rect 872 203 906 205
rect 872 167 906 169
rect 872 95 906 101
rect 872 23 906 33
rect 5230 349 5231 407
rect 5345 546 5379 565
rect 5345 478 5379 480
rect 5345 442 5379 444
rect 5345 357 5379 376
rect 5603 546 5637 565
rect 5603 478 5637 480
rect 5603 442 5637 444
rect 5603 357 5637 376
rect 5796 546 5830 565
rect 5796 478 5830 480
rect 5796 442 5830 444
rect 5796 357 5830 376
rect 6054 546 6088 565
rect 6054 478 6088 480
rect 6054 442 6088 444
rect 6054 357 6088 376
rect 6312 546 6346 565
rect 6312 478 6346 480
rect 6312 442 6346 444
rect 6312 357 6346 376
rect 6570 546 6604 565
rect 6570 478 6604 480
rect 6570 442 6604 444
rect 6570 357 6604 376
rect 6828 546 6862 565
rect 6828 478 6862 480
rect 6828 442 6862 444
rect 6828 357 6862 376
rect 7022 546 7056 565
rect 7022 478 7056 480
rect 7022 442 7056 444
rect 7022 357 7056 376
rect 7280 546 7314 565
rect 7280 478 7314 480
rect 7280 442 7314 444
rect 7280 357 7314 376
rect 7538 546 7572 565
rect 7538 478 7572 480
rect 7538 442 7572 444
rect 7538 357 7572 376
rect 7796 546 7830 565
rect 7796 478 7830 480
rect 7796 442 7830 444
rect 7796 357 7830 376
rect 7990 546 8024 565
rect 7990 478 8024 480
rect 7990 442 8024 444
rect 7990 357 8024 376
rect 8248 546 8282 565
rect 8248 478 8282 480
rect 8248 442 8282 444
rect 8248 357 8282 376
rect 8506 546 8540 565
rect 8506 478 8540 480
rect 8506 442 8540 444
rect 8506 357 8540 376
rect 8764 546 8798 565
rect 8764 478 8798 480
rect 8764 442 8798 444
rect 8764 357 8798 376
rect 9022 546 9056 565
rect 9022 478 9056 480
rect 9022 442 9056 444
rect 9022 357 9056 376
rect 9216 546 9250 565
rect 9216 478 9250 480
rect 9216 442 9250 444
rect 9216 357 9250 376
rect 9474 546 9508 565
rect 9474 478 9508 480
rect 9474 442 9508 444
rect 9474 357 9508 376
rect 9589 543 9623 565
rect 9589 475 9623 493
rect 9589 407 9623 421
rect 5230 339 5265 349
rect 5230 277 5231 339
rect 5230 271 5265 277
rect 5230 205 5231 271
rect 5230 203 5265 205
rect 5230 169 5231 203
rect 5230 167 5265 169
rect 5230 101 5231 167
rect 5230 95 5265 101
rect 5230 33 5231 95
rect 5230 23 5265 33
rect 5230 -35 5231 23
rect 9589 339 9623 349
rect 9589 271 9623 277
rect 9589 203 9623 205
rect 9589 167 9623 169
rect 9589 95 9623 101
rect 9589 23 9623 33
rect 872 -49 993 -35
rect 906 -69 993 -49
rect 1027 -69 1061 -35
rect 1095 -69 1129 -35
rect 1163 -69 1197 -35
rect 1231 -69 1265 -35
rect 1299 -69 1333 -35
rect 1367 -69 1401 -35
rect 1435 -69 1469 -35
rect 1503 -69 1537 -35
rect 1571 -69 1605 -35
rect 1639 -69 1673 -35
rect 1707 -69 1741 -35
rect 1775 -69 1809 -35
rect 1843 -69 1877 -35
rect 1911 -69 1945 -35
rect 1979 -69 2013 -35
rect 2047 -69 2081 -35
rect 2115 -69 2149 -35
rect 2183 -69 2217 -35
rect 2251 -69 2285 -35
rect 2319 -69 2353 -35
rect 2387 -69 2421 -35
rect 2455 -69 2489 -35
rect 2523 -69 2557 -35
rect 2591 -69 2625 -35
rect 2659 -69 2693 -35
rect 2727 -69 2761 -35
rect 2795 -69 2829 -35
rect 2863 -69 2897 -35
rect 2931 -69 2965 -35
rect 2999 -69 3033 -35
rect 3067 -69 3101 -35
rect 3135 -69 3169 -35
rect 3203 -69 3237 -35
rect 3271 -69 3305 -35
rect 3339 -69 3373 -35
rect 3407 -69 3441 -35
rect 3475 -69 3509 -35
rect 3543 -69 3577 -35
rect 3611 -69 3645 -35
rect 3679 -69 3713 -35
rect 3747 -69 3781 -35
rect 3815 -69 3849 -35
rect 3883 -69 3917 -35
rect 3951 -69 3985 -35
rect 4019 -69 4053 -35
rect 4087 -69 4121 -35
rect 4155 -69 4189 -35
rect 4223 -69 4257 -35
rect 4291 -69 4325 -35
rect 4359 -69 4393 -35
rect 4427 -69 4461 -35
rect 4495 -69 4529 -35
rect 4563 -69 4597 -35
rect 4631 -69 4665 -35
rect 4699 -69 4733 -35
rect 4767 -69 4801 -35
rect 4835 -69 4869 -35
rect 4903 -69 4937 -35
rect 4971 -69 5005 -35
rect 5039 -69 5073 -35
rect 5107 -49 5388 -35
rect 5107 -69 5231 -49
rect 5265 -69 5388 -49
rect 5422 -69 5456 -35
rect 5490 -69 5524 -35
rect 5558 -69 5592 -35
rect 5626 -69 5660 -35
rect 5694 -69 5728 -35
rect 5762 -69 5796 -35
rect 5830 -69 5864 -35
rect 5898 -69 5932 -35
rect 5966 -69 6000 -35
rect 6034 -69 6068 -35
rect 6102 -69 6136 -35
rect 6170 -69 6204 -35
rect 6238 -69 6272 -35
rect 6306 -69 6340 -35
rect 6374 -69 6408 -35
rect 6442 -69 6476 -35
rect 6510 -69 6544 -35
rect 6578 -69 6612 -35
rect 6646 -69 6680 -35
rect 6714 -69 6748 -35
rect 6782 -69 6816 -35
rect 6850 -69 6884 -35
rect 6918 -69 6952 -35
rect 6986 -69 7020 -35
rect 7054 -69 7088 -35
rect 7122 -69 7156 -35
rect 7190 -69 7224 -35
rect 7258 -69 7292 -35
rect 7326 -69 7360 -35
rect 7394 -69 7428 -35
rect 7462 -69 7496 -35
rect 7530 -69 7564 -35
rect 7598 -69 7632 -35
rect 7666 -69 7700 -35
rect 7734 -69 7768 -35
rect 7802 -69 7836 -35
rect 7870 -69 7904 -35
rect 7938 -69 7972 -35
rect 8006 -69 8040 -35
rect 8074 -69 8108 -35
rect 8142 -69 8176 -35
rect 8210 -69 8244 -35
rect 8278 -69 8312 -35
rect 8346 -69 8380 -35
rect 8414 -69 8448 -35
rect 8482 -69 8516 -35
rect 8550 -69 8584 -35
rect 8618 -69 8652 -35
rect 8686 -69 8720 -35
rect 8754 -69 8788 -35
rect 8822 -69 8856 -35
rect 8890 -69 8924 -35
rect 8958 -69 8992 -35
rect 9026 -69 9060 -35
rect 9094 -69 9128 -35
rect 9162 -69 9196 -35
rect 9230 -69 9264 -35
rect 9298 -69 9332 -35
rect 9366 -69 9400 -35
rect 9434 -69 9468 -35
rect 9502 -49 9623 -35
rect 9502 -69 9589 -49
rect 872 -121 906 -103
rect 872 -193 906 -171
rect 872 -265 906 -239
rect 872 -337 906 -307
rect 872 -409 906 -375
rect 5230 -103 5231 -69
rect 5230 -121 5265 -103
rect 5230 -171 5231 -121
rect 5230 -193 5265 -171
rect 5230 -239 5231 -193
rect 5230 -265 5265 -239
rect 5230 -307 5231 -265
rect 5230 -337 5265 -307
rect 5230 -375 5231 -337
rect 872 -477 906 -443
rect 872 -545 906 -515
rect 987 -398 1021 -379
rect 987 -466 1021 -464
rect 987 -502 1021 -500
rect 987 -587 1021 -568
rect 1245 -398 1279 -379
rect 1245 -466 1279 -464
rect 1245 -502 1279 -500
rect 1245 -587 1279 -568
rect 1439 -398 1473 -379
rect 1439 -466 1473 -464
rect 1439 -502 1473 -500
rect 1439 -587 1473 -568
rect 1697 -398 1731 -379
rect 1697 -466 1731 -464
rect 1697 -502 1731 -500
rect 1697 -587 1731 -568
rect 1955 -398 1989 -379
rect 1955 -466 1989 -464
rect 1955 -502 1989 -500
rect 1955 -587 1989 -568
rect 2213 -398 2247 -379
rect 2213 -466 2247 -464
rect 2213 -502 2247 -500
rect 2213 -587 2247 -568
rect 2471 -398 2505 -379
rect 2471 -466 2505 -464
rect 2471 -502 2505 -500
rect 2471 -587 2505 -568
rect 2665 -398 2699 -379
rect 2665 -466 2699 -464
rect 2665 -502 2699 -500
rect 2665 -587 2699 -568
rect 2923 -398 2957 -379
rect 2923 -466 2957 -464
rect 2923 -502 2957 -500
rect 2923 -587 2957 -568
rect 3181 -398 3215 -379
rect 3181 -466 3215 -464
rect 3181 -502 3215 -500
rect 3181 -587 3215 -568
rect 3439 -398 3473 -379
rect 3439 -466 3473 -464
rect 3439 -502 3473 -500
rect 3439 -587 3473 -568
rect 3633 -398 3667 -379
rect 3633 -466 3667 -464
rect 3633 -502 3667 -500
rect 3633 -587 3667 -568
rect 3891 -398 3925 -379
rect 3891 -466 3925 -464
rect 3891 -502 3925 -500
rect 3891 -587 3925 -568
rect 4149 -398 4183 -379
rect 4149 -466 4183 -464
rect 4149 -502 4183 -500
rect 4149 -587 4183 -568
rect 4407 -398 4441 -379
rect 4407 -466 4441 -464
rect 4407 -502 4441 -500
rect 4407 -587 4441 -568
rect 4665 -398 4699 -379
rect 4665 -466 4699 -464
rect 4665 -502 4699 -500
rect 4665 -587 4699 -568
rect 4859 -398 4893 -379
rect 4859 -466 4893 -464
rect 4859 -502 4893 -500
rect 4859 -587 4893 -568
rect 5117 -398 5151 -379
rect 5117 -466 5151 -464
rect 5117 -502 5151 -500
rect 5117 -587 5151 -568
rect 5230 -409 5265 -375
rect 9589 -121 9623 -103
rect 9589 -193 9623 -171
rect 9589 -265 9623 -239
rect 9589 -337 9623 -307
rect 5230 -443 5231 -409
rect 5230 -477 5265 -443
rect 5230 -515 5231 -477
rect 5230 -545 5265 -515
rect 5230 -587 5231 -545
rect 5345 -398 5379 -379
rect 5345 -466 5379 -464
rect 5345 -502 5379 -500
rect 5345 -587 5379 -568
rect 5603 -398 5637 -379
rect 5603 -466 5637 -464
rect 5603 -502 5637 -500
rect 5603 -587 5637 -568
rect 5796 -398 5830 -379
rect 5796 -466 5830 -464
rect 5796 -502 5830 -500
rect 5796 -587 5830 -568
rect 6054 -398 6088 -379
rect 6054 -466 6088 -464
rect 6054 -502 6088 -500
rect 6054 -587 6088 -568
rect 6312 -398 6346 -379
rect 6312 -466 6346 -464
rect 6312 -502 6346 -500
rect 6312 -587 6346 -568
rect 6570 -398 6604 -379
rect 6570 -466 6604 -464
rect 6570 -502 6604 -500
rect 6570 -587 6604 -568
rect 6828 -398 6862 -379
rect 6828 -466 6862 -464
rect 6828 -502 6862 -500
rect 6828 -587 6862 -568
rect 7022 -398 7056 -379
rect 7022 -466 7056 -464
rect 7022 -502 7056 -500
rect 7022 -587 7056 -568
rect 7280 -398 7314 -379
rect 7280 -466 7314 -464
rect 7280 -502 7314 -500
rect 7280 -587 7314 -568
rect 7538 -398 7572 -379
rect 7538 -466 7572 -464
rect 7538 -502 7572 -500
rect 7538 -587 7572 -568
rect 7796 -398 7830 -379
rect 7796 -466 7830 -464
rect 7796 -502 7830 -500
rect 7796 -587 7830 -568
rect 7990 -398 8024 -379
rect 7990 -466 8024 -464
rect 7990 -502 8024 -500
rect 7990 -587 8024 -568
rect 8248 -398 8282 -379
rect 8248 -466 8282 -464
rect 8248 -502 8282 -500
rect 8248 -587 8282 -568
rect 8506 -398 8540 -379
rect 8506 -466 8540 -464
rect 8506 -502 8540 -500
rect 8506 -587 8540 -568
rect 8764 -398 8798 -379
rect 8764 -466 8798 -464
rect 8764 -502 8798 -500
rect 8764 -587 8798 -568
rect 9022 -398 9056 -379
rect 9022 -466 9056 -464
rect 9022 -502 9056 -500
rect 9022 -587 9056 -568
rect 9216 -398 9250 -379
rect 9216 -466 9250 -464
rect 9216 -502 9250 -500
rect 9216 -587 9250 -568
rect 9474 -398 9508 -379
rect 9474 -466 9508 -464
rect 9474 -502 9508 -500
rect 9474 -587 9508 -568
rect 9589 -409 9623 -375
rect 9589 -477 9623 -443
rect 9589 -545 9623 -515
rect 872 -613 906 -587
rect 5230 -613 5265 -587
rect 872 -681 906 -659
rect 1033 -664 1080 -630
rect 1116 -664 1150 -630
rect 1186 -664 1233 -630
rect 1485 -664 1532 -630
rect 1568 -664 1602 -630
rect 1638 -664 1685 -630
rect 1743 -664 1790 -630
rect 1826 -664 1860 -630
rect 1896 -664 1943 -630
rect 2001 -664 2048 -630
rect 2084 -664 2118 -630
rect 2154 -664 2201 -630
rect 2259 -664 2306 -630
rect 2342 -664 2376 -630
rect 2412 -664 2459 -630
rect 2711 -664 2758 -630
rect 2794 -664 2828 -630
rect 2864 -664 2911 -630
rect 2969 -664 3016 -630
rect 3052 -664 3086 -630
rect 3122 -664 3169 -630
rect 3227 -664 3274 -630
rect 3310 -664 3344 -630
rect 3380 -664 3427 -630
rect 3679 -664 3726 -630
rect 3762 -664 3796 -630
rect 3832 -664 3879 -630
rect 3937 -664 3984 -630
rect 4020 -664 4054 -630
rect 4090 -664 4137 -630
rect 4195 -664 4242 -630
rect 4278 -664 4312 -630
rect 4348 -664 4395 -630
rect 4453 -664 4500 -630
rect 4536 -664 4570 -630
rect 4606 -664 4653 -630
rect 4905 -664 4952 -630
rect 4988 -664 5022 -630
rect 5058 -664 5105 -630
rect 5230 -659 5231 -613
rect 9589 -613 9623 -587
rect 872 -749 906 -731
rect 872 -817 906 -803
rect 872 -885 906 -875
rect 872 -953 906 -947
rect 5230 -681 5265 -659
rect 5391 -664 5438 -630
rect 5474 -664 5508 -630
rect 5544 -664 5591 -630
rect 5842 -664 5889 -630
rect 5925 -664 5959 -630
rect 5995 -664 6042 -630
rect 6100 -664 6147 -630
rect 6183 -664 6217 -630
rect 6253 -664 6300 -630
rect 6358 -664 6405 -630
rect 6441 -664 6475 -630
rect 6511 -664 6558 -630
rect 6616 -664 6663 -630
rect 6699 -664 6733 -630
rect 6769 -664 6816 -630
rect 7068 -664 7115 -630
rect 7151 -664 7185 -630
rect 7221 -664 7268 -630
rect 7326 -664 7373 -630
rect 7409 -664 7443 -630
rect 7479 -664 7526 -630
rect 7584 -664 7631 -630
rect 7667 -664 7701 -630
rect 7737 -664 7784 -630
rect 8036 -664 8083 -630
rect 8119 -664 8153 -630
rect 8189 -664 8236 -630
rect 8294 -664 8341 -630
rect 8377 -664 8411 -630
rect 8447 -664 8494 -630
rect 8552 -664 8599 -630
rect 8635 -664 8669 -630
rect 8705 -664 8752 -630
rect 8810 -664 8857 -630
rect 8893 -664 8927 -630
rect 8963 -664 9010 -630
rect 9262 -664 9309 -630
rect 9345 -664 9379 -630
rect 9415 -664 9462 -630
rect 5230 -731 5231 -681
rect 5230 -749 5265 -731
rect 5230 -803 5231 -749
rect 5230 -817 5265 -803
rect 5230 -875 5231 -817
rect 5230 -885 5265 -875
rect 5230 -947 5231 -885
rect 5230 -953 5265 -947
rect 872 -1021 906 -1019
rect 1033 -1027 1080 -993
rect 1116 -1027 1150 -993
rect 1186 -1027 1233 -993
rect 1485 -1027 1532 -993
rect 1568 -1027 1602 -993
rect 1638 -1027 1685 -993
rect 1743 -1027 1790 -993
rect 1826 -1027 1860 -993
rect 1896 -1027 1943 -993
rect 2001 -1027 2048 -993
rect 2084 -1027 2118 -993
rect 2154 -1027 2201 -993
rect 2259 -1027 2306 -993
rect 2342 -1027 2376 -993
rect 2412 -1027 2459 -993
rect 2711 -1027 2758 -993
rect 2794 -1027 2828 -993
rect 2864 -1027 2911 -993
rect 2969 -1027 3016 -993
rect 3052 -1027 3086 -993
rect 3122 -1027 3169 -993
rect 3227 -1027 3274 -993
rect 3310 -1027 3344 -993
rect 3380 -1027 3427 -993
rect 3679 -1027 3726 -993
rect 3762 -1027 3796 -993
rect 3832 -1027 3879 -993
rect 3937 -1027 3984 -993
rect 4020 -1027 4054 -993
rect 4090 -1027 4137 -993
rect 4195 -1027 4242 -993
rect 4278 -1027 4312 -993
rect 4348 -1027 4395 -993
rect 4453 -1027 4500 -993
rect 4536 -1027 4570 -993
rect 4606 -1027 4653 -993
rect 4905 -1027 4952 -993
rect 4988 -1027 5022 -993
rect 5058 -1027 5105 -993
rect 5230 -1019 5231 -953
rect 9589 -681 9623 -659
rect 9589 -749 9623 -731
rect 9589 -817 9623 -803
rect 9589 -885 9623 -875
rect 9589 -953 9623 -947
rect 5230 -1021 5265 -1019
rect 872 -1057 906 -1055
rect 5230 -1055 5231 -1021
rect 5391 -1027 5438 -993
rect 5474 -1027 5508 -993
rect 5544 -1027 5591 -993
rect 5842 -1027 5889 -993
rect 5925 -1027 5959 -993
rect 5995 -1027 6042 -993
rect 6100 -1027 6147 -993
rect 6183 -1027 6217 -993
rect 6253 -1027 6300 -993
rect 6358 -1027 6405 -993
rect 6441 -1027 6475 -993
rect 6511 -1027 6558 -993
rect 6616 -1027 6663 -993
rect 6699 -1027 6733 -993
rect 6769 -1027 6816 -993
rect 7068 -1027 7115 -993
rect 7151 -1027 7185 -993
rect 7221 -1027 7268 -993
rect 7326 -1027 7373 -993
rect 7409 -1027 7443 -993
rect 7479 -1027 7526 -993
rect 7584 -1027 7631 -993
rect 7667 -1027 7701 -993
rect 7737 -1027 7784 -993
rect 8036 -1027 8083 -993
rect 8119 -1027 8153 -993
rect 8189 -1027 8236 -993
rect 8294 -1027 8341 -993
rect 8377 -1027 8411 -993
rect 8447 -1027 8494 -993
rect 8552 -1027 8599 -993
rect 8635 -1027 8669 -993
rect 8705 -1027 8752 -993
rect 8810 -1027 8857 -993
rect 8893 -1027 8927 -993
rect 8963 -1027 9010 -993
rect 9262 -1027 9309 -993
rect 9345 -1027 9379 -993
rect 9415 -1027 9462 -993
rect 9589 -1021 9623 -1019
rect 5230 -1057 5265 -1055
rect 872 -1129 906 -1123
rect 872 -1201 906 -1191
rect 872 -1273 906 -1259
rect 987 -1089 1021 -1070
rect 987 -1157 1021 -1155
rect 987 -1193 1021 -1191
rect 987 -1278 1021 -1259
rect 1245 -1089 1279 -1070
rect 1245 -1157 1279 -1155
rect 1245 -1193 1279 -1191
rect 1245 -1278 1279 -1259
rect 1439 -1089 1473 -1070
rect 1439 -1157 1473 -1155
rect 1439 -1193 1473 -1191
rect 1439 -1278 1473 -1259
rect 1697 -1089 1731 -1070
rect 1697 -1157 1731 -1155
rect 1697 -1193 1731 -1191
rect 1697 -1278 1731 -1259
rect 1955 -1089 1989 -1070
rect 1955 -1157 1989 -1155
rect 1955 -1193 1989 -1191
rect 1955 -1278 1989 -1259
rect 2213 -1089 2247 -1070
rect 2213 -1157 2247 -1155
rect 2213 -1193 2247 -1191
rect 2213 -1278 2247 -1259
rect 2471 -1089 2505 -1070
rect 2471 -1157 2505 -1155
rect 2471 -1193 2505 -1191
rect 2471 -1278 2505 -1259
rect 2665 -1089 2699 -1070
rect 2665 -1157 2699 -1155
rect 2665 -1193 2699 -1191
rect 2665 -1278 2699 -1259
rect 2923 -1089 2957 -1070
rect 2923 -1157 2957 -1155
rect 2923 -1193 2957 -1191
rect 2923 -1278 2957 -1259
rect 3181 -1089 3215 -1070
rect 3181 -1157 3215 -1155
rect 3181 -1193 3215 -1191
rect 3181 -1278 3215 -1259
rect 3439 -1089 3473 -1070
rect 3439 -1157 3473 -1155
rect 3439 -1193 3473 -1191
rect 3439 -1278 3473 -1259
rect 3633 -1089 3667 -1070
rect 3633 -1157 3667 -1155
rect 3633 -1193 3667 -1191
rect 3633 -1278 3667 -1259
rect 3891 -1089 3925 -1070
rect 3891 -1157 3925 -1155
rect 3891 -1193 3925 -1191
rect 3891 -1278 3925 -1259
rect 4149 -1089 4183 -1070
rect 4149 -1157 4183 -1155
rect 4149 -1193 4183 -1191
rect 4149 -1278 4183 -1259
rect 4407 -1089 4441 -1070
rect 4407 -1157 4441 -1155
rect 4407 -1193 4441 -1191
rect 4407 -1278 4441 -1259
rect 4665 -1089 4699 -1070
rect 4665 -1157 4699 -1155
rect 4665 -1193 4699 -1191
rect 4665 -1278 4699 -1259
rect 4859 -1089 4893 -1070
rect 4859 -1157 4893 -1155
rect 4859 -1193 4893 -1191
rect 4859 -1278 4893 -1259
rect 5117 -1089 5151 -1070
rect 5117 -1157 5151 -1155
rect 5117 -1193 5151 -1191
rect 5117 -1278 5151 -1259
rect 5230 -1123 5231 -1057
rect 9589 -1057 9623 -1055
rect 5230 -1129 5265 -1123
rect 5230 -1191 5231 -1129
rect 5230 -1201 5265 -1191
rect 5230 -1259 5231 -1201
rect 5230 -1273 5265 -1259
rect 872 -1345 906 -1327
rect 872 -1417 906 -1395
rect 872 -1489 906 -1463
rect 872 -1561 906 -1531
rect 872 -1633 906 -1595
rect 5230 -1327 5231 -1273
rect 5345 -1089 5379 -1070
rect 5345 -1157 5379 -1155
rect 5345 -1193 5379 -1191
rect 5345 -1278 5379 -1259
rect 5603 -1089 5637 -1070
rect 5603 -1157 5637 -1155
rect 5603 -1193 5637 -1191
rect 5603 -1278 5637 -1259
rect 5796 -1089 5830 -1070
rect 5796 -1157 5830 -1155
rect 5796 -1193 5830 -1191
rect 5796 -1278 5830 -1259
rect 6054 -1089 6088 -1070
rect 6054 -1157 6088 -1155
rect 6054 -1193 6088 -1191
rect 6054 -1278 6088 -1259
rect 6312 -1089 6346 -1070
rect 6312 -1157 6346 -1155
rect 6312 -1193 6346 -1191
rect 6312 -1278 6346 -1259
rect 6570 -1089 6604 -1070
rect 6570 -1157 6604 -1155
rect 6570 -1193 6604 -1191
rect 6570 -1278 6604 -1259
rect 6828 -1089 6862 -1070
rect 6828 -1157 6862 -1155
rect 6828 -1193 6862 -1191
rect 6828 -1278 6862 -1259
rect 7022 -1089 7056 -1070
rect 7022 -1157 7056 -1155
rect 7022 -1193 7056 -1191
rect 7022 -1278 7056 -1259
rect 7280 -1089 7314 -1070
rect 7280 -1157 7314 -1155
rect 7280 -1193 7314 -1191
rect 7280 -1278 7314 -1259
rect 7538 -1089 7572 -1070
rect 7538 -1157 7572 -1155
rect 7538 -1193 7572 -1191
rect 7538 -1278 7572 -1259
rect 7796 -1089 7830 -1070
rect 7796 -1157 7830 -1155
rect 7796 -1193 7830 -1191
rect 7796 -1278 7830 -1259
rect 7990 -1089 8024 -1070
rect 7990 -1157 8024 -1155
rect 7990 -1193 8024 -1191
rect 7990 -1278 8024 -1259
rect 8248 -1089 8282 -1070
rect 8248 -1157 8282 -1155
rect 8248 -1193 8282 -1191
rect 8248 -1278 8282 -1259
rect 8506 -1089 8540 -1070
rect 8506 -1157 8540 -1155
rect 8506 -1193 8540 -1191
rect 8506 -1278 8540 -1259
rect 8764 -1089 8798 -1070
rect 8764 -1157 8798 -1155
rect 8764 -1193 8798 -1191
rect 8764 -1278 8798 -1259
rect 9022 -1089 9056 -1070
rect 9022 -1157 9056 -1155
rect 9022 -1193 9056 -1191
rect 9022 -1278 9056 -1259
rect 9216 -1089 9250 -1070
rect 9216 -1157 9250 -1155
rect 9216 -1193 9250 -1191
rect 9216 -1278 9250 -1259
rect 9474 -1089 9508 -1070
rect 9474 -1157 9508 -1155
rect 9474 -1193 9508 -1191
rect 9474 -1278 9508 -1259
rect 9589 -1129 9623 -1123
rect 9589 -1201 9623 -1191
rect 9589 -1273 9623 -1259
rect 5230 -1345 5265 -1327
rect 5230 -1395 5231 -1345
rect 5230 -1417 5265 -1395
rect 5230 -1463 5231 -1417
rect 5230 -1489 5265 -1463
rect 5230 -1531 5231 -1489
rect 5230 -1561 5265 -1531
rect 5230 -1595 5231 -1561
rect 5230 -1633 5265 -1595
rect 9589 -1345 9623 -1327
rect 9589 -1417 9623 -1395
rect 9589 -1489 9623 -1463
rect 9589 -1561 9623 -1531
rect 9589 -1633 9623 -1595
rect 906 -1667 993 -1633
rect 1027 -1667 1061 -1633
rect 1095 -1667 1129 -1633
rect 1163 -1667 1197 -1633
rect 1231 -1667 1265 -1633
rect 1299 -1667 1333 -1633
rect 1367 -1667 1401 -1633
rect 1435 -1667 1469 -1633
rect 1503 -1667 1537 -1633
rect 1571 -1667 1605 -1633
rect 1639 -1667 1673 -1633
rect 1707 -1667 1741 -1633
rect 1775 -1667 1809 -1633
rect 1843 -1667 1877 -1633
rect 1911 -1667 1945 -1633
rect 1979 -1667 2013 -1633
rect 2047 -1667 2081 -1633
rect 2115 -1667 2149 -1633
rect 2183 -1667 2217 -1633
rect 2251 -1667 2285 -1633
rect 2319 -1667 2353 -1633
rect 2387 -1667 2421 -1633
rect 2455 -1667 2489 -1633
rect 2523 -1667 2557 -1633
rect 2591 -1667 2625 -1633
rect 2659 -1667 2693 -1633
rect 2727 -1667 2761 -1633
rect 2795 -1667 2829 -1633
rect 2863 -1667 2897 -1633
rect 2931 -1667 2965 -1633
rect 2999 -1667 3033 -1633
rect 3067 -1667 3101 -1633
rect 3135 -1667 3169 -1633
rect 3203 -1667 3237 -1633
rect 3271 -1667 3305 -1633
rect 3339 -1667 3373 -1633
rect 3407 -1667 3441 -1633
rect 3475 -1667 3509 -1633
rect 3543 -1667 3577 -1633
rect 3611 -1667 3645 -1633
rect 3679 -1667 3713 -1633
rect 3747 -1667 3781 -1633
rect 3815 -1667 3849 -1633
rect 3883 -1667 3917 -1633
rect 3951 -1667 3985 -1633
rect 4019 -1667 4053 -1633
rect 4087 -1667 4121 -1633
rect 4155 -1667 4189 -1633
rect 4223 -1667 4257 -1633
rect 4291 -1667 4325 -1633
rect 4359 -1667 4393 -1633
rect 4427 -1667 4461 -1633
rect 4495 -1667 4529 -1633
rect 4563 -1667 4597 -1633
rect 4631 -1667 4665 -1633
rect 4699 -1667 4733 -1633
rect 4767 -1667 4801 -1633
rect 4835 -1667 4869 -1633
rect 4903 -1667 4937 -1633
rect 4971 -1667 5005 -1633
rect 5039 -1667 5073 -1633
rect 5107 -1667 5231 -1633
rect 5265 -1667 5388 -1633
rect 5422 -1667 5456 -1633
rect 5490 -1667 5524 -1633
rect 5558 -1667 5592 -1633
rect 5626 -1667 5660 -1633
rect 5694 -1667 5728 -1633
rect 5762 -1667 5796 -1633
rect 5830 -1667 5864 -1633
rect 5898 -1667 5932 -1633
rect 5966 -1667 6000 -1633
rect 6034 -1667 6068 -1633
rect 6102 -1667 6136 -1633
rect 6170 -1667 6204 -1633
rect 6238 -1667 6272 -1633
rect 6306 -1667 6340 -1633
rect 6374 -1667 6408 -1633
rect 6442 -1667 6476 -1633
rect 6510 -1667 6544 -1633
rect 6578 -1667 6612 -1633
rect 6646 -1667 6680 -1633
rect 6714 -1667 6748 -1633
rect 6782 -1667 6816 -1633
rect 6850 -1667 6884 -1633
rect 6918 -1667 6952 -1633
rect 6986 -1667 7020 -1633
rect 7054 -1667 7088 -1633
rect 7122 -1667 7156 -1633
rect 7190 -1667 7224 -1633
rect 7258 -1667 7292 -1633
rect 7326 -1667 7360 -1633
rect 7394 -1667 7428 -1633
rect 7462 -1667 7496 -1633
rect 7530 -1667 7564 -1633
rect 7598 -1667 7632 -1633
rect 7666 -1667 7700 -1633
rect 7734 -1667 7768 -1633
rect 7802 -1667 7836 -1633
rect 7870 -1667 7904 -1633
rect 7938 -1667 7972 -1633
rect 8006 -1667 8040 -1633
rect 8074 -1667 8108 -1633
rect 8142 -1667 8176 -1633
rect 8210 -1667 8244 -1633
rect 8278 -1667 8312 -1633
rect 8346 -1667 8380 -1633
rect 8414 -1667 8448 -1633
rect 8482 -1667 8516 -1633
rect 8550 -1667 8584 -1633
rect 8618 -1667 8652 -1633
rect 8686 -1667 8720 -1633
rect 8754 -1667 8788 -1633
rect 8822 -1667 8856 -1633
rect 8890 -1667 8924 -1633
rect 8958 -1667 8992 -1633
rect 9026 -1667 9060 -1633
rect 9094 -1667 9128 -1633
rect 9162 -1667 9196 -1633
rect 9230 -1667 9264 -1633
rect 9298 -1667 9332 -1633
rect 9366 -1667 9400 -1633
rect 9434 -1667 9468 -1633
rect 9502 -1667 9589 -1633
rect 872 -1705 906 -1667
rect 872 -1769 906 -1739
rect 872 -1837 906 -1811
rect 872 -1905 906 -1883
rect 872 -1973 906 -1955
rect 5230 -1705 5265 -1667
rect 5230 -1739 5231 -1705
rect 5230 -1769 5265 -1739
rect 5230 -1811 5231 -1769
rect 5230 -1837 5265 -1811
rect 5230 -1883 5231 -1837
rect 5230 -1905 5265 -1883
rect 5230 -1955 5231 -1905
rect 5230 -1973 5265 -1955
rect 872 -2041 906 -2027
rect 872 -2109 906 -2099
rect 872 -2177 906 -2171
rect 987 -2045 1021 -2026
rect 987 -2113 1021 -2111
rect 987 -2149 1021 -2147
rect 987 -2234 1021 -2215
rect 1245 -2045 1279 -2026
rect 1245 -2113 1279 -2111
rect 1245 -2149 1279 -2147
rect 1245 -2234 1279 -2215
rect 1439 -2045 1473 -2026
rect 1439 -2113 1473 -2111
rect 1439 -2149 1473 -2147
rect 1439 -2234 1473 -2215
rect 1697 -2045 1731 -2026
rect 1697 -2113 1731 -2111
rect 1697 -2149 1731 -2147
rect 1697 -2234 1731 -2215
rect 1955 -2045 1989 -2026
rect 1955 -2113 1989 -2111
rect 1955 -2149 1989 -2147
rect 1955 -2234 1989 -2215
rect 2213 -2045 2247 -2026
rect 2213 -2113 2247 -2111
rect 2213 -2149 2247 -2147
rect 2213 -2234 2247 -2215
rect 2471 -2045 2505 -2026
rect 2471 -2113 2505 -2111
rect 2471 -2149 2505 -2147
rect 2471 -2234 2505 -2215
rect 2665 -2045 2699 -2026
rect 2665 -2113 2699 -2111
rect 2665 -2149 2699 -2147
rect 2665 -2234 2699 -2215
rect 2923 -2045 2957 -2026
rect 2923 -2113 2957 -2111
rect 2923 -2149 2957 -2147
rect 2923 -2234 2957 -2215
rect 3181 -2045 3215 -2026
rect 3181 -2113 3215 -2111
rect 3181 -2149 3215 -2147
rect 3181 -2234 3215 -2215
rect 3439 -2045 3473 -2026
rect 3439 -2113 3473 -2111
rect 3439 -2149 3473 -2147
rect 3439 -2234 3473 -2215
rect 3633 -2045 3667 -2026
rect 3633 -2113 3667 -2111
rect 3633 -2149 3667 -2147
rect 3633 -2234 3667 -2215
rect 3891 -2045 3925 -2026
rect 3891 -2113 3925 -2111
rect 3891 -2149 3925 -2147
rect 3891 -2234 3925 -2215
rect 4149 -2045 4183 -2026
rect 4149 -2113 4183 -2111
rect 4149 -2149 4183 -2147
rect 4149 -2234 4183 -2215
rect 4407 -2045 4441 -2026
rect 4407 -2113 4441 -2111
rect 4407 -2149 4441 -2147
rect 4407 -2234 4441 -2215
rect 4665 -2045 4699 -2026
rect 4665 -2113 4699 -2111
rect 4665 -2149 4699 -2147
rect 4665 -2234 4699 -2215
rect 4859 -2045 4893 -2026
rect 4859 -2113 4893 -2111
rect 4859 -2149 4893 -2147
rect 4859 -2234 4893 -2215
rect 5117 -2045 5151 -2026
rect 5117 -2113 5151 -2111
rect 5117 -2149 5151 -2147
rect 5117 -2234 5151 -2215
rect 5230 -2027 5231 -1973
rect 9589 -1705 9623 -1667
rect 9589 -1769 9623 -1739
rect 9589 -1837 9623 -1811
rect 9589 -1905 9623 -1883
rect 9589 -1973 9623 -1955
rect 5230 -2041 5265 -2027
rect 5230 -2099 5231 -2041
rect 5230 -2109 5265 -2099
rect 5230 -2171 5231 -2109
rect 5230 -2177 5265 -2171
rect 872 -2245 906 -2243
rect 5230 -2243 5231 -2177
rect 5345 -2045 5379 -2026
rect 5345 -2113 5379 -2111
rect 5345 -2149 5379 -2147
rect 5345 -2234 5379 -2215
rect 5603 -2045 5637 -2026
rect 5603 -2113 5637 -2111
rect 5603 -2149 5637 -2147
rect 5603 -2234 5637 -2215
rect 5796 -2045 5830 -2026
rect 5796 -2113 5830 -2111
rect 5796 -2149 5830 -2147
rect 5796 -2234 5830 -2215
rect 6054 -2045 6088 -2026
rect 6054 -2113 6088 -2111
rect 6054 -2149 6088 -2147
rect 6054 -2234 6088 -2215
rect 6312 -2045 6346 -2026
rect 6312 -2113 6346 -2111
rect 6312 -2149 6346 -2147
rect 6312 -2234 6346 -2215
rect 6570 -2045 6604 -2026
rect 6570 -2113 6604 -2111
rect 6570 -2149 6604 -2147
rect 6570 -2234 6604 -2215
rect 6828 -2045 6862 -2026
rect 6828 -2113 6862 -2111
rect 6828 -2149 6862 -2147
rect 6828 -2234 6862 -2215
rect 7022 -2045 7056 -2026
rect 7022 -2113 7056 -2111
rect 7022 -2149 7056 -2147
rect 7022 -2234 7056 -2215
rect 7280 -2045 7314 -2026
rect 7280 -2113 7314 -2111
rect 7280 -2149 7314 -2147
rect 7280 -2234 7314 -2215
rect 7538 -2045 7572 -2026
rect 7538 -2113 7572 -2111
rect 7538 -2149 7572 -2147
rect 7538 -2234 7572 -2215
rect 7796 -2045 7830 -2026
rect 7796 -2113 7830 -2111
rect 7796 -2149 7830 -2147
rect 7796 -2234 7830 -2215
rect 7990 -2045 8024 -2026
rect 7990 -2113 8024 -2111
rect 7990 -2149 8024 -2147
rect 7990 -2234 8024 -2215
rect 8248 -2045 8282 -2026
rect 8248 -2113 8282 -2111
rect 8248 -2149 8282 -2147
rect 8248 -2234 8282 -2215
rect 8506 -2045 8540 -2026
rect 8506 -2113 8540 -2111
rect 8506 -2149 8540 -2147
rect 8506 -2234 8540 -2215
rect 8764 -2045 8798 -2026
rect 8764 -2113 8798 -2111
rect 8764 -2149 8798 -2147
rect 8764 -2234 8798 -2215
rect 9022 -2045 9056 -2026
rect 9022 -2113 9056 -2111
rect 9022 -2149 9056 -2147
rect 9022 -2234 9056 -2215
rect 9216 -2045 9250 -2026
rect 9216 -2113 9250 -2111
rect 9216 -2149 9250 -2147
rect 9216 -2234 9250 -2215
rect 9474 -2045 9508 -2026
rect 9474 -2113 9508 -2111
rect 9474 -2149 9508 -2147
rect 9474 -2234 9508 -2215
rect 9589 -2041 9623 -2027
rect 9589 -2109 9623 -2099
rect 9589 -2177 9623 -2171
rect 5230 -2245 5265 -2243
rect 872 -2281 906 -2279
rect 1033 -2311 1080 -2277
rect 1116 -2311 1150 -2277
rect 1186 -2311 1233 -2277
rect 1485 -2311 1532 -2277
rect 1568 -2311 1602 -2277
rect 1638 -2311 1685 -2277
rect 1743 -2311 1790 -2277
rect 1826 -2311 1860 -2277
rect 1896 -2311 1943 -2277
rect 2001 -2311 2048 -2277
rect 2084 -2311 2118 -2277
rect 2154 -2311 2201 -2277
rect 2259 -2311 2306 -2277
rect 2342 -2311 2376 -2277
rect 2412 -2311 2459 -2277
rect 2711 -2311 2758 -2277
rect 2794 -2311 2828 -2277
rect 2864 -2311 2911 -2277
rect 2969 -2311 3016 -2277
rect 3052 -2311 3086 -2277
rect 3122 -2311 3169 -2277
rect 3227 -2311 3274 -2277
rect 3310 -2311 3344 -2277
rect 3380 -2311 3427 -2277
rect 3679 -2311 3726 -2277
rect 3762 -2311 3796 -2277
rect 3832 -2311 3879 -2277
rect 3937 -2311 3984 -2277
rect 4020 -2311 4054 -2277
rect 4090 -2311 4137 -2277
rect 4195 -2311 4242 -2277
rect 4278 -2311 4312 -2277
rect 4348 -2311 4395 -2277
rect 4453 -2311 4500 -2277
rect 4536 -2311 4570 -2277
rect 4606 -2311 4653 -2277
rect 4905 -2311 4952 -2277
rect 4988 -2311 5022 -2277
rect 5058 -2311 5105 -2277
rect 5230 -2279 5231 -2245
rect 9589 -2245 9623 -2243
rect 5230 -2281 5265 -2279
rect 872 -2353 906 -2347
rect 872 -2425 906 -2415
rect 872 -2497 906 -2483
rect 872 -2569 906 -2551
rect 872 -2641 906 -2619
rect 5230 -2347 5231 -2281
rect 5391 -2311 5438 -2277
rect 5474 -2311 5508 -2277
rect 5544 -2311 5591 -2277
rect 5842 -2311 5889 -2277
rect 5925 -2311 5959 -2277
rect 5995 -2311 6042 -2277
rect 6100 -2311 6147 -2277
rect 6183 -2311 6217 -2277
rect 6253 -2311 6300 -2277
rect 6358 -2311 6405 -2277
rect 6441 -2311 6475 -2277
rect 6511 -2311 6558 -2277
rect 6616 -2311 6663 -2277
rect 6699 -2311 6733 -2277
rect 6769 -2311 6816 -2277
rect 7068 -2311 7115 -2277
rect 7151 -2311 7185 -2277
rect 7221 -2311 7268 -2277
rect 7326 -2311 7373 -2277
rect 7409 -2311 7443 -2277
rect 7479 -2311 7526 -2277
rect 7584 -2311 7631 -2277
rect 7667 -2311 7701 -2277
rect 7737 -2311 7784 -2277
rect 8036 -2311 8083 -2277
rect 8119 -2311 8153 -2277
rect 8189 -2311 8236 -2277
rect 8294 -2311 8341 -2277
rect 8377 -2311 8411 -2277
rect 8447 -2311 8494 -2277
rect 8552 -2311 8599 -2277
rect 8635 -2311 8669 -2277
rect 8705 -2311 8752 -2277
rect 8810 -2311 8857 -2277
rect 8893 -2311 8927 -2277
rect 8963 -2311 9010 -2277
rect 9262 -2311 9309 -2277
rect 9345 -2311 9379 -2277
rect 9415 -2311 9462 -2277
rect 9589 -2281 9623 -2279
rect 5230 -2353 5265 -2347
rect 5230 -2415 5231 -2353
rect 5230 -2425 5265 -2415
rect 5230 -2483 5231 -2425
rect 5230 -2497 5265 -2483
rect 5230 -2551 5231 -2497
rect 5230 -2569 5265 -2551
rect 5230 -2619 5231 -2569
rect 1033 -2674 1080 -2640
rect 1116 -2674 1150 -2640
rect 1186 -2674 1233 -2640
rect 1485 -2674 1532 -2640
rect 1568 -2674 1602 -2640
rect 1638 -2674 1685 -2640
rect 1743 -2674 1790 -2640
rect 1826 -2674 1860 -2640
rect 1896 -2674 1943 -2640
rect 2001 -2674 2048 -2640
rect 2084 -2674 2118 -2640
rect 2154 -2674 2201 -2640
rect 2259 -2674 2306 -2640
rect 2342 -2674 2376 -2640
rect 2412 -2674 2459 -2640
rect 2711 -2674 2758 -2640
rect 2794 -2674 2828 -2640
rect 2864 -2674 2911 -2640
rect 2969 -2674 3016 -2640
rect 3052 -2674 3086 -2640
rect 3122 -2674 3169 -2640
rect 3227 -2674 3274 -2640
rect 3310 -2674 3344 -2640
rect 3380 -2674 3427 -2640
rect 3679 -2674 3726 -2640
rect 3762 -2674 3796 -2640
rect 3832 -2674 3879 -2640
rect 3937 -2674 3984 -2640
rect 4020 -2674 4054 -2640
rect 4090 -2674 4137 -2640
rect 4195 -2674 4242 -2640
rect 4278 -2674 4312 -2640
rect 4348 -2674 4395 -2640
rect 4453 -2674 4500 -2640
rect 4536 -2674 4570 -2640
rect 4606 -2674 4653 -2640
rect 4905 -2674 4952 -2640
rect 4988 -2674 5022 -2640
rect 5058 -2674 5105 -2640
rect 5230 -2641 5265 -2619
rect 9589 -2353 9623 -2347
rect 9589 -2425 9623 -2415
rect 9589 -2497 9623 -2483
rect 9589 -2569 9623 -2551
rect 872 -2713 906 -2687
rect 5230 -2687 5231 -2641
rect 5391 -2674 5438 -2640
rect 5474 -2674 5508 -2640
rect 5544 -2674 5591 -2640
rect 5842 -2674 5889 -2640
rect 5925 -2674 5959 -2640
rect 5995 -2674 6042 -2640
rect 6100 -2674 6147 -2640
rect 6183 -2674 6217 -2640
rect 6253 -2674 6300 -2640
rect 6358 -2674 6405 -2640
rect 6441 -2674 6475 -2640
rect 6511 -2674 6558 -2640
rect 6616 -2674 6663 -2640
rect 6699 -2674 6733 -2640
rect 6769 -2674 6816 -2640
rect 7068 -2674 7115 -2640
rect 7151 -2674 7185 -2640
rect 7221 -2674 7268 -2640
rect 7326 -2674 7373 -2640
rect 7409 -2674 7443 -2640
rect 7479 -2674 7526 -2640
rect 7584 -2674 7631 -2640
rect 7667 -2674 7701 -2640
rect 7737 -2674 7784 -2640
rect 8036 -2674 8083 -2640
rect 8119 -2674 8153 -2640
rect 8189 -2674 8236 -2640
rect 8294 -2674 8341 -2640
rect 8377 -2674 8411 -2640
rect 8447 -2674 8494 -2640
rect 8552 -2674 8599 -2640
rect 8635 -2674 8669 -2640
rect 8705 -2674 8752 -2640
rect 8810 -2674 8857 -2640
rect 8893 -2674 8927 -2640
rect 8963 -2674 9010 -2640
rect 9262 -2674 9309 -2640
rect 9345 -2674 9379 -2640
rect 9415 -2674 9462 -2640
rect 9589 -2641 9623 -2619
rect 5230 -2713 5265 -2687
rect 872 -2785 906 -2755
rect 872 -2857 906 -2823
rect 872 -2925 906 -2891
rect 987 -2736 1021 -2717
rect 987 -2804 1021 -2802
rect 987 -2840 1021 -2838
rect 987 -2925 1021 -2906
rect 1245 -2736 1279 -2717
rect 1245 -2804 1279 -2802
rect 1245 -2840 1279 -2838
rect 1245 -2925 1279 -2906
rect 1439 -2736 1473 -2717
rect 1439 -2804 1473 -2802
rect 1439 -2840 1473 -2838
rect 1439 -2925 1473 -2906
rect 1697 -2736 1731 -2717
rect 1697 -2804 1731 -2802
rect 1697 -2840 1731 -2838
rect 1697 -2925 1731 -2906
rect 1955 -2736 1989 -2717
rect 1955 -2804 1989 -2802
rect 1955 -2840 1989 -2838
rect 1955 -2925 1989 -2906
rect 2213 -2736 2247 -2717
rect 2213 -2804 2247 -2802
rect 2213 -2840 2247 -2838
rect 2213 -2925 2247 -2906
rect 2471 -2736 2505 -2717
rect 2471 -2804 2505 -2802
rect 2471 -2840 2505 -2838
rect 2471 -2925 2505 -2906
rect 2665 -2736 2699 -2717
rect 2665 -2804 2699 -2802
rect 2665 -2840 2699 -2838
rect 2665 -2925 2699 -2906
rect 2923 -2736 2957 -2717
rect 2923 -2804 2957 -2802
rect 2923 -2840 2957 -2838
rect 2923 -2925 2957 -2906
rect 3181 -2736 3215 -2717
rect 3181 -2804 3215 -2802
rect 3181 -2840 3215 -2838
rect 3181 -2925 3215 -2906
rect 3439 -2736 3473 -2717
rect 3439 -2804 3473 -2802
rect 3439 -2840 3473 -2838
rect 3439 -2925 3473 -2906
rect 3633 -2736 3667 -2717
rect 3633 -2804 3667 -2802
rect 3633 -2840 3667 -2838
rect 3633 -2925 3667 -2906
rect 3891 -2736 3925 -2717
rect 3891 -2804 3925 -2802
rect 3891 -2840 3925 -2838
rect 3891 -2925 3925 -2906
rect 4149 -2736 4183 -2717
rect 4149 -2804 4183 -2802
rect 4149 -2840 4183 -2838
rect 4149 -2925 4183 -2906
rect 4407 -2736 4441 -2717
rect 4407 -2804 4441 -2802
rect 4407 -2840 4441 -2838
rect 4407 -2925 4441 -2906
rect 4665 -2736 4699 -2717
rect 4665 -2804 4699 -2802
rect 4665 -2840 4699 -2838
rect 4665 -2925 4699 -2906
rect 4859 -2736 4893 -2717
rect 4859 -2804 4893 -2802
rect 4859 -2840 4893 -2838
rect 4859 -2925 4893 -2906
rect 5117 -2736 5151 -2717
rect 5117 -2804 5151 -2802
rect 5117 -2840 5151 -2838
rect 5117 -2925 5151 -2906
rect 5230 -2755 5231 -2713
rect 9589 -2713 9623 -2687
rect 5230 -2785 5265 -2755
rect 5230 -2823 5231 -2785
rect 5230 -2857 5265 -2823
rect 5230 -2891 5231 -2857
rect 5230 -2925 5265 -2891
rect 5345 -2736 5379 -2717
rect 5345 -2804 5379 -2802
rect 5345 -2840 5379 -2838
rect 5345 -2925 5379 -2906
rect 5603 -2736 5637 -2717
rect 5603 -2804 5637 -2802
rect 5603 -2840 5637 -2838
rect 5603 -2925 5637 -2906
rect 5796 -2736 5830 -2717
rect 5796 -2804 5830 -2802
rect 5796 -2840 5830 -2838
rect 5796 -2925 5830 -2906
rect 6054 -2736 6088 -2717
rect 6054 -2804 6088 -2802
rect 6054 -2840 6088 -2838
rect 6054 -2925 6088 -2906
rect 6312 -2736 6346 -2717
rect 6312 -2804 6346 -2802
rect 6312 -2840 6346 -2838
rect 6312 -2925 6346 -2906
rect 6570 -2736 6604 -2717
rect 6570 -2804 6604 -2802
rect 6570 -2840 6604 -2838
rect 6570 -2925 6604 -2906
rect 6828 -2736 6862 -2717
rect 6828 -2804 6862 -2802
rect 6828 -2840 6862 -2838
rect 6828 -2925 6862 -2906
rect 7022 -2736 7056 -2717
rect 7022 -2804 7056 -2802
rect 7022 -2840 7056 -2838
rect 7022 -2925 7056 -2906
rect 7280 -2736 7314 -2717
rect 7280 -2804 7314 -2802
rect 7280 -2840 7314 -2838
rect 7280 -2925 7314 -2906
rect 7538 -2736 7572 -2717
rect 7538 -2804 7572 -2802
rect 7538 -2840 7572 -2838
rect 7538 -2925 7572 -2906
rect 7796 -2736 7830 -2717
rect 7796 -2804 7830 -2802
rect 7796 -2840 7830 -2838
rect 7796 -2925 7830 -2906
rect 7990 -2736 8024 -2717
rect 7990 -2804 8024 -2802
rect 7990 -2840 8024 -2838
rect 7990 -2925 8024 -2906
rect 8248 -2736 8282 -2717
rect 8248 -2804 8282 -2802
rect 8248 -2840 8282 -2838
rect 8248 -2925 8282 -2906
rect 8506 -2736 8540 -2717
rect 8506 -2804 8540 -2802
rect 8506 -2840 8540 -2838
rect 8506 -2925 8540 -2906
rect 8764 -2736 8798 -2717
rect 8764 -2804 8798 -2802
rect 8764 -2840 8798 -2838
rect 8764 -2925 8798 -2906
rect 9022 -2736 9056 -2717
rect 9022 -2804 9056 -2802
rect 9022 -2840 9056 -2838
rect 9022 -2925 9056 -2906
rect 9216 -2736 9250 -2717
rect 9216 -2804 9250 -2802
rect 9216 -2840 9250 -2838
rect 9216 -2925 9250 -2906
rect 9474 -2736 9508 -2717
rect 9474 -2804 9508 -2802
rect 9474 -2840 9508 -2838
rect 9474 -2925 9508 -2906
rect 9589 -2785 9623 -2755
rect 9589 -2857 9623 -2823
rect 9589 -2925 9623 -2891
rect 872 -2993 906 -2963
rect 872 -3061 906 -3035
rect 872 -3129 906 -3107
rect 872 -3197 906 -3179
rect 872 -3265 906 -3251
rect 5230 -2963 5231 -2925
rect 5230 -2993 5265 -2963
rect 5230 -3035 5231 -2993
rect 5230 -3061 5265 -3035
rect 5230 -3107 5231 -3061
rect 5230 -3129 5265 -3107
rect 5230 -3179 5231 -3129
rect 5230 -3197 5265 -3179
rect 5230 -3251 5231 -3197
rect 5230 -3265 5265 -3251
rect 5230 -3299 5231 -3265
rect 9589 -2993 9623 -2963
rect 9589 -3061 9623 -3035
rect 9589 -3129 9623 -3107
rect 9589 -3197 9623 -3179
rect 9589 -3265 9623 -3251
rect 906 -3323 993 -3299
rect 872 -3333 993 -3323
rect 1027 -3333 1061 -3299
rect 1095 -3333 1129 -3299
rect 1163 -3333 1197 -3299
rect 1231 -3333 1265 -3299
rect 1299 -3333 1333 -3299
rect 1367 -3333 1401 -3299
rect 1435 -3333 1469 -3299
rect 1503 -3333 1537 -3299
rect 1571 -3333 1605 -3299
rect 1639 -3333 1673 -3299
rect 1707 -3333 1741 -3299
rect 1775 -3333 1809 -3299
rect 1843 -3333 1877 -3299
rect 1911 -3333 1945 -3299
rect 1979 -3333 2013 -3299
rect 2047 -3333 2081 -3299
rect 2115 -3333 2149 -3299
rect 2183 -3333 2217 -3299
rect 2251 -3333 2285 -3299
rect 2319 -3333 2353 -3299
rect 2387 -3333 2421 -3299
rect 2455 -3333 2489 -3299
rect 2523 -3333 2557 -3299
rect 2591 -3333 2625 -3299
rect 2659 -3333 2693 -3299
rect 2727 -3333 2761 -3299
rect 2795 -3333 2829 -3299
rect 2863 -3333 2897 -3299
rect 2931 -3333 2965 -3299
rect 2999 -3333 3033 -3299
rect 3067 -3333 3101 -3299
rect 3135 -3333 3169 -3299
rect 3203 -3333 3237 -3299
rect 3271 -3333 3305 -3299
rect 3339 -3333 3373 -3299
rect 3407 -3333 3441 -3299
rect 3475 -3333 3509 -3299
rect 3543 -3333 3577 -3299
rect 3611 -3333 3645 -3299
rect 3679 -3333 3713 -3299
rect 3747 -3333 3781 -3299
rect 3815 -3333 3849 -3299
rect 3883 -3333 3917 -3299
rect 3951 -3333 3985 -3299
rect 4019 -3333 4053 -3299
rect 4087 -3333 4121 -3299
rect 4155 -3333 4189 -3299
rect 4223 -3333 4257 -3299
rect 4291 -3333 4325 -3299
rect 4359 -3333 4393 -3299
rect 4427 -3333 4461 -3299
rect 4495 -3333 4529 -3299
rect 4563 -3333 4597 -3299
rect 4631 -3333 4665 -3299
rect 4699 -3333 4733 -3299
rect 4767 -3333 4801 -3299
rect 4835 -3333 4869 -3299
rect 4903 -3333 4937 -3299
rect 4971 -3333 5005 -3299
rect 5039 -3333 5073 -3299
rect 5107 -3323 5231 -3299
rect 5265 -3323 5388 -3299
rect 5107 -3333 5388 -3323
rect 5422 -3333 5456 -3299
rect 5490 -3333 5524 -3299
rect 5558 -3333 5592 -3299
rect 5626 -3333 5660 -3299
rect 5694 -3333 5728 -3299
rect 5762 -3333 5796 -3299
rect 5830 -3333 5864 -3299
rect 5898 -3333 5932 -3299
rect 5966 -3333 6000 -3299
rect 6034 -3333 6068 -3299
rect 6102 -3333 6136 -3299
rect 6170 -3333 6204 -3299
rect 6238 -3333 6272 -3299
rect 6306 -3333 6340 -3299
rect 6374 -3333 6408 -3299
rect 6442 -3333 6476 -3299
rect 6510 -3333 6544 -3299
rect 6578 -3333 6612 -3299
rect 6646 -3333 6680 -3299
rect 6714 -3333 6748 -3299
rect 6782 -3333 6816 -3299
rect 6850 -3333 6884 -3299
rect 6918 -3333 6952 -3299
rect 6986 -3333 7020 -3299
rect 7054 -3333 7088 -3299
rect 7122 -3333 7156 -3299
rect 7190 -3333 7224 -3299
rect 7258 -3333 7292 -3299
rect 7326 -3333 7360 -3299
rect 7394 -3333 7428 -3299
rect 7462 -3333 7496 -3299
rect 7530 -3333 7564 -3299
rect 7598 -3333 7632 -3299
rect 7666 -3333 7700 -3299
rect 7734 -3333 7768 -3299
rect 7802 -3333 7836 -3299
rect 7870 -3333 7904 -3299
rect 7938 -3333 7972 -3299
rect 8006 -3333 8040 -3299
rect 8074 -3333 8108 -3299
rect 8142 -3333 8176 -3299
rect 8210 -3333 8244 -3299
rect 8278 -3333 8312 -3299
rect 8346 -3333 8380 -3299
rect 8414 -3333 8448 -3299
rect 8482 -3333 8516 -3299
rect 8550 -3333 8584 -3299
rect 8618 -3333 8652 -3299
rect 8686 -3333 8720 -3299
rect 8754 -3333 8788 -3299
rect 8822 -3333 8856 -3299
rect 8890 -3333 8924 -3299
rect 8958 -3333 8992 -3299
rect 9026 -3333 9060 -3299
rect 9094 -3333 9128 -3299
rect 9162 -3333 9196 -3299
rect 9230 -3333 9264 -3299
rect 9298 -3333 9332 -3299
rect 9366 -3333 9400 -3299
rect 9434 -3333 9468 -3299
rect 9502 -3323 9589 -3299
rect 9502 -3333 9623 -3323
rect 872 -3401 906 -3395
rect 872 -3469 906 -3467
rect 872 -3505 906 -3503
rect 872 -3577 906 -3571
rect 872 -3649 906 -3639
rect 5230 -3395 5231 -3333
rect 5230 -3401 5265 -3395
rect 5230 -3467 5231 -3401
rect 5230 -3469 5265 -3467
rect 5230 -3503 5231 -3469
rect 5230 -3505 5265 -3503
rect 5230 -3571 5231 -3505
rect 5230 -3577 5265 -3571
rect 5230 -3639 5231 -3577
rect 5230 -3649 5265 -3639
rect 5230 -3707 5231 -3649
rect 9589 -3401 9623 -3395
rect 9589 -3469 9623 -3467
rect 9589 -3505 9623 -3503
rect 9589 -3577 9623 -3571
rect 9589 -3649 9623 -3639
rect 872 -3721 906 -3707
rect 872 -3793 906 -3775
rect 872 -3865 906 -3843
rect 872 -3937 906 -3899
rect 987 -3726 1021 -3707
rect 987 -3794 1021 -3792
rect 987 -3830 1021 -3828
rect 987 -3915 1021 -3896
rect 1245 -3726 1279 -3707
rect 1245 -3794 1279 -3792
rect 1245 -3830 1279 -3828
rect 1245 -3915 1279 -3896
rect 1439 -3726 1473 -3707
rect 1439 -3794 1473 -3792
rect 1439 -3830 1473 -3828
rect 1439 -3915 1473 -3896
rect 1697 -3726 1731 -3707
rect 1697 -3794 1731 -3792
rect 1697 -3830 1731 -3828
rect 1697 -3915 1731 -3896
rect 1955 -3726 1989 -3707
rect 1955 -3794 1989 -3792
rect 1955 -3830 1989 -3828
rect 1955 -3915 1989 -3896
rect 2213 -3726 2247 -3707
rect 2213 -3794 2247 -3792
rect 2213 -3830 2247 -3828
rect 2213 -3915 2247 -3896
rect 2471 -3726 2505 -3707
rect 2471 -3794 2505 -3792
rect 2471 -3830 2505 -3828
rect 2471 -3915 2505 -3896
rect 2665 -3726 2699 -3707
rect 2665 -3794 2699 -3792
rect 2665 -3830 2699 -3828
rect 2665 -3915 2699 -3896
rect 2923 -3726 2957 -3707
rect 2923 -3794 2957 -3792
rect 2923 -3830 2957 -3828
rect 2923 -3915 2957 -3896
rect 3181 -3726 3215 -3707
rect 3181 -3794 3215 -3792
rect 3181 -3830 3215 -3828
rect 3181 -3915 3215 -3896
rect 3439 -3726 3473 -3707
rect 3439 -3794 3473 -3792
rect 3439 -3830 3473 -3828
rect 3439 -3915 3473 -3896
rect 3633 -3726 3667 -3707
rect 3633 -3794 3667 -3792
rect 3633 -3830 3667 -3828
rect 3633 -3915 3667 -3896
rect 3891 -3726 3925 -3707
rect 3891 -3794 3925 -3792
rect 3891 -3830 3925 -3828
rect 3891 -3915 3925 -3896
rect 4149 -3726 4183 -3707
rect 4149 -3794 4183 -3792
rect 4149 -3830 4183 -3828
rect 4149 -3915 4183 -3896
rect 4407 -3726 4441 -3707
rect 4407 -3794 4441 -3792
rect 4407 -3830 4441 -3828
rect 4407 -3915 4441 -3896
rect 4665 -3726 4699 -3707
rect 4665 -3794 4699 -3792
rect 4665 -3830 4699 -3828
rect 4665 -3915 4699 -3896
rect 4859 -3726 4893 -3707
rect 4859 -3794 4893 -3792
rect 4859 -3830 4893 -3828
rect 4859 -3915 4893 -3896
rect 5117 -3726 5151 -3707
rect 5117 -3794 5151 -3792
rect 5117 -3830 5151 -3828
rect 5117 -3915 5151 -3896
rect 5230 -3721 5265 -3707
rect 5230 -3775 5231 -3721
rect 5230 -3793 5265 -3775
rect 5230 -3843 5231 -3793
rect 5230 -3865 5265 -3843
rect 5230 -3899 5231 -3865
rect 5230 -3937 5265 -3899
rect 5345 -3726 5379 -3707
rect 5345 -3794 5379 -3792
rect 5345 -3830 5379 -3828
rect 5345 -3915 5379 -3896
rect 5603 -3726 5637 -3707
rect 5603 -3794 5637 -3792
rect 5603 -3830 5637 -3828
rect 5603 -3915 5637 -3896
rect 5796 -3726 5830 -3707
rect 5796 -3794 5830 -3792
rect 5796 -3830 5830 -3828
rect 5796 -3915 5830 -3896
rect 6054 -3726 6088 -3707
rect 6054 -3794 6088 -3792
rect 6054 -3830 6088 -3828
rect 6054 -3915 6088 -3896
rect 6312 -3726 6346 -3707
rect 6312 -3794 6346 -3792
rect 6312 -3830 6346 -3828
rect 6312 -3915 6346 -3896
rect 6570 -3726 6604 -3707
rect 6570 -3794 6604 -3792
rect 6570 -3830 6604 -3828
rect 6570 -3915 6604 -3896
rect 6828 -3726 6862 -3707
rect 6828 -3794 6862 -3792
rect 6828 -3830 6862 -3828
rect 6828 -3915 6862 -3896
rect 7022 -3726 7056 -3707
rect 7022 -3794 7056 -3792
rect 7022 -3830 7056 -3828
rect 7022 -3915 7056 -3896
rect 7280 -3726 7314 -3707
rect 7280 -3794 7314 -3792
rect 7280 -3830 7314 -3828
rect 7280 -3915 7314 -3896
rect 7538 -3726 7572 -3707
rect 7538 -3794 7572 -3792
rect 7538 -3830 7572 -3828
rect 7538 -3915 7572 -3896
rect 7796 -3726 7830 -3707
rect 7796 -3794 7830 -3792
rect 7796 -3830 7830 -3828
rect 7796 -3915 7830 -3896
rect 7990 -3726 8024 -3707
rect 7990 -3794 8024 -3792
rect 7990 -3830 8024 -3828
rect 7990 -3915 8024 -3896
rect 8248 -3726 8282 -3707
rect 8248 -3794 8282 -3792
rect 8248 -3830 8282 -3828
rect 8248 -3915 8282 -3896
rect 8506 -3726 8540 -3707
rect 8506 -3794 8540 -3792
rect 8506 -3830 8540 -3828
rect 8506 -3915 8540 -3896
rect 8764 -3726 8798 -3707
rect 8764 -3794 8798 -3792
rect 8764 -3830 8798 -3828
rect 8764 -3915 8798 -3896
rect 9022 -3726 9056 -3707
rect 9022 -3794 9056 -3792
rect 9022 -3830 9056 -3828
rect 9022 -3915 9056 -3896
rect 9216 -3726 9250 -3707
rect 9216 -3794 9250 -3792
rect 9216 -3830 9250 -3828
rect 9216 -3915 9250 -3896
rect 9474 -3726 9508 -3707
rect 9474 -3794 9508 -3792
rect 9474 -3830 9508 -3828
rect 9474 -3915 9508 -3896
rect 9589 -3721 9623 -3707
rect 9589 -3793 9623 -3775
rect 9589 -3865 9623 -3843
rect 872 -4009 906 -3971
rect 1033 -3992 1080 -3958
rect 1116 -3992 1150 -3958
rect 1186 -3992 1233 -3958
rect 1485 -3992 1532 -3958
rect 1568 -3992 1602 -3958
rect 1638 -3992 1685 -3958
rect 1743 -3992 1790 -3958
rect 1826 -3992 1860 -3958
rect 1896 -3992 1943 -3958
rect 2001 -3992 2048 -3958
rect 2084 -3992 2118 -3958
rect 2154 -3992 2201 -3958
rect 2259 -3992 2306 -3958
rect 2342 -3992 2376 -3958
rect 2412 -3992 2459 -3958
rect 2711 -3992 2758 -3958
rect 2794 -3992 2828 -3958
rect 2864 -3992 2911 -3958
rect 2969 -3992 3016 -3958
rect 3052 -3992 3086 -3958
rect 3122 -3992 3169 -3958
rect 3227 -3992 3274 -3958
rect 3310 -3992 3344 -3958
rect 3380 -3992 3427 -3958
rect 3679 -3992 3726 -3958
rect 3762 -3992 3796 -3958
rect 3832 -3992 3879 -3958
rect 3937 -3992 3984 -3958
rect 4020 -3992 4054 -3958
rect 4090 -3992 4137 -3958
rect 4195 -3992 4242 -3958
rect 4278 -3992 4312 -3958
rect 4348 -3992 4395 -3958
rect 4453 -3992 4500 -3958
rect 4536 -3992 4570 -3958
rect 4606 -3992 4653 -3958
rect 4905 -3992 4952 -3958
rect 4988 -3992 5022 -3958
rect 5058 -3992 5105 -3958
rect 5230 -3971 5231 -3937
rect 9589 -3937 9623 -3899
rect 872 -4072 906 -4043
rect 5230 -4009 5265 -3971
rect 5391 -3992 5438 -3958
rect 5474 -3992 5508 -3958
rect 5544 -3992 5591 -3958
rect 5842 -3992 5889 -3958
rect 5925 -3992 5959 -3958
rect 5995 -3992 6042 -3958
rect 6100 -3992 6147 -3958
rect 6183 -3992 6217 -3958
rect 6253 -3992 6300 -3958
rect 6358 -3992 6405 -3958
rect 6441 -3992 6475 -3958
rect 6511 -3992 6558 -3958
rect 6616 -3992 6663 -3958
rect 6699 -3992 6733 -3958
rect 6769 -3992 6816 -3958
rect 7068 -3992 7115 -3958
rect 7151 -3992 7185 -3958
rect 7221 -3992 7268 -3958
rect 7326 -3992 7373 -3958
rect 7409 -3992 7443 -3958
rect 7479 -3992 7526 -3958
rect 7584 -3992 7631 -3958
rect 7667 -3992 7701 -3958
rect 7737 -3992 7784 -3958
rect 8036 -3992 8083 -3958
rect 8119 -3992 8153 -3958
rect 8189 -3992 8236 -3958
rect 8294 -3992 8341 -3958
rect 8377 -3992 8411 -3958
rect 8447 -3992 8494 -3958
rect 8552 -3992 8599 -3958
rect 8635 -3992 8669 -3958
rect 8705 -3992 8752 -3958
rect 8810 -3992 8857 -3958
rect 8893 -3992 8927 -3958
rect 8963 -3992 9010 -3958
rect 9262 -3992 9309 -3958
rect 9345 -3992 9379 -3958
rect 9415 -3992 9462 -3958
rect 5230 -4043 5231 -4009
rect 5230 -4072 5265 -4043
rect 9589 -4009 9623 -3971
rect 9589 -4072 9623 -4043
rect 872 -4106 946 -4072
rect 980 -4106 993 -4072
rect 1052 -4106 1061 -4072
rect 1124 -4106 1129 -4072
rect 1196 -4106 1197 -4072
rect 1231 -4106 1234 -4072
rect 1299 -4106 1306 -4072
rect 1367 -4106 1378 -4072
rect 1435 -4106 1450 -4072
rect 1503 -4106 1522 -4072
rect 1571 -4106 1594 -4072
rect 1639 -4106 1666 -4072
rect 1707 -4106 1738 -4072
rect 1775 -4106 1809 -4072
rect 1844 -4106 1877 -4072
rect 1916 -4106 1945 -4072
rect 1988 -4106 2013 -4072
rect 2060 -4106 2081 -4072
rect 2132 -4106 2149 -4072
rect 2204 -4106 2217 -4072
rect 2276 -4106 2285 -4072
rect 2348 -4106 2353 -4072
rect 2420 -4106 2421 -4072
rect 2455 -4106 2458 -4072
rect 2523 -4106 2530 -4072
rect 2591 -4106 2602 -4072
rect 2659 -4106 2674 -4072
rect 2727 -4106 2746 -4072
rect 2795 -4106 2818 -4072
rect 2863 -4106 2890 -4072
rect 2931 -4106 2962 -4072
rect 2999 -4106 3033 -4072
rect 3068 -4106 3101 -4072
rect 3140 -4106 3169 -4072
rect 3212 -4106 3237 -4072
rect 3284 -4106 3305 -4072
rect 3356 -4106 3373 -4072
rect 3428 -4106 3441 -4072
rect 3500 -4106 3509 -4072
rect 3572 -4106 3577 -4072
rect 3644 -4106 3645 -4072
rect 3679 -4106 3682 -4072
rect 3747 -4106 3754 -4072
rect 3815 -4106 3826 -4072
rect 3883 -4106 3898 -4072
rect 3951 -4106 3970 -4072
rect 4019 -4106 4042 -4072
rect 4087 -4106 4114 -4072
rect 4155 -4106 4186 -4072
rect 4223 -4106 4257 -4072
rect 4292 -4106 4325 -4072
rect 4364 -4106 4393 -4072
rect 4436 -4106 4461 -4072
rect 4508 -4106 4529 -4072
rect 4580 -4106 4597 -4072
rect 4652 -4106 4665 -4072
rect 4724 -4106 4733 -4072
rect 4796 -4106 4801 -4072
rect 4868 -4106 4869 -4072
rect 4903 -4106 4906 -4072
rect 4971 -4106 4978 -4072
rect 5039 -4106 5050 -4072
rect 5107 -4106 5122 -4072
rect 5156 -4106 5339 -4072
rect 5373 -4106 5388 -4072
rect 5445 -4106 5456 -4072
rect 5517 -4106 5524 -4072
rect 5589 -4106 5592 -4072
rect 5626 -4106 5627 -4072
rect 5694 -4106 5699 -4072
rect 5762 -4106 5771 -4072
rect 5830 -4106 5843 -4072
rect 5898 -4106 5915 -4072
rect 5966 -4106 5987 -4072
rect 6034 -4106 6059 -4072
rect 6102 -4106 6131 -4072
rect 6170 -4106 6203 -4072
rect 6238 -4106 6272 -4072
rect 6309 -4106 6340 -4072
rect 6381 -4106 6408 -4072
rect 6453 -4106 6476 -4072
rect 6525 -4106 6544 -4072
rect 6597 -4106 6612 -4072
rect 6669 -4106 6680 -4072
rect 6741 -4106 6748 -4072
rect 6813 -4106 6816 -4072
rect 6850 -4106 6851 -4072
rect 6918 -4106 6923 -4072
rect 6986 -4106 6995 -4072
rect 7054 -4106 7067 -4072
rect 7122 -4106 7139 -4072
rect 7190 -4106 7211 -4072
rect 7258 -4106 7283 -4072
rect 7326 -4106 7355 -4072
rect 7394 -4106 7427 -4072
rect 7462 -4106 7496 -4072
rect 7533 -4106 7564 -4072
rect 7605 -4106 7632 -4072
rect 7677 -4106 7700 -4072
rect 7749 -4106 7768 -4072
rect 7821 -4106 7836 -4072
rect 7893 -4106 7904 -4072
rect 7965 -4106 7972 -4072
rect 8037 -4106 8040 -4072
rect 8074 -4106 8075 -4072
rect 8142 -4106 8147 -4072
rect 8210 -4106 8219 -4072
rect 8278 -4106 8291 -4072
rect 8346 -4106 8363 -4072
rect 8414 -4106 8435 -4072
rect 8482 -4106 8507 -4072
rect 8550 -4106 8579 -4072
rect 8618 -4106 8651 -4072
rect 8686 -4106 8720 -4072
rect 8757 -4106 8788 -4072
rect 8829 -4106 8856 -4072
rect 8901 -4106 8924 -4072
rect 8973 -4106 8992 -4072
rect 9045 -4106 9060 -4072
rect 9117 -4106 9128 -4072
rect 9189 -4106 9196 -4072
rect 9261 -4106 9264 -4072
rect 9298 -4106 9299 -4072
rect 9366 -4106 9371 -4072
rect 9434 -4106 9443 -4072
rect 9502 -4106 9515 -4072
rect 9549 -4106 9623 -4072
rect 872 -4135 906 -4106
rect 872 -4207 906 -4169
rect 5230 -4135 5265 -4106
rect 5230 -4169 5231 -4135
rect 1033 -4220 1080 -4186
rect 1116 -4220 1150 -4186
rect 1186 -4220 1233 -4186
rect 1485 -4220 1532 -4186
rect 1568 -4220 1602 -4186
rect 1638 -4220 1685 -4186
rect 1743 -4220 1790 -4186
rect 1826 -4220 1860 -4186
rect 1896 -4220 1943 -4186
rect 2001 -4220 2048 -4186
rect 2084 -4220 2118 -4186
rect 2154 -4220 2201 -4186
rect 2259 -4220 2306 -4186
rect 2342 -4220 2376 -4186
rect 2412 -4220 2459 -4186
rect 2711 -4220 2758 -4186
rect 2794 -4220 2828 -4186
rect 2864 -4220 2911 -4186
rect 2969 -4220 3016 -4186
rect 3052 -4220 3086 -4186
rect 3122 -4220 3169 -4186
rect 3227 -4220 3274 -4186
rect 3310 -4220 3344 -4186
rect 3380 -4220 3427 -4186
rect 3679 -4220 3726 -4186
rect 3762 -4220 3796 -4186
rect 3832 -4220 3879 -4186
rect 3937 -4220 3984 -4186
rect 4020 -4220 4054 -4186
rect 4090 -4220 4137 -4186
rect 4195 -4220 4242 -4186
rect 4278 -4220 4312 -4186
rect 4348 -4220 4395 -4186
rect 4453 -4220 4500 -4186
rect 4536 -4220 4570 -4186
rect 4606 -4220 4653 -4186
rect 4905 -4220 4952 -4186
rect 4988 -4220 5022 -4186
rect 5058 -4220 5105 -4186
rect 5230 -4207 5265 -4169
rect 9589 -4135 9623 -4106
rect 872 -4279 906 -4241
rect 5230 -4241 5231 -4207
rect 5391 -4220 5438 -4186
rect 5474 -4220 5508 -4186
rect 5544 -4220 5591 -4186
rect 5842 -4220 5889 -4186
rect 5925 -4220 5959 -4186
rect 5995 -4220 6042 -4186
rect 6100 -4220 6147 -4186
rect 6183 -4220 6217 -4186
rect 6253 -4220 6300 -4186
rect 6358 -4220 6405 -4186
rect 6441 -4220 6475 -4186
rect 6511 -4220 6558 -4186
rect 6616 -4220 6663 -4186
rect 6699 -4220 6733 -4186
rect 6769 -4220 6816 -4186
rect 7068 -4220 7115 -4186
rect 7151 -4220 7185 -4186
rect 7221 -4220 7268 -4186
rect 7326 -4220 7373 -4186
rect 7409 -4220 7443 -4186
rect 7479 -4220 7526 -4186
rect 7584 -4220 7631 -4186
rect 7667 -4220 7701 -4186
rect 7737 -4220 7784 -4186
rect 8036 -4220 8083 -4186
rect 8119 -4220 8153 -4186
rect 8189 -4220 8236 -4186
rect 8294 -4220 8341 -4186
rect 8377 -4220 8411 -4186
rect 8447 -4220 8494 -4186
rect 8552 -4220 8599 -4186
rect 8635 -4220 8669 -4186
rect 8705 -4220 8752 -4186
rect 8810 -4220 8857 -4186
rect 8893 -4220 8927 -4186
rect 8963 -4220 9010 -4186
rect 9262 -4220 9309 -4186
rect 9345 -4220 9379 -4186
rect 9415 -4220 9462 -4186
rect 9589 -4207 9623 -4169
rect 872 -4335 906 -4313
rect 872 -4403 906 -4385
rect 872 -4471 906 -4457
rect 987 -4282 1021 -4263
rect 987 -4350 1021 -4348
rect 987 -4386 1021 -4384
rect 987 -4471 1021 -4452
rect 1245 -4282 1279 -4263
rect 1245 -4350 1279 -4348
rect 1245 -4386 1279 -4384
rect 1245 -4471 1279 -4452
rect 1439 -4282 1473 -4263
rect 1439 -4350 1473 -4348
rect 1439 -4386 1473 -4384
rect 1439 -4471 1473 -4452
rect 1697 -4282 1731 -4263
rect 1697 -4350 1731 -4348
rect 1697 -4386 1731 -4384
rect 1697 -4471 1731 -4452
rect 1955 -4282 1989 -4263
rect 1955 -4350 1989 -4348
rect 1955 -4386 1989 -4384
rect 1955 -4471 1989 -4452
rect 2213 -4282 2247 -4263
rect 2213 -4350 2247 -4348
rect 2213 -4386 2247 -4384
rect 2213 -4471 2247 -4452
rect 2471 -4282 2505 -4263
rect 2471 -4350 2505 -4348
rect 2471 -4386 2505 -4384
rect 2471 -4471 2505 -4452
rect 2665 -4282 2699 -4263
rect 2665 -4350 2699 -4348
rect 2665 -4386 2699 -4384
rect 2665 -4471 2699 -4452
rect 2923 -4282 2957 -4263
rect 2923 -4350 2957 -4348
rect 2923 -4386 2957 -4384
rect 2923 -4471 2957 -4452
rect 3181 -4282 3215 -4263
rect 3181 -4350 3215 -4348
rect 3181 -4386 3215 -4384
rect 3181 -4471 3215 -4452
rect 3439 -4282 3473 -4263
rect 3439 -4350 3473 -4348
rect 3439 -4386 3473 -4384
rect 3439 -4471 3473 -4452
rect 3633 -4282 3667 -4263
rect 3633 -4350 3667 -4348
rect 3633 -4386 3667 -4384
rect 3633 -4471 3667 -4452
rect 3891 -4282 3925 -4263
rect 3891 -4350 3925 -4348
rect 3891 -4386 3925 -4384
rect 3891 -4471 3925 -4452
rect 4149 -4282 4183 -4263
rect 4149 -4350 4183 -4348
rect 4149 -4386 4183 -4384
rect 4149 -4471 4183 -4452
rect 4407 -4282 4441 -4263
rect 4407 -4350 4441 -4348
rect 4407 -4386 4441 -4384
rect 4407 -4471 4441 -4452
rect 4665 -4282 4699 -4263
rect 4665 -4350 4699 -4348
rect 4665 -4386 4699 -4384
rect 4665 -4471 4699 -4452
rect 4859 -4282 4893 -4263
rect 4859 -4350 4893 -4348
rect 4859 -4386 4893 -4384
rect 4859 -4471 4893 -4452
rect 5117 -4282 5151 -4263
rect 5117 -4350 5151 -4348
rect 5117 -4386 5151 -4384
rect 5117 -4471 5151 -4452
rect 5230 -4279 5265 -4241
rect 5230 -4313 5231 -4279
rect 5230 -4335 5265 -4313
rect 5230 -4385 5231 -4335
rect 5230 -4403 5265 -4385
rect 5230 -4457 5231 -4403
rect 5230 -4471 5265 -4457
rect 5345 -4282 5379 -4263
rect 5345 -4350 5379 -4348
rect 5345 -4386 5379 -4384
rect 5345 -4471 5379 -4452
rect 5603 -4282 5637 -4263
rect 5603 -4350 5637 -4348
rect 5603 -4386 5637 -4384
rect 5603 -4471 5637 -4452
rect 5796 -4282 5830 -4263
rect 5796 -4350 5830 -4348
rect 5796 -4386 5830 -4384
rect 5796 -4471 5830 -4452
rect 6054 -4282 6088 -4263
rect 6054 -4350 6088 -4348
rect 6054 -4386 6088 -4384
rect 6054 -4471 6088 -4452
rect 6312 -4282 6346 -4263
rect 6312 -4350 6346 -4348
rect 6312 -4386 6346 -4384
rect 6312 -4471 6346 -4452
rect 6570 -4282 6604 -4263
rect 6570 -4350 6604 -4348
rect 6570 -4386 6604 -4384
rect 6570 -4471 6604 -4452
rect 6828 -4282 6862 -4263
rect 6828 -4350 6862 -4348
rect 6828 -4386 6862 -4384
rect 6828 -4471 6862 -4452
rect 7022 -4282 7056 -4263
rect 7022 -4350 7056 -4348
rect 7022 -4386 7056 -4384
rect 7022 -4471 7056 -4452
rect 7280 -4282 7314 -4263
rect 7280 -4350 7314 -4348
rect 7280 -4386 7314 -4384
rect 7280 -4471 7314 -4452
rect 7538 -4282 7572 -4263
rect 7538 -4350 7572 -4348
rect 7538 -4386 7572 -4384
rect 7538 -4471 7572 -4452
rect 7796 -4282 7830 -4263
rect 7796 -4350 7830 -4348
rect 7796 -4386 7830 -4384
rect 7796 -4471 7830 -4452
rect 7990 -4282 8024 -4263
rect 7990 -4350 8024 -4348
rect 7990 -4386 8024 -4384
rect 7990 -4471 8024 -4452
rect 8248 -4282 8282 -4263
rect 8248 -4350 8282 -4348
rect 8248 -4386 8282 -4384
rect 8248 -4471 8282 -4452
rect 8506 -4282 8540 -4263
rect 8506 -4350 8540 -4348
rect 8506 -4386 8540 -4384
rect 8506 -4471 8540 -4452
rect 8764 -4282 8798 -4263
rect 8764 -4350 8798 -4348
rect 8764 -4386 8798 -4384
rect 8764 -4471 8798 -4452
rect 9022 -4282 9056 -4263
rect 9022 -4350 9056 -4348
rect 9022 -4386 9056 -4384
rect 9022 -4471 9056 -4452
rect 9216 -4282 9250 -4263
rect 9216 -4350 9250 -4348
rect 9216 -4386 9250 -4384
rect 9216 -4471 9250 -4452
rect 9474 -4282 9508 -4263
rect 9474 -4350 9508 -4348
rect 9474 -4386 9508 -4384
rect 9474 -4471 9508 -4452
rect 9589 -4279 9623 -4241
rect 9589 -4335 9623 -4313
rect 9589 -4403 9623 -4385
rect 9589 -4471 9623 -4457
rect 872 -4539 906 -4529
rect 872 -4607 906 -4601
rect 872 -4675 906 -4673
rect 872 -4711 906 -4709
rect 872 -4783 906 -4777
rect 5230 -4529 5231 -4471
rect 5230 -4539 5265 -4529
rect 5230 -4601 5231 -4539
rect 5230 -4607 5265 -4601
rect 5230 -4673 5231 -4607
rect 5230 -4675 5265 -4673
rect 5230 -4709 5231 -4675
rect 5230 -4711 5265 -4709
rect 5230 -4777 5231 -4711
rect 5230 -4783 5265 -4777
rect 5230 -4845 5231 -4783
rect 9589 -4539 9623 -4529
rect 9589 -4607 9623 -4601
rect 9589 -4675 9623 -4673
rect 9589 -4711 9623 -4709
rect 9589 -4783 9623 -4777
rect 872 -4855 993 -4845
rect 906 -4879 993 -4855
rect 1027 -4879 1061 -4845
rect 1095 -4879 1129 -4845
rect 1163 -4879 1197 -4845
rect 1231 -4879 1265 -4845
rect 1299 -4879 1333 -4845
rect 1367 -4879 1401 -4845
rect 1435 -4879 1469 -4845
rect 1503 -4879 1537 -4845
rect 1571 -4879 1605 -4845
rect 1639 -4879 1673 -4845
rect 1707 -4879 1741 -4845
rect 1775 -4879 1809 -4845
rect 1843 -4879 1877 -4845
rect 1911 -4879 1945 -4845
rect 1979 -4879 2013 -4845
rect 2047 -4879 2081 -4845
rect 2115 -4879 2149 -4845
rect 2183 -4879 2217 -4845
rect 2251 -4879 2285 -4845
rect 2319 -4879 2353 -4845
rect 2387 -4879 2421 -4845
rect 2455 -4879 2489 -4845
rect 2523 -4879 2557 -4845
rect 2591 -4879 2625 -4845
rect 2659 -4879 2693 -4845
rect 2727 -4879 2761 -4845
rect 2795 -4879 2829 -4845
rect 2863 -4879 2897 -4845
rect 2931 -4879 2965 -4845
rect 2999 -4879 3033 -4845
rect 3067 -4879 3101 -4845
rect 3135 -4879 3169 -4845
rect 3203 -4879 3237 -4845
rect 3271 -4879 3305 -4845
rect 3339 -4879 3373 -4845
rect 3407 -4879 3441 -4845
rect 3475 -4879 3509 -4845
rect 3543 -4879 3577 -4845
rect 3611 -4879 3645 -4845
rect 3679 -4879 3713 -4845
rect 3747 -4879 3781 -4845
rect 3815 -4879 3849 -4845
rect 3883 -4879 3917 -4845
rect 3951 -4879 3985 -4845
rect 4019 -4879 4053 -4845
rect 4087 -4879 4121 -4845
rect 4155 -4879 4189 -4845
rect 4223 -4879 4257 -4845
rect 4291 -4879 4325 -4845
rect 4359 -4879 4393 -4845
rect 4427 -4879 4461 -4845
rect 4495 -4879 4529 -4845
rect 4563 -4879 4597 -4845
rect 4631 -4879 4665 -4845
rect 4699 -4879 4733 -4845
rect 4767 -4879 4801 -4845
rect 4835 -4879 4869 -4845
rect 4903 -4879 4937 -4845
rect 4971 -4879 5005 -4845
rect 5039 -4879 5073 -4845
rect 5107 -4855 5388 -4845
rect 5107 -4879 5231 -4855
rect 5265 -4879 5388 -4855
rect 5422 -4879 5456 -4845
rect 5490 -4879 5524 -4845
rect 5558 -4879 5592 -4845
rect 5626 -4879 5660 -4845
rect 5694 -4879 5728 -4845
rect 5762 -4879 5796 -4845
rect 5830 -4879 5864 -4845
rect 5898 -4879 5932 -4845
rect 5966 -4879 6000 -4845
rect 6034 -4879 6068 -4845
rect 6102 -4879 6136 -4845
rect 6170 -4879 6204 -4845
rect 6238 -4879 6272 -4845
rect 6306 -4879 6340 -4845
rect 6374 -4879 6408 -4845
rect 6442 -4879 6476 -4845
rect 6510 -4879 6544 -4845
rect 6578 -4879 6612 -4845
rect 6646 -4879 6680 -4845
rect 6714 -4879 6748 -4845
rect 6782 -4879 6816 -4845
rect 6850 -4879 6884 -4845
rect 6918 -4879 6952 -4845
rect 6986 -4879 7020 -4845
rect 7054 -4879 7088 -4845
rect 7122 -4879 7156 -4845
rect 7190 -4879 7224 -4845
rect 7258 -4879 7292 -4845
rect 7326 -4879 7360 -4845
rect 7394 -4879 7428 -4845
rect 7462 -4879 7496 -4845
rect 7530 -4879 7564 -4845
rect 7598 -4879 7632 -4845
rect 7666 -4879 7700 -4845
rect 7734 -4879 7768 -4845
rect 7802 -4879 7836 -4845
rect 7870 -4879 7904 -4845
rect 7938 -4879 7972 -4845
rect 8006 -4879 8040 -4845
rect 8074 -4879 8108 -4845
rect 8142 -4879 8176 -4845
rect 8210 -4879 8244 -4845
rect 8278 -4879 8312 -4845
rect 8346 -4879 8380 -4845
rect 8414 -4879 8448 -4845
rect 8482 -4879 8516 -4845
rect 8550 -4879 8584 -4845
rect 8618 -4879 8652 -4845
rect 8686 -4879 8720 -4845
rect 8754 -4879 8788 -4845
rect 8822 -4879 8856 -4845
rect 8890 -4879 8924 -4845
rect 8958 -4879 8992 -4845
rect 9026 -4879 9060 -4845
rect 9094 -4879 9128 -4845
rect 9162 -4879 9196 -4845
rect 9230 -4879 9264 -4845
rect 9298 -4879 9332 -4845
rect 9366 -4879 9400 -4845
rect 9434 -4879 9468 -4845
rect 9502 -4855 9623 -4845
rect 9502 -4879 9589 -4855
rect 872 -4927 906 -4913
rect 872 -4999 906 -4981
rect 872 -5071 906 -5049
rect 872 -5143 906 -5117
rect 872 -5215 906 -5185
rect 5230 -4913 5231 -4879
rect 5230 -4927 5265 -4913
rect 5230 -4981 5231 -4927
rect 5230 -4999 5265 -4981
rect 5230 -5049 5231 -4999
rect 5230 -5071 5265 -5049
rect 5230 -5117 5231 -5071
rect 5230 -5143 5265 -5117
rect 5230 -5185 5231 -5143
rect 5230 -5215 5265 -5185
rect 5230 -5253 5231 -5215
rect 9589 -4927 9623 -4913
rect 9589 -4999 9623 -4981
rect 9589 -5071 9623 -5049
rect 9589 -5143 9623 -5117
rect 9589 -5215 9623 -5185
rect 872 -5287 906 -5253
rect 872 -5355 906 -5321
rect 872 -5423 906 -5393
rect 987 -5272 1021 -5253
rect 987 -5340 1021 -5338
rect 987 -5376 1021 -5374
rect 987 -5461 1021 -5442
rect 1245 -5272 1279 -5253
rect 1245 -5340 1279 -5338
rect 1245 -5376 1279 -5374
rect 1245 -5461 1279 -5442
rect 1439 -5272 1473 -5253
rect 1439 -5340 1473 -5338
rect 1439 -5376 1473 -5374
rect 1439 -5461 1473 -5442
rect 1697 -5272 1731 -5253
rect 1697 -5340 1731 -5338
rect 1697 -5376 1731 -5374
rect 1697 -5461 1731 -5442
rect 1955 -5272 1989 -5253
rect 1955 -5340 1989 -5338
rect 1955 -5376 1989 -5374
rect 1955 -5461 1989 -5442
rect 2213 -5272 2247 -5253
rect 2213 -5340 2247 -5338
rect 2213 -5376 2247 -5374
rect 2213 -5461 2247 -5442
rect 2471 -5272 2505 -5253
rect 2471 -5340 2505 -5338
rect 2471 -5376 2505 -5374
rect 2471 -5461 2505 -5442
rect 2665 -5272 2699 -5253
rect 2665 -5340 2699 -5338
rect 2665 -5376 2699 -5374
rect 2665 -5461 2699 -5442
rect 2923 -5272 2957 -5253
rect 2923 -5340 2957 -5338
rect 2923 -5376 2957 -5374
rect 2923 -5461 2957 -5442
rect 3181 -5272 3215 -5253
rect 3181 -5340 3215 -5338
rect 3181 -5376 3215 -5374
rect 3181 -5461 3215 -5442
rect 3439 -5272 3473 -5253
rect 3439 -5340 3473 -5338
rect 3439 -5376 3473 -5374
rect 3439 -5461 3473 -5442
rect 3633 -5272 3667 -5253
rect 3633 -5340 3667 -5338
rect 3633 -5376 3667 -5374
rect 3633 -5461 3667 -5442
rect 3891 -5272 3925 -5253
rect 3891 -5340 3925 -5338
rect 3891 -5376 3925 -5374
rect 3891 -5461 3925 -5442
rect 4149 -5272 4183 -5253
rect 4149 -5340 4183 -5338
rect 4149 -5376 4183 -5374
rect 4149 -5461 4183 -5442
rect 4407 -5272 4441 -5253
rect 4407 -5340 4441 -5338
rect 4407 -5376 4441 -5374
rect 4407 -5461 4441 -5442
rect 4665 -5272 4699 -5253
rect 4665 -5340 4699 -5338
rect 4665 -5376 4699 -5374
rect 4665 -5461 4699 -5442
rect 4859 -5272 4893 -5253
rect 4859 -5340 4893 -5338
rect 4859 -5376 4893 -5374
rect 4859 -5461 4893 -5442
rect 5117 -5272 5151 -5253
rect 5117 -5340 5151 -5338
rect 5117 -5376 5151 -5374
rect 5117 -5461 5151 -5442
rect 5230 -5287 5265 -5253
rect 5230 -5321 5231 -5287
rect 5230 -5355 5265 -5321
rect 5230 -5393 5231 -5355
rect 5230 -5423 5265 -5393
rect 872 -5491 906 -5465
rect 5230 -5465 5231 -5423
rect 5345 -5272 5379 -5253
rect 5345 -5340 5379 -5338
rect 5345 -5376 5379 -5374
rect 5345 -5461 5379 -5442
rect 5603 -5272 5637 -5253
rect 5603 -5340 5637 -5338
rect 5603 -5376 5637 -5374
rect 5603 -5461 5637 -5442
rect 5796 -5272 5830 -5253
rect 5796 -5340 5830 -5338
rect 5796 -5376 5830 -5374
rect 5796 -5461 5830 -5442
rect 6054 -5272 6088 -5253
rect 6054 -5340 6088 -5338
rect 6054 -5376 6088 -5374
rect 6054 -5461 6088 -5442
rect 6312 -5272 6346 -5253
rect 6312 -5340 6346 -5338
rect 6312 -5376 6346 -5374
rect 6312 -5461 6346 -5442
rect 6570 -5272 6604 -5253
rect 6570 -5340 6604 -5338
rect 6570 -5376 6604 -5374
rect 6570 -5461 6604 -5442
rect 6828 -5272 6862 -5253
rect 6828 -5340 6862 -5338
rect 6828 -5376 6862 -5374
rect 6828 -5461 6862 -5442
rect 7022 -5272 7056 -5253
rect 7022 -5340 7056 -5338
rect 7022 -5376 7056 -5374
rect 7022 -5461 7056 -5442
rect 7280 -5272 7314 -5253
rect 7280 -5340 7314 -5338
rect 7280 -5376 7314 -5374
rect 7280 -5461 7314 -5442
rect 7538 -5272 7572 -5253
rect 7538 -5340 7572 -5338
rect 7538 -5376 7572 -5374
rect 7538 -5461 7572 -5442
rect 7796 -5272 7830 -5253
rect 7796 -5340 7830 -5338
rect 7796 -5376 7830 -5374
rect 7796 -5461 7830 -5442
rect 7990 -5272 8024 -5253
rect 7990 -5340 8024 -5338
rect 7990 -5376 8024 -5374
rect 7990 -5461 8024 -5442
rect 8248 -5272 8282 -5253
rect 8248 -5340 8282 -5338
rect 8248 -5376 8282 -5374
rect 8248 -5461 8282 -5442
rect 8506 -5272 8540 -5253
rect 8506 -5340 8540 -5338
rect 8506 -5376 8540 -5374
rect 8506 -5461 8540 -5442
rect 8764 -5272 8798 -5253
rect 8764 -5340 8798 -5338
rect 8764 -5376 8798 -5374
rect 8764 -5461 8798 -5442
rect 9022 -5272 9056 -5253
rect 9022 -5340 9056 -5338
rect 9022 -5376 9056 -5374
rect 9022 -5461 9056 -5442
rect 9216 -5272 9250 -5253
rect 9216 -5340 9250 -5338
rect 9216 -5376 9250 -5374
rect 9216 -5461 9250 -5442
rect 9474 -5272 9508 -5253
rect 9474 -5340 9508 -5338
rect 9474 -5376 9508 -5374
rect 9474 -5461 9508 -5442
rect 9589 -5287 9623 -5253
rect 9589 -5355 9623 -5321
rect 9589 -5423 9623 -5393
rect 5230 -5491 5265 -5465
rect 872 -5559 906 -5537
rect 1033 -5538 1080 -5504
rect 1116 -5538 1150 -5504
rect 1186 -5538 1233 -5504
rect 1485 -5538 1532 -5504
rect 1568 -5538 1602 -5504
rect 1638 -5538 1685 -5504
rect 1743 -5538 1790 -5504
rect 1826 -5538 1860 -5504
rect 1896 -5538 1943 -5504
rect 2001 -5538 2048 -5504
rect 2084 -5538 2118 -5504
rect 2154 -5538 2201 -5504
rect 2259 -5538 2306 -5504
rect 2342 -5538 2376 -5504
rect 2412 -5538 2459 -5504
rect 2711 -5538 2758 -5504
rect 2794 -5538 2828 -5504
rect 2864 -5538 2911 -5504
rect 2969 -5538 3016 -5504
rect 3052 -5538 3086 -5504
rect 3122 -5538 3169 -5504
rect 3227 -5538 3274 -5504
rect 3310 -5538 3344 -5504
rect 3380 -5538 3427 -5504
rect 3679 -5538 3726 -5504
rect 3762 -5538 3796 -5504
rect 3832 -5538 3879 -5504
rect 3937 -5538 3984 -5504
rect 4020 -5538 4054 -5504
rect 4090 -5538 4137 -5504
rect 4195 -5538 4242 -5504
rect 4278 -5538 4312 -5504
rect 4348 -5538 4395 -5504
rect 4453 -5538 4500 -5504
rect 4536 -5538 4570 -5504
rect 4606 -5538 4653 -5504
rect 4905 -5538 4952 -5504
rect 4988 -5538 5022 -5504
rect 5058 -5538 5105 -5504
rect 5230 -5537 5231 -5491
rect 9589 -5491 9623 -5465
rect 872 -5627 906 -5609
rect 872 -5695 906 -5681
rect 872 -5763 906 -5753
rect 872 -5831 906 -5825
rect 5230 -5559 5265 -5537
rect 5391 -5538 5438 -5504
rect 5474 -5538 5508 -5504
rect 5544 -5538 5591 -5504
rect 5842 -5538 5889 -5504
rect 5925 -5538 5959 -5504
rect 5995 -5538 6042 -5504
rect 6100 -5538 6147 -5504
rect 6183 -5538 6217 -5504
rect 6253 -5538 6300 -5504
rect 6358 -5538 6405 -5504
rect 6441 -5538 6475 -5504
rect 6511 -5538 6558 -5504
rect 6616 -5538 6663 -5504
rect 6699 -5538 6733 -5504
rect 6769 -5538 6816 -5504
rect 7068 -5538 7115 -5504
rect 7151 -5538 7185 -5504
rect 7221 -5538 7268 -5504
rect 7326 -5538 7373 -5504
rect 7409 -5538 7443 -5504
rect 7479 -5538 7526 -5504
rect 7584 -5538 7631 -5504
rect 7667 -5538 7701 -5504
rect 7737 -5538 7784 -5504
rect 8036 -5538 8083 -5504
rect 8119 -5538 8153 -5504
rect 8189 -5538 8236 -5504
rect 8294 -5538 8341 -5504
rect 8377 -5538 8411 -5504
rect 8447 -5538 8494 -5504
rect 8552 -5538 8599 -5504
rect 8635 -5538 8669 -5504
rect 8705 -5538 8752 -5504
rect 8810 -5538 8857 -5504
rect 8893 -5538 8927 -5504
rect 8963 -5538 9010 -5504
rect 9262 -5538 9309 -5504
rect 9345 -5538 9379 -5504
rect 9415 -5538 9462 -5504
rect 5230 -5609 5231 -5559
rect 5230 -5627 5265 -5609
rect 5230 -5681 5231 -5627
rect 5230 -5695 5265 -5681
rect 5230 -5753 5231 -5695
rect 5230 -5763 5265 -5753
rect 5230 -5825 5231 -5763
rect 5230 -5831 5265 -5825
rect 872 -5899 906 -5897
rect 1033 -5900 1080 -5866
rect 1116 -5900 1150 -5866
rect 1186 -5900 1233 -5866
rect 1485 -5900 1532 -5866
rect 1568 -5900 1602 -5866
rect 1638 -5900 1685 -5866
rect 1743 -5900 1790 -5866
rect 1826 -5900 1860 -5866
rect 1896 -5900 1943 -5866
rect 2001 -5900 2048 -5866
rect 2084 -5900 2118 -5866
rect 2154 -5900 2201 -5866
rect 2259 -5900 2306 -5866
rect 2342 -5900 2376 -5866
rect 2412 -5900 2459 -5866
rect 2711 -5900 2758 -5866
rect 2794 -5900 2828 -5866
rect 2864 -5900 2911 -5866
rect 2969 -5900 3016 -5866
rect 3052 -5900 3086 -5866
rect 3122 -5900 3169 -5866
rect 3227 -5900 3274 -5866
rect 3310 -5900 3344 -5866
rect 3380 -5900 3427 -5866
rect 3679 -5900 3726 -5866
rect 3762 -5900 3796 -5866
rect 3832 -5900 3879 -5866
rect 3937 -5900 3984 -5866
rect 4020 -5900 4054 -5866
rect 4090 -5900 4137 -5866
rect 4195 -5900 4242 -5866
rect 4278 -5900 4312 -5866
rect 4348 -5900 4395 -5866
rect 4453 -5900 4500 -5866
rect 4536 -5900 4570 -5866
rect 4606 -5900 4653 -5866
rect 4905 -5900 4952 -5866
rect 4988 -5900 5022 -5866
rect 5058 -5900 5105 -5866
rect 5230 -5897 5231 -5831
rect 9589 -5559 9623 -5537
rect 9589 -5627 9623 -5609
rect 9589 -5695 9623 -5681
rect 9589 -5763 9623 -5753
rect 9589 -5831 9623 -5825
rect 5230 -5899 5265 -5897
rect 872 -5935 906 -5933
rect 5230 -5933 5231 -5899
rect 5391 -5900 5438 -5866
rect 5474 -5900 5508 -5866
rect 5544 -5900 5591 -5866
rect 5842 -5900 5889 -5866
rect 5925 -5900 5959 -5866
rect 5995 -5900 6042 -5866
rect 6100 -5900 6147 -5866
rect 6183 -5900 6217 -5866
rect 6253 -5900 6300 -5866
rect 6358 -5900 6405 -5866
rect 6441 -5900 6475 -5866
rect 6511 -5900 6558 -5866
rect 6616 -5900 6663 -5866
rect 6699 -5900 6733 -5866
rect 6769 -5900 6816 -5866
rect 7068 -5900 7115 -5866
rect 7151 -5900 7185 -5866
rect 7221 -5900 7268 -5866
rect 7326 -5900 7373 -5866
rect 7409 -5900 7443 -5866
rect 7479 -5900 7526 -5866
rect 7584 -5900 7631 -5866
rect 7667 -5900 7701 -5866
rect 7737 -5900 7784 -5866
rect 8036 -5900 8083 -5866
rect 8119 -5900 8153 -5866
rect 8189 -5900 8236 -5866
rect 8294 -5900 8341 -5866
rect 8377 -5900 8411 -5866
rect 8447 -5900 8494 -5866
rect 8552 -5900 8599 -5866
rect 8635 -5900 8669 -5866
rect 8705 -5900 8752 -5866
rect 8810 -5900 8857 -5866
rect 8893 -5900 8927 -5866
rect 8963 -5900 9010 -5866
rect 9262 -5900 9309 -5866
rect 9345 -5900 9379 -5866
rect 9415 -5900 9462 -5866
rect 9589 -5899 9623 -5897
rect 5230 -5935 5265 -5933
rect 872 -6007 906 -6001
rect 872 -6079 906 -6069
rect 872 -6151 906 -6137
rect 987 -5962 1021 -5943
rect 987 -6030 1021 -6028
rect 987 -6066 1021 -6064
rect 987 -6151 1021 -6132
rect 1245 -5962 1279 -5943
rect 1245 -6030 1279 -6028
rect 1245 -6066 1279 -6064
rect 1245 -6151 1279 -6132
rect 1439 -5962 1473 -5943
rect 1439 -6030 1473 -6028
rect 1439 -6066 1473 -6064
rect 1439 -6151 1473 -6132
rect 1697 -5962 1731 -5943
rect 1697 -6030 1731 -6028
rect 1697 -6066 1731 -6064
rect 1697 -6151 1731 -6132
rect 1955 -5962 1989 -5943
rect 1955 -6030 1989 -6028
rect 1955 -6066 1989 -6064
rect 1955 -6151 1989 -6132
rect 2213 -5962 2247 -5943
rect 2213 -6030 2247 -6028
rect 2213 -6066 2247 -6064
rect 2213 -6151 2247 -6132
rect 2471 -5962 2505 -5943
rect 2471 -6030 2505 -6028
rect 2471 -6066 2505 -6064
rect 2471 -6151 2505 -6132
rect 2665 -5962 2699 -5943
rect 2665 -6030 2699 -6028
rect 2665 -6066 2699 -6064
rect 2665 -6151 2699 -6132
rect 2923 -5962 2957 -5943
rect 2923 -6030 2957 -6028
rect 2923 -6066 2957 -6064
rect 2923 -6151 2957 -6132
rect 3181 -5962 3215 -5943
rect 3181 -6030 3215 -6028
rect 3181 -6066 3215 -6064
rect 3181 -6151 3215 -6132
rect 3439 -5962 3473 -5943
rect 3439 -6030 3473 -6028
rect 3439 -6066 3473 -6064
rect 3439 -6151 3473 -6132
rect 3633 -5962 3667 -5943
rect 3633 -6030 3667 -6028
rect 3633 -6066 3667 -6064
rect 3633 -6151 3667 -6132
rect 3891 -5962 3925 -5943
rect 3891 -6030 3925 -6028
rect 3891 -6066 3925 -6064
rect 3891 -6151 3925 -6132
rect 4149 -5962 4183 -5943
rect 4149 -6030 4183 -6028
rect 4149 -6066 4183 -6064
rect 4149 -6151 4183 -6132
rect 4407 -5962 4441 -5943
rect 4407 -6030 4441 -6028
rect 4407 -6066 4441 -6064
rect 4407 -6151 4441 -6132
rect 4665 -5962 4699 -5943
rect 4665 -6030 4699 -6028
rect 4665 -6066 4699 -6064
rect 4665 -6151 4699 -6132
rect 4859 -5962 4893 -5943
rect 4859 -6030 4893 -6028
rect 4859 -6066 4893 -6064
rect 4859 -6151 4893 -6132
rect 5117 -5962 5151 -5943
rect 5117 -6030 5151 -6028
rect 5117 -6066 5151 -6064
rect 5117 -6151 5151 -6132
rect 5230 -6001 5231 -5935
rect 9589 -5935 9623 -5933
rect 5230 -6007 5265 -6001
rect 5230 -6069 5231 -6007
rect 5230 -6079 5265 -6069
rect 5230 -6137 5231 -6079
rect 5230 -6151 5265 -6137
rect 5345 -5962 5379 -5943
rect 5345 -6030 5379 -6028
rect 5345 -6066 5379 -6064
rect 5345 -6151 5379 -6132
rect 5603 -5962 5637 -5943
rect 5603 -6030 5637 -6028
rect 5603 -6066 5637 -6064
rect 5603 -6151 5637 -6132
rect 5796 -5962 5830 -5943
rect 5796 -6030 5830 -6028
rect 5796 -6066 5830 -6064
rect 5796 -6151 5830 -6132
rect 6054 -5962 6088 -5943
rect 6054 -6030 6088 -6028
rect 6054 -6066 6088 -6064
rect 6054 -6151 6088 -6132
rect 6312 -5962 6346 -5943
rect 6312 -6030 6346 -6028
rect 6312 -6066 6346 -6064
rect 6312 -6151 6346 -6132
rect 6570 -5962 6604 -5943
rect 6570 -6030 6604 -6028
rect 6570 -6066 6604 -6064
rect 6570 -6151 6604 -6132
rect 6828 -5962 6862 -5943
rect 6828 -6030 6862 -6028
rect 6828 -6066 6862 -6064
rect 6828 -6151 6862 -6132
rect 7022 -5962 7056 -5943
rect 7022 -6030 7056 -6028
rect 7022 -6066 7056 -6064
rect 7022 -6151 7056 -6132
rect 7280 -5962 7314 -5943
rect 7280 -6030 7314 -6028
rect 7280 -6066 7314 -6064
rect 7280 -6151 7314 -6132
rect 7538 -5962 7572 -5943
rect 7538 -6030 7572 -6028
rect 7538 -6066 7572 -6064
rect 7538 -6151 7572 -6132
rect 7796 -5962 7830 -5943
rect 7796 -6030 7830 -6028
rect 7796 -6066 7830 -6064
rect 7796 -6151 7830 -6132
rect 7990 -5962 8024 -5943
rect 7990 -6030 8024 -6028
rect 7990 -6066 8024 -6064
rect 7990 -6151 8024 -6132
rect 8248 -5962 8282 -5943
rect 8248 -6030 8282 -6028
rect 8248 -6066 8282 -6064
rect 8248 -6151 8282 -6132
rect 8506 -5962 8540 -5943
rect 8506 -6030 8540 -6028
rect 8506 -6066 8540 -6064
rect 8506 -6151 8540 -6132
rect 8764 -5962 8798 -5943
rect 8764 -6030 8798 -6028
rect 8764 -6066 8798 -6064
rect 8764 -6151 8798 -6132
rect 9022 -5962 9056 -5943
rect 9022 -6030 9056 -6028
rect 9022 -6066 9056 -6064
rect 9022 -6151 9056 -6132
rect 9216 -5962 9250 -5943
rect 9216 -6030 9250 -6028
rect 9216 -6066 9250 -6064
rect 9216 -6151 9250 -6132
rect 9474 -5962 9508 -5943
rect 9474 -6030 9508 -6028
rect 9474 -6066 9508 -6064
rect 9474 -6151 9508 -6132
rect 9589 -6007 9623 -6001
rect 9589 -6079 9623 -6069
rect 9589 -6151 9623 -6137
rect 872 -6223 906 -6205
rect 872 -6295 906 -6273
rect 872 -6367 906 -6341
rect 872 -6439 906 -6409
rect 872 -6511 906 -6473
rect 5230 -6205 5231 -6151
rect 5230 -6223 5265 -6205
rect 5230 -6273 5231 -6223
rect 5230 -6295 5265 -6273
rect 5230 -6341 5231 -6295
rect 5230 -6367 5265 -6341
rect 5230 -6409 5231 -6367
rect 5230 -6439 5265 -6409
rect 5230 -6473 5231 -6439
rect 5230 -6511 5265 -6473
rect 9589 -6223 9623 -6205
rect 9589 -6295 9623 -6273
rect 9589 -6367 9623 -6341
rect 9589 -6439 9623 -6409
rect 9589 -6511 9623 -6473
rect 906 -6545 993 -6511
rect 1027 -6545 1061 -6511
rect 1095 -6545 1129 -6511
rect 1163 -6545 1197 -6511
rect 1231 -6545 1265 -6511
rect 1299 -6545 1333 -6511
rect 1367 -6545 1401 -6511
rect 1435 -6545 1469 -6511
rect 1503 -6545 1537 -6511
rect 1571 -6545 1605 -6511
rect 1639 -6545 1673 -6511
rect 1707 -6545 1741 -6511
rect 1775 -6545 1809 -6511
rect 1843 -6545 1877 -6511
rect 1911 -6545 1945 -6511
rect 1979 -6545 2013 -6511
rect 2047 -6545 2081 -6511
rect 2115 -6545 2149 -6511
rect 2183 -6545 2217 -6511
rect 2251 -6545 2285 -6511
rect 2319 -6545 2353 -6511
rect 2387 -6545 2421 -6511
rect 2455 -6545 2489 -6511
rect 2523 -6545 2557 -6511
rect 2591 -6545 2625 -6511
rect 2659 -6545 2693 -6511
rect 2727 -6545 2761 -6511
rect 2795 -6545 2829 -6511
rect 2863 -6545 2897 -6511
rect 2931 -6545 2965 -6511
rect 2999 -6545 3033 -6511
rect 3067 -6545 3101 -6511
rect 3135 -6545 3169 -6511
rect 3203 -6545 3237 -6511
rect 3271 -6545 3305 -6511
rect 3339 -6545 3373 -6511
rect 3407 -6545 3441 -6511
rect 3475 -6545 3509 -6511
rect 3543 -6545 3577 -6511
rect 3611 -6545 3645 -6511
rect 3679 -6545 3713 -6511
rect 3747 -6545 3781 -6511
rect 3815 -6545 3849 -6511
rect 3883 -6545 3917 -6511
rect 3951 -6545 3985 -6511
rect 4019 -6545 4053 -6511
rect 4087 -6545 4121 -6511
rect 4155 -6545 4189 -6511
rect 4223 -6545 4257 -6511
rect 4291 -6545 4325 -6511
rect 4359 -6545 4393 -6511
rect 4427 -6545 4461 -6511
rect 4495 -6545 4529 -6511
rect 4563 -6545 4597 -6511
rect 4631 -6545 4665 -6511
rect 4699 -6545 4733 -6511
rect 4767 -6545 4801 -6511
rect 4835 -6545 4869 -6511
rect 4903 -6545 4937 -6511
rect 4971 -6545 5005 -6511
rect 5039 -6545 5073 -6511
rect 5107 -6545 5231 -6511
rect 5265 -6545 5388 -6511
rect 5422 -6545 5456 -6511
rect 5490 -6545 5524 -6511
rect 5558 -6545 5592 -6511
rect 5626 -6545 5660 -6511
rect 5694 -6545 5728 -6511
rect 5762 -6545 5796 -6511
rect 5830 -6545 5864 -6511
rect 5898 -6545 5932 -6511
rect 5966 -6545 6000 -6511
rect 6034 -6545 6068 -6511
rect 6102 -6545 6136 -6511
rect 6170 -6545 6204 -6511
rect 6238 -6545 6272 -6511
rect 6306 -6545 6340 -6511
rect 6374 -6545 6408 -6511
rect 6442 -6545 6476 -6511
rect 6510 -6545 6544 -6511
rect 6578 -6545 6612 -6511
rect 6646 -6545 6680 -6511
rect 6714 -6545 6748 -6511
rect 6782 -6545 6816 -6511
rect 6850 -6545 6884 -6511
rect 6918 -6545 6952 -6511
rect 6986 -6545 7020 -6511
rect 7054 -6545 7088 -6511
rect 7122 -6545 7156 -6511
rect 7190 -6545 7224 -6511
rect 7258 -6545 7292 -6511
rect 7326 -6545 7360 -6511
rect 7394 -6545 7428 -6511
rect 7462 -6545 7496 -6511
rect 7530 -6545 7564 -6511
rect 7598 -6545 7632 -6511
rect 7666 -6545 7700 -6511
rect 7734 -6545 7768 -6511
rect 7802 -6545 7836 -6511
rect 7870 -6545 7904 -6511
rect 7938 -6545 7972 -6511
rect 8006 -6545 8040 -6511
rect 8074 -6545 8108 -6511
rect 8142 -6545 8176 -6511
rect 8210 -6545 8244 -6511
rect 8278 -6545 8312 -6511
rect 8346 -6545 8380 -6511
rect 8414 -6545 8448 -6511
rect 8482 -6545 8516 -6511
rect 8550 -6545 8584 -6511
rect 8618 -6545 8652 -6511
rect 8686 -6545 8720 -6511
rect 8754 -6545 8788 -6511
rect 8822 -6545 8856 -6511
rect 8890 -6545 8924 -6511
rect 8958 -6545 8992 -6511
rect 9026 -6545 9060 -6511
rect 9094 -6545 9128 -6511
rect 9162 -6545 9196 -6511
rect 9230 -6545 9264 -6511
rect 9298 -6545 9332 -6511
rect 9366 -6545 9400 -6511
rect 9434 -6545 9468 -6511
rect 9502 -6545 9589 -6511
rect 872 -6583 906 -6545
rect 872 -6647 906 -6617
rect 872 -6715 906 -6689
rect 872 -6783 906 -6761
rect 872 -6851 906 -6833
rect 5230 -6583 5265 -6545
rect 5230 -6617 5231 -6583
rect 5230 -6647 5265 -6617
rect 5230 -6689 5231 -6647
rect 5230 -6715 5265 -6689
rect 5230 -6761 5231 -6715
rect 5230 -6783 5265 -6761
rect 5230 -6833 5231 -6783
rect 5230 -6851 5265 -6833
rect 872 -6919 906 -6905
rect 872 -6987 906 -6977
rect 872 -7055 906 -7049
rect 987 -6919 1021 -6900
rect 987 -6987 1021 -6985
rect 987 -7023 1021 -7021
rect 987 -7108 1021 -7089
rect 1245 -6919 1279 -6900
rect 1245 -6987 1279 -6985
rect 1245 -7023 1279 -7021
rect 1245 -7108 1279 -7089
rect 1439 -6919 1473 -6900
rect 1439 -6987 1473 -6985
rect 1439 -7023 1473 -7021
rect 1439 -7108 1473 -7089
rect 1697 -6919 1731 -6900
rect 1697 -6987 1731 -6985
rect 1697 -7023 1731 -7021
rect 1697 -7108 1731 -7089
rect 1955 -6919 1989 -6900
rect 1955 -6987 1989 -6985
rect 1955 -7023 1989 -7021
rect 1955 -7108 1989 -7089
rect 2213 -6919 2247 -6900
rect 2213 -6987 2247 -6985
rect 2213 -7023 2247 -7021
rect 2213 -7108 2247 -7089
rect 2471 -6919 2505 -6900
rect 2471 -6987 2505 -6985
rect 2471 -7023 2505 -7021
rect 2471 -7108 2505 -7089
rect 2665 -6919 2699 -6900
rect 2665 -6987 2699 -6985
rect 2665 -7023 2699 -7021
rect 2665 -7108 2699 -7089
rect 2923 -6919 2957 -6900
rect 2923 -6987 2957 -6985
rect 2923 -7023 2957 -7021
rect 2923 -7108 2957 -7089
rect 3181 -6919 3215 -6900
rect 3181 -6987 3215 -6985
rect 3181 -7023 3215 -7021
rect 3181 -7108 3215 -7089
rect 3439 -6919 3473 -6900
rect 3439 -6987 3473 -6985
rect 3439 -7023 3473 -7021
rect 3439 -7108 3473 -7089
rect 3633 -6919 3667 -6900
rect 3633 -6987 3667 -6985
rect 3633 -7023 3667 -7021
rect 3633 -7108 3667 -7089
rect 3891 -6919 3925 -6900
rect 3891 -6987 3925 -6985
rect 3891 -7023 3925 -7021
rect 3891 -7108 3925 -7089
rect 4149 -6919 4183 -6900
rect 4149 -6987 4183 -6985
rect 4149 -7023 4183 -7021
rect 4149 -7108 4183 -7089
rect 4407 -6919 4441 -6900
rect 4407 -6987 4441 -6985
rect 4407 -7023 4441 -7021
rect 4407 -7108 4441 -7089
rect 4665 -6919 4699 -6900
rect 4665 -6987 4699 -6985
rect 4665 -7023 4699 -7021
rect 4665 -7108 4699 -7089
rect 4859 -6919 4893 -6900
rect 4859 -6987 4893 -6985
rect 4859 -7023 4893 -7021
rect 4859 -7108 4893 -7089
rect 5117 -6919 5151 -6900
rect 5117 -6987 5151 -6985
rect 5117 -7023 5151 -7021
rect 5117 -7108 5151 -7089
rect 5230 -6905 5231 -6851
rect 9589 -6583 9623 -6545
rect 9589 -6647 9623 -6617
rect 9589 -6715 9623 -6689
rect 9589 -6783 9623 -6761
rect 9589 -6851 9623 -6833
rect 5230 -6919 5265 -6905
rect 5230 -6977 5231 -6919
rect 5230 -6987 5265 -6977
rect 5230 -7049 5231 -6987
rect 5230 -7055 5265 -7049
rect 872 -7123 906 -7121
rect 5230 -7121 5231 -7055
rect 5345 -6919 5379 -6900
rect 5345 -6987 5379 -6985
rect 5345 -7023 5379 -7021
rect 5345 -7108 5379 -7089
rect 5603 -6919 5637 -6900
rect 5603 -6987 5637 -6985
rect 5603 -7023 5637 -7021
rect 5603 -7108 5637 -7089
rect 5796 -6919 5830 -6900
rect 5796 -6987 5830 -6985
rect 5796 -7023 5830 -7021
rect 5796 -7108 5830 -7089
rect 6054 -6919 6088 -6900
rect 6054 -6987 6088 -6985
rect 6054 -7023 6088 -7021
rect 6054 -7108 6088 -7089
rect 6312 -6919 6346 -6900
rect 6312 -6987 6346 -6985
rect 6312 -7023 6346 -7021
rect 6312 -7108 6346 -7089
rect 6570 -6919 6604 -6900
rect 6570 -6987 6604 -6985
rect 6570 -7023 6604 -7021
rect 6570 -7108 6604 -7089
rect 6828 -6919 6862 -6900
rect 6828 -6987 6862 -6985
rect 6828 -7023 6862 -7021
rect 6828 -7108 6862 -7089
rect 7022 -6919 7056 -6900
rect 7022 -6987 7056 -6985
rect 7022 -7023 7056 -7021
rect 7022 -7108 7056 -7089
rect 7280 -6919 7314 -6900
rect 7280 -6987 7314 -6985
rect 7280 -7023 7314 -7021
rect 7280 -7108 7314 -7089
rect 7538 -6919 7572 -6900
rect 7538 -6987 7572 -6985
rect 7538 -7023 7572 -7021
rect 7538 -7108 7572 -7089
rect 7796 -6919 7830 -6900
rect 7796 -6987 7830 -6985
rect 7796 -7023 7830 -7021
rect 7796 -7108 7830 -7089
rect 7990 -6919 8024 -6900
rect 7990 -6987 8024 -6985
rect 7990 -7023 8024 -7021
rect 7990 -7108 8024 -7089
rect 8248 -6919 8282 -6900
rect 8248 -6987 8282 -6985
rect 8248 -7023 8282 -7021
rect 8248 -7108 8282 -7089
rect 8506 -6919 8540 -6900
rect 8506 -6987 8540 -6985
rect 8506 -7023 8540 -7021
rect 8506 -7108 8540 -7089
rect 8764 -6919 8798 -6900
rect 8764 -6987 8798 -6985
rect 8764 -7023 8798 -7021
rect 8764 -7108 8798 -7089
rect 9022 -6919 9056 -6900
rect 9022 -6987 9056 -6985
rect 9022 -7023 9056 -7021
rect 9022 -7108 9056 -7089
rect 9216 -6919 9250 -6900
rect 9216 -6987 9250 -6985
rect 9216 -7023 9250 -7021
rect 9216 -7108 9250 -7089
rect 9474 -6919 9508 -6900
rect 9474 -6987 9508 -6985
rect 9474 -7023 9508 -7021
rect 9474 -7108 9508 -7089
rect 9589 -6919 9623 -6905
rect 9589 -6987 9623 -6977
rect 9589 -7055 9623 -7049
rect 5230 -7123 5265 -7121
rect 872 -7159 906 -7157
rect 1033 -7185 1080 -7151
rect 1116 -7185 1150 -7151
rect 1186 -7185 1233 -7151
rect 1485 -7185 1532 -7151
rect 1568 -7185 1602 -7151
rect 1638 -7185 1685 -7151
rect 1743 -7185 1790 -7151
rect 1826 -7185 1860 -7151
rect 1896 -7185 1943 -7151
rect 2001 -7185 2048 -7151
rect 2084 -7185 2118 -7151
rect 2154 -7185 2201 -7151
rect 2259 -7185 2306 -7151
rect 2342 -7185 2376 -7151
rect 2412 -7185 2459 -7151
rect 2711 -7185 2758 -7151
rect 2794 -7185 2828 -7151
rect 2864 -7185 2911 -7151
rect 2969 -7185 3016 -7151
rect 3052 -7185 3086 -7151
rect 3122 -7185 3169 -7151
rect 3227 -7185 3274 -7151
rect 3310 -7185 3344 -7151
rect 3380 -7185 3427 -7151
rect 3679 -7185 3726 -7151
rect 3762 -7185 3796 -7151
rect 3832 -7185 3879 -7151
rect 3937 -7185 3984 -7151
rect 4020 -7185 4054 -7151
rect 4090 -7185 4137 -7151
rect 4195 -7185 4242 -7151
rect 4278 -7185 4312 -7151
rect 4348 -7185 4395 -7151
rect 4453 -7185 4500 -7151
rect 4536 -7185 4570 -7151
rect 4606 -7185 4653 -7151
rect 4905 -7185 4952 -7151
rect 4988 -7185 5022 -7151
rect 5058 -7185 5105 -7151
rect 5230 -7157 5231 -7123
rect 9589 -7123 9623 -7121
rect 5230 -7159 5265 -7157
rect 872 -7231 906 -7225
rect 872 -7303 906 -7293
rect 872 -7375 906 -7361
rect 872 -7447 906 -7429
rect 872 -7519 906 -7497
rect 5230 -7225 5231 -7159
rect 5391 -7185 5438 -7151
rect 5474 -7185 5508 -7151
rect 5544 -7185 5591 -7151
rect 5842 -7185 5889 -7151
rect 5925 -7185 5959 -7151
rect 5995 -7185 6042 -7151
rect 6100 -7185 6147 -7151
rect 6183 -7185 6217 -7151
rect 6253 -7185 6300 -7151
rect 6358 -7185 6405 -7151
rect 6441 -7185 6475 -7151
rect 6511 -7185 6558 -7151
rect 6616 -7185 6663 -7151
rect 6699 -7185 6733 -7151
rect 6769 -7185 6816 -7151
rect 7068 -7185 7115 -7151
rect 7151 -7185 7185 -7151
rect 7221 -7185 7268 -7151
rect 7326 -7185 7373 -7151
rect 7409 -7185 7443 -7151
rect 7479 -7185 7526 -7151
rect 7584 -7185 7631 -7151
rect 7667 -7185 7701 -7151
rect 7737 -7185 7784 -7151
rect 8036 -7185 8083 -7151
rect 8119 -7185 8153 -7151
rect 8189 -7185 8236 -7151
rect 8294 -7185 8341 -7151
rect 8377 -7185 8411 -7151
rect 8447 -7185 8494 -7151
rect 8552 -7185 8599 -7151
rect 8635 -7185 8669 -7151
rect 8705 -7185 8752 -7151
rect 8810 -7185 8857 -7151
rect 8893 -7185 8927 -7151
rect 8963 -7185 9010 -7151
rect 9262 -7185 9309 -7151
rect 9345 -7185 9379 -7151
rect 9415 -7185 9462 -7151
rect 9589 -7159 9623 -7157
rect 5230 -7231 5265 -7225
rect 5230 -7293 5231 -7231
rect 5230 -7303 5265 -7293
rect 5230 -7361 5231 -7303
rect 5230 -7375 5265 -7361
rect 5230 -7429 5231 -7375
rect 5230 -7447 5265 -7429
rect 5230 -7497 5231 -7447
rect 1033 -7547 1080 -7513
rect 1116 -7547 1150 -7513
rect 1186 -7547 1233 -7513
rect 1485 -7547 1532 -7513
rect 1568 -7547 1602 -7513
rect 1638 -7547 1685 -7513
rect 1743 -7547 1790 -7513
rect 1826 -7547 1860 -7513
rect 1896 -7547 1943 -7513
rect 2001 -7547 2048 -7513
rect 2084 -7547 2118 -7513
rect 2154 -7547 2201 -7513
rect 2259 -7547 2306 -7513
rect 2342 -7547 2376 -7513
rect 2412 -7547 2459 -7513
rect 2711 -7547 2758 -7513
rect 2794 -7547 2828 -7513
rect 2864 -7547 2911 -7513
rect 2969 -7547 3016 -7513
rect 3052 -7547 3086 -7513
rect 3122 -7547 3169 -7513
rect 3227 -7547 3274 -7513
rect 3310 -7547 3344 -7513
rect 3380 -7547 3427 -7513
rect 3679 -7547 3726 -7513
rect 3762 -7547 3796 -7513
rect 3832 -7547 3879 -7513
rect 3937 -7547 3984 -7513
rect 4020 -7547 4054 -7513
rect 4090 -7547 4137 -7513
rect 4195 -7547 4242 -7513
rect 4278 -7547 4312 -7513
rect 4348 -7547 4395 -7513
rect 4453 -7547 4500 -7513
rect 4536 -7547 4570 -7513
rect 4606 -7547 4653 -7513
rect 4905 -7547 4952 -7513
rect 4988 -7547 5022 -7513
rect 5058 -7547 5105 -7513
rect 5230 -7519 5265 -7497
rect 9589 -7231 9623 -7225
rect 9589 -7303 9623 -7293
rect 9589 -7375 9623 -7361
rect 9589 -7447 9623 -7429
rect 872 -7591 906 -7565
rect 5230 -7565 5231 -7519
rect 5391 -7547 5438 -7513
rect 5474 -7547 5508 -7513
rect 5544 -7547 5591 -7513
rect 5842 -7547 5889 -7513
rect 5925 -7547 5959 -7513
rect 5995 -7547 6042 -7513
rect 6100 -7547 6147 -7513
rect 6183 -7547 6217 -7513
rect 6253 -7547 6300 -7513
rect 6358 -7547 6405 -7513
rect 6441 -7547 6475 -7513
rect 6511 -7547 6558 -7513
rect 6616 -7547 6663 -7513
rect 6699 -7547 6733 -7513
rect 6769 -7547 6816 -7513
rect 7068 -7547 7115 -7513
rect 7151 -7547 7185 -7513
rect 7221 -7547 7268 -7513
rect 7326 -7547 7373 -7513
rect 7409 -7547 7443 -7513
rect 7479 -7547 7526 -7513
rect 7584 -7547 7631 -7513
rect 7667 -7547 7701 -7513
rect 7737 -7547 7784 -7513
rect 8036 -7547 8083 -7513
rect 8119 -7547 8153 -7513
rect 8189 -7547 8236 -7513
rect 8294 -7547 8341 -7513
rect 8377 -7547 8411 -7513
rect 8447 -7547 8494 -7513
rect 8552 -7547 8599 -7513
rect 8635 -7547 8669 -7513
rect 8705 -7547 8752 -7513
rect 8810 -7547 8857 -7513
rect 8893 -7547 8927 -7513
rect 8963 -7547 9010 -7513
rect 9262 -7547 9309 -7513
rect 9345 -7547 9379 -7513
rect 9415 -7547 9462 -7513
rect 9589 -7519 9623 -7497
rect 872 -7663 906 -7633
rect 872 -7735 906 -7701
rect 872 -7803 906 -7769
rect 987 -7609 1021 -7590
rect 987 -7677 1021 -7675
rect 987 -7713 1021 -7711
rect 987 -7798 1021 -7779
rect 1245 -7609 1279 -7590
rect 1245 -7677 1279 -7675
rect 1245 -7713 1279 -7711
rect 1245 -7798 1279 -7779
rect 1439 -7609 1473 -7590
rect 1439 -7677 1473 -7675
rect 1439 -7713 1473 -7711
rect 1439 -7798 1473 -7779
rect 1697 -7609 1731 -7590
rect 1697 -7677 1731 -7675
rect 1697 -7713 1731 -7711
rect 1697 -7798 1731 -7779
rect 1955 -7609 1989 -7590
rect 1955 -7677 1989 -7675
rect 1955 -7713 1989 -7711
rect 1955 -7798 1989 -7779
rect 2213 -7609 2247 -7590
rect 2213 -7677 2247 -7675
rect 2213 -7713 2247 -7711
rect 2213 -7798 2247 -7779
rect 2471 -7609 2505 -7590
rect 2471 -7677 2505 -7675
rect 2471 -7713 2505 -7711
rect 2471 -7798 2505 -7779
rect 2665 -7609 2699 -7590
rect 2665 -7677 2699 -7675
rect 2665 -7713 2699 -7711
rect 2665 -7798 2699 -7779
rect 2923 -7609 2957 -7590
rect 2923 -7677 2957 -7675
rect 2923 -7713 2957 -7711
rect 2923 -7798 2957 -7779
rect 3181 -7609 3215 -7590
rect 3181 -7677 3215 -7675
rect 3181 -7713 3215 -7711
rect 3181 -7798 3215 -7779
rect 3439 -7609 3473 -7590
rect 3439 -7677 3473 -7675
rect 3439 -7713 3473 -7711
rect 3439 -7798 3473 -7779
rect 3633 -7609 3667 -7590
rect 3633 -7677 3667 -7675
rect 3633 -7713 3667 -7711
rect 3633 -7798 3667 -7779
rect 3891 -7609 3925 -7590
rect 3891 -7677 3925 -7675
rect 3891 -7713 3925 -7711
rect 3891 -7798 3925 -7779
rect 4149 -7609 4183 -7590
rect 4149 -7677 4183 -7675
rect 4149 -7713 4183 -7711
rect 4149 -7798 4183 -7779
rect 4407 -7609 4441 -7590
rect 4407 -7677 4441 -7675
rect 4407 -7713 4441 -7711
rect 4407 -7798 4441 -7779
rect 4665 -7609 4699 -7590
rect 4665 -7677 4699 -7675
rect 4665 -7713 4699 -7711
rect 4665 -7798 4699 -7779
rect 4859 -7609 4893 -7590
rect 4859 -7677 4893 -7675
rect 4859 -7713 4893 -7711
rect 4859 -7798 4893 -7779
rect 5117 -7609 5151 -7590
rect 5117 -7677 5151 -7675
rect 5117 -7713 5151 -7711
rect 5117 -7798 5151 -7779
rect 5230 -7591 5265 -7565
rect 5230 -7633 5231 -7591
rect 5230 -7663 5265 -7633
rect 5230 -7701 5231 -7663
rect 5230 -7735 5265 -7701
rect 5230 -7769 5231 -7735
rect 872 -7871 906 -7841
rect 872 -7939 906 -7913
rect 872 -8007 906 -7985
rect 872 -8075 906 -8057
rect 5230 -7803 5265 -7769
rect 5345 -7609 5379 -7590
rect 5345 -7677 5379 -7675
rect 5345 -7713 5379 -7711
rect 5345 -7798 5379 -7779
rect 5603 -7609 5637 -7590
rect 5603 -7677 5637 -7675
rect 5603 -7713 5637 -7711
rect 5603 -7798 5637 -7779
rect 5796 -7609 5830 -7590
rect 5796 -7677 5830 -7675
rect 5796 -7713 5830 -7711
rect 5796 -7798 5830 -7779
rect 6054 -7609 6088 -7590
rect 6054 -7677 6088 -7675
rect 6054 -7713 6088 -7711
rect 6054 -7798 6088 -7779
rect 6312 -7609 6346 -7590
rect 6312 -7677 6346 -7675
rect 6312 -7713 6346 -7711
rect 6312 -7798 6346 -7779
rect 6570 -7609 6604 -7590
rect 6570 -7677 6604 -7675
rect 6570 -7713 6604 -7711
rect 6570 -7798 6604 -7779
rect 6828 -7609 6862 -7590
rect 6828 -7677 6862 -7675
rect 6828 -7713 6862 -7711
rect 6828 -7798 6862 -7779
rect 7022 -7609 7056 -7590
rect 7022 -7677 7056 -7675
rect 7022 -7713 7056 -7711
rect 7022 -7798 7056 -7779
rect 7280 -7609 7314 -7590
rect 7280 -7677 7314 -7675
rect 7280 -7713 7314 -7711
rect 7280 -7798 7314 -7779
rect 7538 -7609 7572 -7590
rect 7538 -7677 7572 -7675
rect 7538 -7713 7572 -7711
rect 7538 -7798 7572 -7779
rect 7796 -7609 7830 -7590
rect 7796 -7677 7830 -7675
rect 7796 -7713 7830 -7711
rect 7796 -7798 7830 -7779
rect 7990 -7609 8024 -7590
rect 7990 -7677 8024 -7675
rect 7990 -7713 8024 -7711
rect 7990 -7798 8024 -7779
rect 8248 -7609 8282 -7590
rect 8248 -7677 8282 -7675
rect 8248 -7713 8282 -7711
rect 8248 -7798 8282 -7779
rect 8506 -7609 8540 -7590
rect 8506 -7677 8540 -7675
rect 8506 -7713 8540 -7711
rect 8506 -7798 8540 -7779
rect 8764 -7609 8798 -7590
rect 8764 -7677 8798 -7675
rect 8764 -7713 8798 -7711
rect 8764 -7798 8798 -7779
rect 9022 -7609 9056 -7590
rect 9022 -7677 9056 -7675
rect 9022 -7713 9056 -7711
rect 9022 -7798 9056 -7779
rect 9216 -7609 9250 -7590
rect 9216 -7677 9250 -7675
rect 9216 -7713 9250 -7711
rect 9216 -7798 9250 -7779
rect 9474 -7609 9508 -7590
rect 9474 -7677 9508 -7675
rect 9474 -7713 9508 -7711
rect 9474 -7798 9508 -7779
rect 9589 -7591 9623 -7565
rect 9589 -7663 9623 -7633
rect 9589 -7735 9623 -7701
rect 5230 -7841 5231 -7803
rect 5230 -7871 5265 -7841
rect 5230 -7913 5231 -7871
rect 5230 -7939 5265 -7913
rect 5230 -7985 5231 -7939
rect 5230 -8007 5265 -7985
rect 5230 -8057 5231 -8007
rect 5230 -8075 5265 -8057
rect 5230 -8109 5231 -8075
rect 9589 -7803 9623 -7769
rect 9589 -7871 9623 -7841
rect 9589 -7939 9623 -7913
rect 9589 -8007 9623 -7985
rect 9589 -8075 9623 -8057
rect 906 -8129 993 -8109
rect 872 -8143 993 -8129
rect 1027 -8143 1061 -8109
rect 1095 -8143 1129 -8109
rect 1163 -8143 1197 -8109
rect 1231 -8143 1265 -8109
rect 1299 -8143 1333 -8109
rect 1367 -8143 1401 -8109
rect 1435 -8143 1469 -8109
rect 1503 -8143 1537 -8109
rect 1571 -8143 1605 -8109
rect 1639 -8143 1673 -8109
rect 1707 -8143 1741 -8109
rect 1775 -8143 1809 -8109
rect 1843 -8143 1877 -8109
rect 1911 -8143 1945 -8109
rect 1979 -8143 2013 -8109
rect 2047 -8143 2081 -8109
rect 2115 -8143 2149 -8109
rect 2183 -8143 2217 -8109
rect 2251 -8143 2285 -8109
rect 2319 -8143 2353 -8109
rect 2387 -8143 2421 -8109
rect 2455 -8143 2489 -8109
rect 2523 -8143 2557 -8109
rect 2591 -8143 2625 -8109
rect 2659 -8143 2693 -8109
rect 2727 -8143 2761 -8109
rect 2795 -8143 2829 -8109
rect 2863 -8143 2897 -8109
rect 2931 -8143 2965 -8109
rect 2999 -8143 3033 -8109
rect 3067 -8143 3101 -8109
rect 3135 -8143 3169 -8109
rect 3203 -8143 3237 -8109
rect 3271 -8143 3305 -8109
rect 3339 -8143 3373 -8109
rect 3407 -8143 3441 -8109
rect 3475 -8143 3509 -8109
rect 3543 -8143 3577 -8109
rect 3611 -8143 3645 -8109
rect 3679 -8143 3713 -8109
rect 3747 -8143 3781 -8109
rect 3815 -8143 3849 -8109
rect 3883 -8143 3917 -8109
rect 3951 -8143 3985 -8109
rect 4019 -8143 4053 -8109
rect 4087 -8143 4121 -8109
rect 4155 -8143 4189 -8109
rect 4223 -8143 4257 -8109
rect 4291 -8143 4325 -8109
rect 4359 -8143 4393 -8109
rect 4427 -8143 4461 -8109
rect 4495 -8143 4529 -8109
rect 4563 -8143 4597 -8109
rect 4631 -8143 4665 -8109
rect 4699 -8143 4733 -8109
rect 4767 -8143 4801 -8109
rect 4835 -8143 4869 -8109
rect 4903 -8143 4937 -8109
rect 4971 -8143 5005 -8109
rect 5039 -8143 5073 -8109
rect 5107 -8129 5231 -8109
rect 5265 -8129 5388 -8109
rect 5107 -8143 5388 -8129
rect 5422 -8143 5456 -8109
rect 5490 -8143 5524 -8109
rect 5558 -8143 5592 -8109
rect 5626 -8143 5660 -8109
rect 5694 -8143 5728 -8109
rect 5762 -8143 5796 -8109
rect 5830 -8143 5864 -8109
rect 5898 -8143 5932 -8109
rect 5966 -8143 6000 -8109
rect 6034 -8143 6068 -8109
rect 6102 -8143 6136 -8109
rect 6170 -8143 6204 -8109
rect 6238 -8143 6272 -8109
rect 6306 -8143 6340 -8109
rect 6374 -8143 6408 -8109
rect 6442 -8143 6476 -8109
rect 6510 -8143 6544 -8109
rect 6578 -8143 6612 -8109
rect 6646 -8143 6680 -8109
rect 6714 -8143 6748 -8109
rect 6782 -8143 6816 -8109
rect 6850 -8143 6884 -8109
rect 6918 -8143 6952 -8109
rect 6986 -8143 7020 -8109
rect 7054 -8143 7088 -8109
rect 7122 -8143 7156 -8109
rect 7190 -8143 7224 -8109
rect 7258 -8143 7292 -8109
rect 7326 -8143 7360 -8109
rect 7394 -8143 7428 -8109
rect 7462 -8143 7496 -8109
rect 7530 -8143 7564 -8109
rect 7598 -8143 7632 -8109
rect 7666 -8143 7700 -8109
rect 7734 -8143 7768 -8109
rect 7802 -8143 7836 -8109
rect 7870 -8143 7904 -8109
rect 7938 -8143 7972 -8109
rect 8006 -8143 8040 -8109
rect 8074 -8143 8108 -8109
rect 8142 -8143 8176 -8109
rect 8210 -8143 8244 -8109
rect 8278 -8143 8312 -8109
rect 8346 -8143 8380 -8109
rect 8414 -8143 8448 -8109
rect 8482 -8143 8516 -8109
rect 8550 -8143 8584 -8109
rect 8618 -8143 8652 -8109
rect 8686 -8143 8720 -8109
rect 8754 -8143 8788 -8109
rect 8822 -8143 8856 -8109
rect 8890 -8143 8924 -8109
rect 8958 -8143 8992 -8109
rect 9026 -8143 9060 -8109
rect 9094 -8143 9128 -8109
rect 9162 -8143 9196 -8109
rect 9230 -8143 9264 -8109
rect 9298 -8143 9332 -8109
rect 9366 -8143 9400 -8109
rect 9434 -8143 9468 -8109
rect 9502 -8129 9589 -8109
rect 9502 -8143 9623 -8129
rect 872 -8211 906 -8201
rect 872 -8279 906 -8273
rect 872 -8347 906 -8345
rect 872 -8383 906 -8381
rect 872 -8455 906 -8449
rect 872 -8527 906 -8517
rect 5230 -8201 5231 -8143
rect 5230 -8211 5265 -8201
rect 5230 -8273 5231 -8211
rect 5230 -8279 5265 -8273
rect 5230 -8345 5231 -8279
rect 5230 -8347 5265 -8345
rect 5230 -8381 5231 -8347
rect 5230 -8383 5265 -8381
rect 5230 -8449 5231 -8383
rect 5230 -8455 5265 -8449
rect 5230 -8517 5231 -8455
rect 5230 -8527 5265 -8517
rect 872 -8599 906 -8585
rect 872 -8671 906 -8653
rect 872 -8743 906 -8721
rect 987 -8553 1021 -8534
rect 987 -8621 1021 -8619
rect 987 -8657 1021 -8655
rect 987 -8742 1021 -8723
rect 1245 -8553 1279 -8534
rect 1245 -8621 1279 -8619
rect 1245 -8657 1279 -8655
rect 1245 -8742 1279 -8723
rect 1439 -8553 1473 -8534
rect 1439 -8621 1473 -8619
rect 1439 -8657 1473 -8655
rect 1439 -8742 1473 -8723
rect 1697 -8553 1731 -8534
rect 1697 -8621 1731 -8619
rect 1697 -8657 1731 -8655
rect 1697 -8742 1731 -8723
rect 1955 -8553 1989 -8534
rect 1955 -8621 1989 -8619
rect 1955 -8657 1989 -8655
rect 1955 -8742 1989 -8723
rect 2213 -8553 2247 -8534
rect 2213 -8621 2247 -8619
rect 2213 -8657 2247 -8655
rect 2213 -8742 2247 -8723
rect 2471 -8553 2505 -8534
rect 2471 -8621 2505 -8619
rect 2471 -8657 2505 -8655
rect 2471 -8742 2505 -8723
rect 2665 -8553 2699 -8534
rect 2665 -8621 2699 -8619
rect 2665 -8657 2699 -8655
rect 2665 -8742 2699 -8723
rect 2923 -8553 2957 -8534
rect 2923 -8621 2957 -8619
rect 2923 -8657 2957 -8655
rect 2923 -8742 2957 -8723
rect 3181 -8553 3215 -8534
rect 3181 -8621 3215 -8619
rect 3181 -8657 3215 -8655
rect 3181 -8742 3215 -8723
rect 3439 -8553 3473 -8534
rect 3439 -8621 3473 -8619
rect 3439 -8657 3473 -8655
rect 3439 -8742 3473 -8723
rect 3633 -8553 3667 -8534
rect 3633 -8621 3667 -8619
rect 3633 -8657 3667 -8655
rect 3633 -8742 3667 -8723
rect 3891 -8553 3925 -8534
rect 3891 -8621 3925 -8619
rect 3891 -8657 3925 -8655
rect 3891 -8742 3925 -8723
rect 4149 -8553 4183 -8534
rect 4149 -8621 4183 -8619
rect 4149 -8657 4183 -8655
rect 4149 -8742 4183 -8723
rect 4407 -8553 4441 -8534
rect 4407 -8621 4441 -8619
rect 4407 -8657 4441 -8655
rect 4407 -8742 4441 -8723
rect 4665 -8553 4699 -8534
rect 4665 -8621 4699 -8619
rect 4665 -8657 4699 -8655
rect 4665 -8742 4699 -8723
rect 4859 -8553 4893 -8534
rect 4859 -8621 4893 -8619
rect 4859 -8657 4893 -8655
rect 4859 -8742 4893 -8723
rect 5117 -8553 5151 -8534
rect 5117 -8621 5151 -8619
rect 5117 -8657 5151 -8655
rect 5117 -8742 5151 -8723
rect 5230 -8585 5231 -8527
rect 9589 -8211 9623 -8201
rect 9589 -8279 9623 -8273
rect 9589 -8347 9623 -8345
rect 9589 -8383 9623 -8381
rect 9589 -8455 9623 -8449
rect 9589 -8527 9623 -8517
rect 5230 -8599 5265 -8585
rect 5230 -8653 5231 -8599
rect 5230 -8671 5265 -8653
rect 5230 -8721 5231 -8671
rect 872 -8899 906 -8777
rect 5230 -8743 5265 -8721
rect 5345 -8553 5379 -8534
rect 5345 -8621 5379 -8619
rect 5345 -8657 5379 -8655
rect 5345 -8742 5379 -8723
rect 5603 -8553 5637 -8534
rect 5603 -8621 5637 -8619
rect 5603 -8657 5637 -8655
rect 5603 -8742 5637 -8723
rect 5796 -8553 5830 -8534
rect 5796 -8621 5830 -8619
rect 5796 -8657 5830 -8655
rect 5796 -8742 5830 -8723
rect 6054 -8553 6088 -8534
rect 6054 -8621 6088 -8619
rect 6054 -8657 6088 -8655
rect 6054 -8742 6088 -8723
rect 6312 -8553 6346 -8534
rect 6312 -8621 6346 -8619
rect 6312 -8657 6346 -8655
rect 6312 -8742 6346 -8723
rect 6570 -8553 6604 -8534
rect 6570 -8621 6604 -8619
rect 6570 -8657 6604 -8655
rect 6570 -8742 6604 -8723
rect 6828 -8553 6862 -8534
rect 6828 -8621 6862 -8619
rect 6828 -8657 6862 -8655
rect 6828 -8742 6862 -8723
rect 7022 -8553 7056 -8534
rect 7022 -8621 7056 -8619
rect 7022 -8657 7056 -8655
rect 7022 -8742 7056 -8723
rect 7280 -8553 7314 -8534
rect 7280 -8621 7314 -8619
rect 7280 -8657 7314 -8655
rect 7280 -8742 7314 -8723
rect 7538 -8553 7572 -8534
rect 7538 -8621 7572 -8619
rect 7538 -8657 7572 -8655
rect 7538 -8742 7572 -8723
rect 7796 -8553 7830 -8534
rect 7796 -8621 7830 -8619
rect 7796 -8657 7830 -8655
rect 7796 -8742 7830 -8723
rect 7990 -8553 8024 -8534
rect 7990 -8621 8024 -8619
rect 7990 -8657 8024 -8655
rect 7990 -8742 8024 -8723
rect 8248 -8553 8282 -8534
rect 8248 -8621 8282 -8619
rect 8248 -8657 8282 -8655
rect 8248 -8742 8282 -8723
rect 8506 -8553 8540 -8534
rect 8506 -8621 8540 -8619
rect 8506 -8657 8540 -8655
rect 8506 -8742 8540 -8723
rect 8764 -8553 8798 -8534
rect 8764 -8621 8798 -8619
rect 8764 -8657 8798 -8655
rect 8764 -8742 8798 -8723
rect 9022 -8553 9056 -8534
rect 9022 -8621 9056 -8619
rect 9022 -8657 9056 -8655
rect 9022 -8742 9056 -8723
rect 9216 -8553 9250 -8534
rect 9216 -8621 9250 -8619
rect 9216 -8657 9250 -8655
rect 9216 -8742 9250 -8723
rect 9474 -8553 9508 -8534
rect 9474 -8621 9508 -8619
rect 9474 -8657 9508 -8655
rect 9474 -8742 9508 -8723
rect 9589 -8599 9623 -8585
rect 9589 -8671 9623 -8653
rect 5230 -8777 5231 -8743
rect 1033 -8819 1080 -8785
rect 1116 -8819 1150 -8785
rect 1186 -8819 1233 -8785
rect 1485 -8819 1532 -8785
rect 1568 -8819 1602 -8785
rect 1638 -8819 1685 -8785
rect 1743 -8819 1790 -8785
rect 1826 -8819 1860 -8785
rect 1896 -8819 1943 -8785
rect 2001 -8819 2048 -8785
rect 2084 -8819 2118 -8785
rect 2154 -8819 2201 -8785
rect 2259 -8819 2306 -8785
rect 2342 -8819 2376 -8785
rect 2412 -8819 2459 -8785
rect 2711 -8819 2758 -8785
rect 2794 -8819 2828 -8785
rect 2864 -8819 2911 -8785
rect 2969 -8819 3016 -8785
rect 3052 -8819 3086 -8785
rect 3122 -8819 3169 -8785
rect 3227 -8819 3274 -8785
rect 3310 -8819 3344 -8785
rect 3380 -8819 3427 -8785
rect 3679 -8819 3726 -8785
rect 3762 -8819 3796 -8785
rect 3832 -8819 3879 -8785
rect 3937 -8819 3984 -8785
rect 4020 -8819 4054 -8785
rect 4090 -8819 4137 -8785
rect 4195 -8819 4242 -8785
rect 4278 -8819 4312 -8785
rect 4348 -8819 4395 -8785
rect 4453 -8819 4500 -8785
rect 4536 -8819 4570 -8785
rect 4606 -8819 4653 -8785
rect 4905 -8819 4952 -8785
rect 4988 -8819 5022 -8785
rect 5058 -8819 5105 -8785
rect 5230 -8899 5265 -8777
rect 9589 -8743 9623 -8721
rect 5391 -8819 5438 -8785
rect 5474 -8819 5508 -8785
rect 5544 -8819 5591 -8785
rect 5842 -8819 5889 -8785
rect 5925 -8819 5959 -8785
rect 5995 -8819 6042 -8785
rect 6100 -8819 6147 -8785
rect 6183 -8819 6217 -8785
rect 6253 -8819 6300 -8785
rect 6358 -8819 6405 -8785
rect 6441 -8819 6475 -8785
rect 6511 -8819 6558 -8785
rect 6616 -8819 6663 -8785
rect 6699 -8819 6733 -8785
rect 6769 -8819 6816 -8785
rect 7068 -8819 7115 -8785
rect 7151 -8819 7185 -8785
rect 7221 -8819 7268 -8785
rect 7326 -8819 7373 -8785
rect 7409 -8819 7443 -8785
rect 7479 -8819 7526 -8785
rect 7584 -8819 7631 -8785
rect 7667 -8819 7701 -8785
rect 7737 -8819 7784 -8785
rect 8036 -8819 8083 -8785
rect 8119 -8819 8153 -8785
rect 8189 -8819 8236 -8785
rect 8294 -8819 8341 -8785
rect 8377 -8819 8411 -8785
rect 8447 -8819 8494 -8785
rect 8552 -8819 8599 -8785
rect 8635 -8819 8669 -8785
rect 8705 -8819 8752 -8785
rect 8810 -8819 8857 -8785
rect 8893 -8819 8927 -8785
rect 8963 -8819 9010 -8785
rect 9262 -8819 9309 -8785
rect 9345 -8819 9379 -8785
rect 9415 -8819 9462 -8785
rect 9589 -8899 9623 -8777
rect 872 -8933 946 -8899
rect 980 -8933 993 -8899
rect 1052 -8933 1061 -8899
rect 1124 -8933 1129 -8899
rect 1196 -8933 1197 -8899
rect 1231 -8933 1234 -8899
rect 1299 -8933 1306 -8899
rect 1367 -8933 1378 -8899
rect 1435 -8933 1450 -8899
rect 1503 -8933 1522 -8899
rect 1571 -8933 1594 -8899
rect 1639 -8933 1666 -8899
rect 1707 -8933 1738 -8899
rect 1775 -8933 1809 -8899
rect 1844 -8933 1877 -8899
rect 1916 -8933 1945 -8899
rect 1988 -8933 2013 -8899
rect 2060 -8933 2081 -8899
rect 2132 -8933 2149 -8899
rect 2204 -8933 2217 -8899
rect 2276 -8933 2285 -8899
rect 2348 -8933 2353 -8899
rect 2420 -8933 2421 -8899
rect 2455 -8933 2458 -8899
rect 2523 -8933 2530 -8899
rect 2591 -8933 2602 -8899
rect 2659 -8933 2674 -8899
rect 2727 -8933 2746 -8899
rect 2795 -8933 2818 -8899
rect 2863 -8933 2890 -8899
rect 2931 -8933 2962 -8899
rect 2999 -8933 3033 -8899
rect 3068 -8933 3101 -8899
rect 3140 -8933 3169 -8899
rect 3212 -8933 3237 -8899
rect 3284 -8933 3305 -8899
rect 3356 -8933 3373 -8899
rect 3428 -8933 3441 -8899
rect 3500 -8933 3509 -8899
rect 3572 -8933 3577 -8899
rect 3644 -8933 3645 -8899
rect 3679 -8933 3682 -8899
rect 3747 -8933 3754 -8899
rect 3815 -8933 3826 -8899
rect 3883 -8933 3898 -8899
rect 3951 -8933 3970 -8899
rect 4019 -8933 4042 -8899
rect 4087 -8933 4114 -8899
rect 4155 -8933 4186 -8899
rect 4223 -8933 4257 -8899
rect 4292 -8933 4325 -8899
rect 4364 -8933 4393 -8899
rect 4436 -8933 4461 -8899
rect 4508 -8933 4529 -8899
rect 4580 -8933 4597 -8899
rect 4652 -8933 4665 -8899
rect 4724 -8933 4733 -8899
rect 4796 -8933 4801 -8899
rect 4868 -8933 4869 -8899
rect 4903 -8933 4906 -8899
rect 4971 -8933 4978 -8899
rect 5039 -8933 5050 -8899
rect 5107 -8933 5122 -8899
rect 5156 -8933 5339 -8899
rect 5373 -8933 5388 -8899
rect 5445 -8933 5456 -8899
rect 5517 -8933 5524 -8899
rect 5589 -8933 5592 -8899
rect 5626 -8933 5627 -8899
rect 5694 -8933 5699 -8899
rect 5762 -8933 5771 -8899
rect 5830 -8933 5843 -8899
rect 5898 -8933 5915 -8899
rect 5966 -8933 5987 -8899
rect 6034 -8933 6059 -8899
rect 6102 -8933 6131 -8899
rect 6170 -8933 6203 -8899
rect 6238 -8933 6272 -8899
rect 6309 -8933 6340 -8899
rect 6381 -8933 6408 -8899
rect 6453 -8933 6476 -8899
rect 6525 -8933 6544 -8899
rect 6597 -8933 6612 -8899
rect 6669 -8933 6680 -8899
rect 6741 -8933 6748 -8899
rect 6813 -8933 6816 -8899
rect 6850 -8933 6851 -8899
rect 6918 -8933 6923 -8899
rect 6986 -8933 6995 -8899
rect 7054 -8933 7067 -8899
rect 7122 -8933 7139 -8899
rect 7190 -8933 7211 -8899
rect 7258 -8933 7283 -8899
rect 7326 -8933 7355 -8899
rect 7394 -8933 7427 -8899
rect 7462 -8933 7496 -8899
rect 7533 -8933 7564 -8899
rect 7605 -8933 7632 -8899
rect 7677 -8933 7700 -8899
rect 7749 -8933 7768 -8899
rect 7821 -8933 7836 -8899
rect 7893 -8933 7904 -8899
rect 7965 -8933 7972 -8899
rect 8037 -8933 8040 -8899
rect 8074 -8933 8075 -8899
rect 8142 -8933 8147 -8899
rect 8210 -8933 8219 -8899
rect 8278 -8933 8291 -8899
rect 8346 -8933 8363 -8899
rect 8414 -8933 8435 -8899
rect 8482 -8933 8507 -8899
rect 8550 -8933 8579 -8899
rect 8618 -8933 8651 -8899
rect 8686 -8933 8720 -8899
rect 8757 -8933 8788 -8899
rect 8829 -8933 8856 -8899
rect 8901 -8933 8924 -8899
rect 8973 -8933 8992 -8899
rect 9045 -8933 9060 -8899
rect 9117 -8933 9128 -8899
rect 9189 -8933 9196 -8899
rect 9261 -8933 9264 -8899
rect 9298 -8933 9299 -8899
rect 9366 -8933 9371 -8899
rect 9434 -8933 9443 -8899
rect 9502 -8933 9515 -8899
rect 9549 -8933 9623 -8899
<< viali >>
rect 946 722 980 756
rect 1018 722 1027 756
rect 1027 722 1052 756
rect 1090 722 1095 756
rect 1095 722 1124 756
rect 1162 722 1163 756
rect 1163 722 1196 756
rect 1234 722 1265 756
rect 1265 722 1268 756
rect 1306 722 1333 756
rect 1333 722 1340 756
rect 1378 722 1401 756
rect 1401 722 1412 756
rect 1450 722 1469 756
rect 1469 722 1484 756
rect 1522 722 1537 756
rect 1537 722 1556 756
rect 1594 722 1605 756
rect 1605 722 1628 756
rect 1666 722 1673 756
rect 1673 722 1700 756
rect 1738 722 1741 756
rect 1741 722 1772 756
rect 1810 722 1843 756
rect 1843 722 1844 756
rect 1882 722 1911 756
rect 1911 722 1916 756
rect 1954 722 1979 756
rect 1979 722 1988 756
rect 2026 722 2047 756
rect 2047 722 2060 756
rect 2098 722 2115 756
rect 2115 722 2132 756
rect 2170 722 2183 756
rect 2183 722 2204 756
rect 2242 722 2251 756
rect 2251 722 2276 756
rect 2314 722 2319 756
rect 2319 722 2348 756
rect 2386 722 2387 756
rect 2387 722 2420 756
rect 2458 722 2489 756
rect 2489 722 2492 756
rect 2530 722 2557 756
rect 2557 722 2564 756
rect 2602 722 2625 756
rect 2625 722 2636 756
rect 2674 722 2693 756
rect 2693 722 2708 756
rect 2746 722 2761 756
rect 2761 722 2780 756
rect 2818 722 2829 756
rect 2829 722 2852 756
rect 2890 722 2897 756
rect 2897 722 2924 756
rect 2962 722 2965 756
rect 2965 722 2996 756
rect 3034 722 3067 756
rect 3067 722 3068 756
rect 3106 722 3135 756
rect 3135 722 3140 756
rect 3178 722 3203 756
rect 3203 722 3212 756
rect 3250 722 3271 756
rect 3271 722 3284 756
rect 3322 722 3339 756
rect 3339 722 3356 756
rect 3394 722 3407 756
rect 3407 722 3428 756
rect 3466 722 3475 756
rect 3475 722 3500 756
rect 3538 722 3543 756
rect 3543 722 3572 756
rect 3610 722 3611 756
rect 3611 722 3644 756
rect 3682 722 3713 756
rect 3713 722 3716 756
rect 3754 722 3781 756
rect 3781 722 3788 756
rect 3826 722 3849 756
rect 3849 722 3860 756
rect 3898 722 3917 756
rect 3917 722 3932 756
rect 3970 722 3985 756
rect 3985 722 4004 756
rect 4042 722 4053 756
rect 4053 722 4076 756
rect 4114 722 4121 756
rect 4121 722 4148 756
rect 4186 722 4189 756
rect 4189 722 4220 756
rect 4258 722 4291 756
rect 4291 722 4292 756
rect 4330 722 4359 756
rect 4359 722 4364 756
rect 4402 722 4427 756
rect 4427 722 4436 756
rect 4474 722 4495 756
rect 4495 722 4508 756
rect 4546 722 4563 756
rect 4563 722 4580 756
rect 4618 722 4631 756
rect 4631 722 4652 756
rect 4690 722 4699 756
rect 4699 722 4724 756
rect 4762 722 4767 756
rect 4767 722 4796 756
rect 4834 722 4835 756
rect 4835 722 4868 756
rect 4906 722 4937 756
rect 4937 722 4940 756
rect 4978 722 5005 756
rect 5005 722 5012 756
rect 5050 722 5073 756
rect 5073 722 5084 756
rect 5122 722 5156 756
rect 5339 722 5373 756
rect 5411 722 5422 756
rect 5422 722 5445 756
rect 5483 722 5490 756
rect 5490 722 5517 756
rect 5555 722 5558 756
rect 5558 722 5589 756
rect 5627 722 5660 756
rect 5660 722 5661 756
rect 5699 722 5728 756
rect 5728 722 5733 756
rect 5771 722 5796 756
rect 5796 722 5805 756
rect 5843 722 5864 756
rect 5864 722 5877 756
rect 5915 722 5932 756
rect 5932 722 5949 756
rect 5987 722 6000 756
rect 6000 722 6021 756
rect 6059 722 6068 756
rect 6068 722 6093 756
rect 6131 722 6136 756
rect 6136 722 6165 756
rect 6203 722 6204 756
rect 6204 722 6237 756
rect 6275 722 6306 756
rect 6306 722 6309 756
rect 6347 722 6374 756
rect 6374 722 6381 756
rect 6419 722 6442 756
rect 6442 722 6453 756
rect 6491 722 6510 756
rect 6510 722 6525 756
rect 6563 722 6578 756
rect 6578 722 6597 756
rect 6635 722 6646 756
rect 6646 722 6669 756
rect 6707 722 6714 756
rect 6714 722 6741 756
rect 6779 722 6782 756
rect 6782 722 6813 756
rect 6851 722 6884 756
rect 6884 722 6885 756
rect 6923 722 6952 756
rect 6952 722 6957 756
rect 6995 722 7020 756
rect 7020 722 7029 756
rect 7067 722 7088 756
rect 7088 722 7101 756
rect 7139 722 7156 756
rect 7156 722 7173 756
rect 7211 722 7224 756
rect 7224 722 7245 756
rect 7283 722 7292 756
rect 7292 722 7317 756
rect 7355 722 7360 756
rect 7360 722 7389 756
rect 7427 722 7428 756
rect 7428 722 7461 756
rect 7499 722 7530 756
rect 7530 722 7533 756
rect 7571 722 7598 756
rect 7598 722 7605 756
rect 7643 722 7666 756
rect 7666 722 7677 756
rect 7715 722 7734 756
rect 7734 722 7749 756
rect 7787 722 7802 756
rect 7802 722 7821 756
rect 7859 722 7870 756
rect 7870 722 7893 756
rect 7931 722 7938 756
rect 7938 722 7965 756
rect 8003 722 8006 756
rect 8006 722 8037 756
rect 8075 722 8108 756
rect 8108 722 8109 756
rect 8147 722 8176 756
rect 8176 722 8181 756
rect 8219 722 8244 756
rect 8244 722 8253 756
rect 8291 722 8312 756
rect 8312 722 8325 756
rect 8363 722 8380 756
rect 8380 722 8397 756
rect 8435 722 8448 756
rect 8448 722 8469 756
rect 8507 722 8516 756
rect 8516 722 8541 756
rect 8579 722 8584 756
rect 8584 722 8613 756
rect 8651 722 8652 756
rect 8652 722 8685 756
rect 8723 722 8754 756
rect 8754 722 8757 756
rect 8795 722 8822 756
rect 8822 722 8829 756
rect 8867 722 8890 756
rect 8890 722 8901 756
rect 8939 722 8958 756
rect 8958 722 8973 756
rect 9011 722 9026 756
rect 9026 722 9045 756
rect 9083 722 9094 756
rect 9094 722 9117 756
rect 9155 722 9162 756
rect 9162 722 9189 756
rect 9227 722 9230 756
rect 9230 722 9261 756
rect 9299 722 9332 756
rect 9332 722 9333 756
rect 9371 722 9400 756
rect 9400 722 9405 756
rect 9443 722 9468 756
rect 9468 722 9477 756
rect 9515 722 9549 756
rect 1080 608 1082 642
rect 1082 608 1114 642
rect 1152 608 1184 642
rect 1184 608 1186 642
rect 1532 608 1534 642
rect 1534 608 1566 642
rect 1604 608 1636 642
rect 1636 608 1638 642
rect 1790 608 1792 642
rect 1792 608 1824 642
rect 1862 608 1894 642
rect 1894 608 1896 642
rect 2048 608 2050 642
rect 2050 608 2082 642
rect 2120 608 2152 642
rect 2152 608 2154 642
rect 2306 608 2308 642
rect 2308 608 2340 642
rect 2378 608 2410 642
rect 2410 608 2412 642
rect 2758 608 2760 642
rect 2760 608 2792 642
rect 2830 608 2862 642
rect 2862 608 2864 642
rect 3016 608 3018 642
rect 3018 608 3050 642
rect 3088 608 3120 642
rect 3120 608 3122 642
rect 3274 608 3276 642
rect 3276 608 3308 642
rect 3346 608 3378 642
rect 3378 608 3380 642
rect 3726 608 3728 642
rect 3728 608 3760 642
rect 3798 608 3830 642
rect 3830 608 3832 642
rect 3984 608 3986 642
rect 3986 608 4018 642
rect 4056 608 4088 642
rect 4088 608 4090 642
rect 4242 608 4244 642
rect 4244 608 4276 642
rect 4314 608 4346 642
rect 4346 608 4348 642
rect 4500 608 4502 642
rect 4502 608 4534 642
rect 4572 608 4604 642
rect 4604 608 4606 642
rect 4952 608 4954 642
rect 4954 608 4986 642
rect 5024 608 5056 642
rect 5056 608 5058 642
rect 872 565 906 599
rect 5438 608 5440 642
rect 5440 608 5472 642
rect 5510 608 5542 642
rect 5542 608 5544 642
rect 5889 608 5891 642
rect 5891 608 5923 642
rect 5961 608 5993 642
rect 5993 608 5995 642
rect 6147 608 6149 642
rect 6149 608 6181 642
rect 6219 608 6251 642
rect 6251 608 6253 642
rect 6405 608 6407 642
rect 6407 608 6439 642
rect 6477 608 6509 642
rect 6509 608 6511 642
rect 6663 608 6665 642
rect 6665 608 6697 642
rect 6735 608 6767 642
rect 6767 608 6769 642
rect 7115 608 7117 642
rect 7117 608 7149 642
rect 7187 608 7219 642
rect 7219 608 7221 642
rect 7373 608 7375 642
rect 7375 608 7407 642
rect 7445 608 7477 642
rect 7477 608 7479 642
rect 7631 608 7633 642
rect 7633 608 7665 642
rect 7703 608 7735 642
rect 7735 608 7737 642
rect 8083 608 8085 642
rect 8085 608 8117 642
rect 8155 608 8187 642
rect 8187 608 8189 642
rect 8341 608 8343 642
rect 8343 608 8375 642
rect 8413 608 8445 642
rect 8445 608 8447 642
rect 8599 608 8601 642
rect 8601 608 8633 642
rect 8671 608 8703 642
rect 8703 608 8705 642
rect 8857 608 8859 642
rect 8859 608 8891 642
rect 8929 608 8961 642
rect 8961 608 8963 642
rect 9309 608 9311 642
rect 9311 608 9343 642
rect 9381 608 9413 642
rect 9413 608 9415 642
rect 5231 565 5265 599
rect 9589 565 9623 599
rect 872 509 906 527
rect 872 493 906 509
rect 872 441 906 455
rect 872 421 906 441
rect 872 373 906 383
rect 872 349 906 373
rect 987 512 1021 514
rect 987 480 1021 512
rect 987 410 1021 442
rect 987 408 1021 410
rect 1245 512 1279 514
rect 1245 480 1279 512
rect 1245 410 1279 442
rect 1245 408 1279 410
rect 1439 512 1473 514
rect 1439 480 1473 512
rect 1439 410 1473 442
rect 1439 408 1473 410
rect 1697 512 1731 514
rect 1697 480 1731 512
rect 1697 410 1731 442
rect 1697 408 1731 410
rect 1955 512 1989 514
rect 1955 480 1989 512
rect 1955 410 1989 442
rect 1955 408 1989 410
rect 2213 512 2247 514
rect 2213 480 2247 512
rect 2213 410 2247 442
rect 2213 408 2247 410
rect 2471 512 2505 514
rect 2471 480 2505 512
rect 2471 410 2505 442
rect 2471 408 2505 410
rect 2665 512 2699 514
rect 2665 480 2699 512
rect 2665 410 2699 442
rect 2665 408 2699 410
rect 2923 512 2957 514
rect 2923 480 2957 512
rect 2923 410 2957 442
rect 2923 408 2957 410
rect 3181 512 3215 514
rect 3181 480 3215 512
rect 3181 410 3215 442
rect 3181 408 3215 410
rect 3439 512 3473 514
rect 3439 480 3473 512
rect 3439 410 3473 442
rect 3439 408 3473 410
rect 3633 512 3667 514
rect 3633 480 3667 512
rect 3633 410 3667 442
rect 3633 408 3667 410
rect 3891 512 3925 514
rect 3891 480 3925 512
rect 3891 410 3925 442
rect 3891 408 3925 410
rect 4149 512 4183 514
rect 4149 480 4183 512
rect 4149 410 4183 442
rect 4149 408 4183 410
rect 4407 512 4441 514
rect 4407 480 4441 512
rect 4407 410 4441 442
rect 4407 408 4441 410
rect 4665 512 4699 514
rect 4665 480 4699 512
rect 4665 410 4699 442
rect 4665 408 4699 410
rect 4859 512 4893 514
rect 4859 480 4893 512
rect 4859 410 4893 442
rect 4859 408 4893 410
rect 5117 512 5151 514
rect 5117 480 5151 512
rect 5117 410 5151 442
rect 5117 408 5151 410
rect 5231 509 5265 527
rect 5231 493 5265 509
rect 5231 441 5265 455
rect 5231 421 5265 441
rect 872 305 906 311
rect 872 277 906 305
rect 872 237 906 239
rect 872 205 906 237
rect 872 135 906 167
rect 872 133 906 135
rect 872 67 906 95
rect 872 61 906 67
rect 872 -1 906 23
rect 872 -11 906 -1
rect 5231 373 5265 383
rect 5231 349 5265 373
rect 5345 512 5379 514
rect 5345 480 5379 512
rect 5345 410 5379 442
rect 5345 408 5379 410
rect 5603 512 5637 514
rect 5603 480 5637 512
rect 5603 410 5637 442
rect 5603 408 5637 410
rect 5796 512 5830 514
rect 5796 480 5830 512
rect 5796 410 5830 442
rect 5796 408 5830 410
rect 6054 512 6088 514
rect 6054 480 6088 512
rect 6054 410 6088 442
rect 6054 408 6088 410
rect 6312 512 6346 514
rect 6312 480 6346 512
rect 6312 410 6346 442
rect 6312 408 6346 410
rect 6570 512 6604 514
rect 6570 480 6604 512
rect 6570 410 6604 442
rect 6570 408 6604 410
rect 6828 512 6862 514
rect 6828 480 6862 512
rect 6828 410 6862 442
rect 6828 408 6862 410
rect 7022 512 7056 514
rect 7022 480 7056 512
rect 7022 410 7056 442
rect 7022 408 7056 410
rect 7280 512 7314 514
rect 7280 480 7314 512
rect 7280 410 7314 442
rect 7280 408 7314 410
rect 7538 512 7572 514
rect 7538 480 7572 512
rect 7538 410 7572 442
rect 7538 408 7572 410
rect 7796 512 7830 514
rect 7796 480 7830 512
rect 7796 410 7830 442
rect 7796 408 7830 410
rect 7990 512 8024 514
rect 7990 480 8024 512
rect 7990 410 8024 442
rect 7990 408 8024 410
rect 8248 512 8282 514
rect 8248 480 8282 512
rect 8248 410 8282 442
rect 8248 408 8282 410
rect 8506 512 8540 514
rect 8506 480 8540 512
rect 8506 410 8540 442
rect 8506 408 8540 410
rect 8764 512 8798 514
rect 8764 480 8798 512
rect 8764 410 8798 442
rect 8764 408 8798 410
rect 9022 512 9056 514
rect 9022 480 9056 512
rect 9022 410 9056 442
rect 9022 408 9056 410
rect 9216 512 9250 514
rect 9216 480 9250 512
rect 9216 410 9250 442
rect 9216 408 9250 410
rect 9474 512 9508 514
rect 9474 480 9508 512
rect 9474 410 9508 442
rect 9474 408 9508 410
rect 9589 509 9623 527
rect 9589 493 9623 509
rect 9589 441 9623 455
rect 9589 421 9623 441
rect 9589 373 9623 383
rect 5231 305 5265 311
rect 5231 277 5265 305
rect 5231 237 5265 239
rect 5231 205 5265 237
rect 5231 135 5265 167
rect 5231 133 5265 135
rect 5231 67 5265 95
rect 5231 61 5265 67
rect 5231 -1 5265 23
rect 5231 -11 5265 -1
rect 9589 349 9623 373
rect 9589 305 9623 311
rect 9589 277 9623 305
rect 9589 237 9623 239
rect 9589 205 9623 237
rect 9589 135 9623 167
rect 9589 133 9623 135
rect 9589 67 9623 95
rect 9589 61 9623 67
rect 9589 -1 9623 23
rect 9589 -11 9623 -1
rect 872 -69 906 -49
rect 5231 -69 5265 -49
rect 9589 -69 9623 -49
rect 872 -83 906 -69
rect 872 -137 906 -121
rect 872 -155 906 -137
rect 872 -205 906 -193
rect 872 -227 906 -205
rect 872 -273 906 -265
rect 872 -299 906 -273
rect 872 -341 906 -337
rect 872 -371 906 -341
rect 5231 -83 5265 -69
rect 5231 -137 5265 -121
rect 5231 -155 5265 -137
rect 5231 -205 5265 -193
rect 5231 -227 5265 -205
rect 5231 -273 5265 -265
rect 5231 -299 5265 -273
rect 5231 -341 5265 -337
rect 5231 -371 5265 -341
rect 872 -443 906 -409
rect 872 -511 906 -481
rect 872 -515 906 -511
rect 872 -579 906 -553
rect 872 -587 906 -579
rect 987 -432 1021 -430
rect 987 -464 1021 -432
rect 987 -534 1021 -502
rect 987 -536 1021 -534
rect 1245 -432 1279 -430
rect 1245 -464 1279 -432
rect 1245 -534 1279 -502
rect 1245 -536 1279 -534
rect 1439 -432 1473 -430
rect 1439 -464 1473 -432
rect 1439 -534 1473 -502
rect 1439 -536 1473 -534
rect 1697 -432 1731 -430
rect 1697 -464 1731 -432
rect 1697 -534 1731 -502
rect 1697 -536 1731 -534
rect 1955 -432 1989 -430
rect 1955 -464 1989 -432
rect 1955 -534 1989 -502
rect 1955 -536 1989 -534
rect 2213 -432 2247 -430
rect 2213 -464 2247 -432
rect 2213 -534 2247 -502
rect 2213 -536 2247 -534
rect 2471 -432 2505 -430
rect 2471 -464 2505 -432
rect 2471 -534 2505 -502
rect 2471 -536 2505 -534
rect 2665 -432 2699 -430
rect 2665 -464 2699 -432
rect 2665 -534 2699 -502
rect 2665 -536 2699 -534
rect 2923 -432 2957 -430
rect 2923 -464 2957 -432
rect 2923 -534 2957 -502
rect 2923 -536 2957 -534
rect 3181 -432 3215 -430
rect 3181 -464 3215 -432
rect 3181 -534 3215 -502
rect 3181 -536 3215 -534
rect 3439 -432 3473 -430
rect 3439 -464 3473 -432
rect 3439 -534 3473 -502
rect 3439 -536 3473 -534
rect 3633 -432 3667 -430
rect 3633 -464 3667 -432
rect 3633 -534 3667 -502
rect 3633 -536 3667 -534
rect 3891 -432 3925 -430
rect 3891 -464 3925 -432
rect 3891 -534 3925 -502
rect 3891 -536 3925 -534
rect 4149 -432 4183 -430
rect 4149 -464 4183 -432
rect 4149 -534 4183 -502
rect 4149 -536 4183 -534
rect 4407 -432 4441 -430
rect 4407 -464 4441 -432
rect 4407 -534 4441 -502
rect 4407 -536 4441 -534
rect 4665 -432 4699 -430
rect 4665 -464 4699 -432
rect 4665 -534 4699 -502
rect 4665 -536 4699 -534
rect 4859 -432 4893 -430
rect 4859 -464 4893 -432
rect 4859 -534 4893 -502
rect 4859 -536 4893 -534
rect 5117 -432 5151 -430
rect 5117 -464 5151 -432
rect 5117 -534 5151 -502
rect 5117 -536 5151 -534
rect 9589 -83 9623 -69
rect 9589 -137 9623 -121
rect 9589 -155 9623 -137
rect 9589 -205 9623 -193
rect 9589 -227 9623 -205
rect 9589 -273 9623 -265
rect 9589 -299 9623 -273
rect 9589 -341 9623 -337
rect 9589 -371 9623 -341
rect 5231 -443 5265 -409
rect 5231 -511 5265 -481
rect 5231 -515 5265 -511
rect 5231 -579 5265 -553
rect 5231 -587 5265 -579
rect 5345 -432 5379 -430
rect 5345 -464 5379 -432
rect 5345 -534 5379 -502
rect 5345 -536 5379 -534
rect 5603 -432 5637 -430
rect 5603 -464 5637 -432
rect 5603 -534 5637 -502
rect 5603 -536 5637 -534
rect 5796 -432 5830 -430
rect 5796 -464 5830 -432
rect 5796 -534 5830 -502
rect 5796 -536 5830 -534
rect 6054 -432 6088 -430
rect 6054 -464 6088 -432
rect 6054 -534 6088 -502
rect 6054 -536 6088 -534
rect 6312 -432 6346 -430
rect 6312 -464 6346 -432
rect 6312 -534 6346 -502
rect 6312 -536 6346 -534
rect 6570 -432 6604 -430
rect 6570 -464 6604 -432
rect 6570 -534 6604 -502
rect 6570 -536 6604 -534
rect 6828 -432 6862 -430
rect 6828 -464 6862 -432
rect 6828 -534 6862 -502
rect 6828 -536 6862 -534
rect 7022 -432 7056 -430
rect 7022 -464 7056 -432
rect 7022 -534 7056 -502
rect 7022 -536 7056 -534
rect 7280 -432 7314 -430
rect 7280 -464 7314 -432
rect 7280 -534 7314 -502
rect 7280 -536 7314 -534
rect 7538 -432 7572 -430
rect 7538 -464 7572 -432
rect 7538 -534 7572 -502
rect 7538 -536 7572 -534
rect 7796 -432 7830 -430
rect 7796 -464 7830 -432
rect 7796 -534 7830 -502
rect 7796 -536 7830 -534
rect 7990 -432 8024 -430
rect 7990 -464 8024 -432
rect 7990 -534 8024 -502
rect 7990 -536 8024 -534
rect 8248 -432 8282 -430
rect 8248 -464 8282 -432
rect 8248 -534 8282 -502
rect 8248 -536 8282 -534
rect 8506 -432 8540 -430
rect 8506 -464 8540 -432
rect 8506 -534 8540 -502
rect 8506 -536 8540 -534
rect 8764 -432 8798 -430
rect 8764 -464 8798 -432
rect 8764 -534 8798 -502
rect 8764 -536 8798 -534
rect 9022 -432 9056 -430
rect 9022 -464 9056 -432
rect 9022 -534 9056 -502
rect 9022 -536 9056 -534
rect 9216 -432 9250 -430
rect 9216 -464 9250 -432
rect 9216 -534 9250 -502
rect 9216 -536 9250 -534
rect 9474 -432 9508 -430
rect 9474 -464 9508 -432
rect 9474 -534 9508 -502
rect 9474 -536 9508 -534
rect 9589 -443 9623 -409
rect 9589 -511 9623 -481
rect 9589 -515 9623 -511
rect 9589 -579 9623 -553
rect 9589 -587 9623 -579
rect 872 -647 906 -625
rect 872 -659 906 -647
rect 1080 -664 1082 -630
rect 1082 -664 1114 -630
rect 1152 -664 1184 -630
rect 1184 -664 1186 -630
rect 1532 -664 1534 -630
rect 1534 -664 1566 -630
rect 1604 -664 1636 -630
rect 1636 -664 1638 -630
rect 1790 -664 1792 -630
rect 1792 -664 1824 -630
rect 1862 -664 1894 -630
rect 1894 -664 1896 -630
rect 2048 -664 2050 -630
rect 2050 -664 2082 -630
rect 2120 -664 2152 -630
rect 2152 -664 2154 -630
rect 2306 -664 2308 -630
rect 2308 -664 2340 -630
rect 2378 -664 2410 -630
rect 2410 -664 2412 -630
rect 2758 -664 2760 -630
rect 2760 -664 2792 -630
rect 2830 -664 2862 -630
rect 2862 -664 2864 -630
rect 3016 -664 3018 -630
rect 3018 -664 3050 -630
rect 3088 -664 3120 -630
rect 3120 -664 3122 -630
rect 3274 -664 3276 -630
rect 3276 -664 3308 -630
rect 3346 -664 3378 -630
rect 3378 -664 3380 -630
rect 3726 -664 3728 -630
rect 3728 -664 3760 -630
rect 3798 -664 3830 -630
rect 3830 -664 3832 -630
rect 3984 -664 3986 -630
rect 3986 -664 4018 -630
rect 4056 -664 4088 -630
rect 4088 -664 4090 -630
rect 4242 -664 4244 -630
rect 4244 -664 4276 -630
rect 4314 -664 4346 -630
rect 4346 -664 4348 -630
rect 4500 -664 4502 -630
rect 4502 -664 4534 -630
rect 4572 -664 4604 -630
rect 4604 -664 4606 -630
rect 4952 -664 4954 -630
rect 4954 -664 4986 -630
rect 5024 -664 5056 -630
rect 5056 -664 5058 -630
rect 5231 -647 5265 -625
rect 5231 -659 5265 -647
rect 872 -715 906 -697
rect 872 -731 906 -715
rect 872 -783 906 -769
rect 872 -803 906 -783
rect 872 -851 906 -841
rect 872 -875 906 -851
rect 872 -919 906 -913
rect 872 -947 906 -919
rect 872 -987 906 -985
rect 872 -1019 906 -987
rect 5438 -664 5440 -630
rect 5440 -664 5472 -630
rect 5510 -664 5542 -630
rect 5542 -664 5544 -630
rect 5889 -664 5891 -630
rect 5891 -664 5923 -630
rect 5961 -664 5993 -630
rect 5993 -664 5995 -630
rect 6147 -664 6149 -630
rect 6149 -664 6181 -630
rect 6219 -664 6251 -630
rect 6251 -664 6253 -630
rect 6405 -664 6407 -630
rect 6407 -664 6439 -630
rect 6477 -664 6509 -630
rect 6509 -664 6511 -630
rect 6663 -664 6665 -630
rect 6665 -664 6697 -630
rect 6735 -664 6767 -630
rect 6767 -664 6769 -630
rect 7115 -664 7117 -630
rect 7117 -664 7149 -630
rect 7187 -664 7219 -630
rect 7219 -664 7221 -630
rect 7373 -664 7375 -630
rect 7375 -664 7407 -630
rect 7445 -664 7477 -630
rect 7477 -664 7479 -630
rect 7631 -664 7633 -630
rect 7633 -664 7665 -630
rect 7703 -664 7735 -630
rect 7735 -664 7737 -630
rect 8083 -664 8085 -630
rect 8085 -664 8117 -630
rect 8155 -664 8187 -630
rect 8187 -664 8189 -630
rect 8341 -664 8343 -630
rect 8343 -664 8375 -630
rect 8413 -664 8445 -630
rect 8445 -664 8447 -630
rect 8599 -664 8601 -630
rect 8601 -664 8633 -630
rect 8671 -664 8703 -630
rect 8703 -664 8705 -630
rect 8857 -664 8859 -630
rect 8859 -664 8891 -630
rect 8929 -664 8961 -630
rect 8961 -664 8963 -630
rect 9309 -664 9311 -630
rect 9311 -664 9343 -630
rect 9381 -664 9413 -630
rect 9413 -664 9415 -630
rect 9589 -647 9623 -625
rect 9589 -659 9623 -647
rect 5231 -715 5265 -697
rect 5231 -731 5265 -715
rect 5231 -783 5265 -769
rect 5231 -803 5265 -783
rect 5231 -851 5265 -841
rect 5231 -875 5265 -851
rect 5231 -919 5265 -913
rect 5231 -947 5265 -919
rect 1080 -1027 1082 -993
rect 1082 -1027 1114 -993
rect 1152 -1027 1184 -993
rect 1184 -1027 1186 -993
rect 1532 -1027 1534 -993
rect 1534 -1027 1566 -993
rect 1604 -1027 1636 -993
rect 1636 -1027 1638 -993
rect 1790 -1027 1792 -993
rect 1792 -1027 1824 -993
rect 1862 -1027 1894 -993
rect 1894 -1027 1896 -993
rect 2048 -1027 2050 -993
rect 2050 -1027 2082 -993
rect 2120 -1027 2152 -993
rect 2152 -1027 2154 -993
rect 2306 -1027 2308 -993
rect 2308 -1027 2340 -993
rect 2378 -1027 2410 -993
rect 2410 -1027 2412 -993
rect 2758 -1027 2760 -993
rect 2760 -1027 2792 -993
rect 2830 -1027 2862 -993
rect 2862 -1027 2864 -993
rect 3016 -1027 3018 -993
rect 3018 -1027 3050 -993
rect 3088 -1027 3120 -993
rect 3120 -1027 3122 -993
rect 3274 -1027 3276 -993
rect 3276 -1027 3308 -993
rect 3346 -1027 3378 -993
rect 3378 -1027 3380 -993
rect 3726 -1027 3728 -993
rect 3728 -1027 3760 -993
rect 3798 -1027 3830 -993
rect 3830 -1027 3832 -993
rect 3984 -1027 3986 -993
rect 3986 -1027 4018 -993
rect 4056 -1027 4088 -993
rect 4088 -1027 4090 -993
rect 4242 -1027 4244 -993
rect 4244 -1027 4276 -993
rect 4314 -1027 4346 -993
rect 4346 -1027 4348 -993
rect 4500 -1027 4502 -993
rect 4502 -1027 4534 -993
rect 4572 -1027 4604 -993
rect 4604 -1027 4606 -993
rect 4952 -1027 4954 -993
rect 4954 -1027 4986 -993
rect 5024 -1027 5056 -993
rect 5056 -1027 5058 -993
rect 5231 -987 5265 -985
rect 5231 -1019 5265 -987
rect 9589 -715 9623 -697
rect 9589 -731 9623 -715
rect 9589 -783 9623 -769
rect 9589 -803 9623 -783
rect 9589 -851 9623 -841
rect 9589 -875 9623 -851
rect 9589 -919 9623 -913
rect 9589 -947 9623 -919
rect 9589 -987 9623 -985
rect 872 -1089 906 -1057
rect 5438 -1027 5440 -993
rect 5440 -1027 5472 -993
rect 5510 -1027 5542 -993
rect 5542 -1027 5544 -993
rect 5889 -1027 5891 -993
rect 5891 -1027 5923 -993
rect 5961 -1027 5993 -993
rect 5993 -1027 5995 -993
rect 6147 -1027 6149 -993
rect 6149 -1027 6181 -993
rect 6219 -1027 6251 -993
rect 6251 -1027 6253 -993
rect 6405 -1027 6407 -993
rect 6407 -1027 6439 -993
rect 6477 -1027 6509 -993
rect 6509 -1027 6511 -993
rect 6663 -1027 6665 -993
rect 6665 -1027 6697 -993
rect 6735 -1027 6767 -993
rect 6767 -1027 6769 -993
rect 7115 -1027 7117 -993
rect 7117 -1027 7149 -993
rect 7187 -1027 7219 -993
rect 7219 -1027 7221 -993
rect 7373 -1027 7375 -993
rect 7375 -1027 7407 -993
rect 7445 -1027 7477 -993
rect 7477 -1027 7479 -993
rect 7631 -1027 7633 -993
rect 7633 -1027 7665 -993
rect 7703 -1027 7735 -993
rect 7735 -1027 7737 -993
rect 8083 -1027 8085 -993
rect 8085 -1027 8117 -993
rect 8155 -1027 8187 -993
rect 8187 -1027 8189 -993
rect 8341 -1027 8343 -993
rect 8343 -1027 8375 -993
rect 8413 -1027 8445 -993
rect 8445 -1027 8447 -993
rect 8599 -1027 8601 -993
rect 8601 -1027 8633 -993
rect 8671 -1027 8703 -993
rect 8703 -1027 8705 -993
rect 8857 -1027 8859 -993
rect 8859 -1027 8891 -993
rect 8929 -1027 8961 -993
rect 8961 -1027 8963 -993
rect 9309 -1027 9311 -993
rect 9311 -1027 9343 -993
rect 9381 -1027 9413 -993
rect 9413 -1027 9415 -993
rect 9589 -1019 9623 -987
rect 872 -1091 906 -1089
rect 872 -1157 906 -1129
rect 872 -1163 906 -1157
rect 872 -1225 906 -1201
rect 872 -1235 906 -1225
rect 872 -1293 906 -1273
rect 987 -1123 1021 -1121
rect 987 -1155 1021 -1123
rect 987 -1225 1021 -1193
rect 987 -1227 1021 -1225
rect 1245 -1123 1279 -1121
rect 1245 -1155 1279 -1123
rect 1245 -1225 1279 -1193
rect 1245 -1227 1279 -1225
rect 1439 -1123 1473 -1121
rect 1439 -1155 1473 -1123
rect 1439 -1225 1473 -1193
rect 1439 -1227 1473 -1225
rect 1697 -1123 1731 -1121
rect 1697 -1155 1731 -1123
rect 1697 -1225 1731 -1193
rect 1697 -1227 1731 -1225
rect 1955 -1123 1989 -1121
rect 1955 -1155 1989 -1123
rect 1955 -1225 1989 -1193
rect 1955 -1227 1989 -1225
rect 2213 -1123 2247 -1121
rect 2213 -1155 2247 -1123
rect 2213 -1225 2247 -1193
rect 2213 -1227 2247 -1225
rect 2471 -1123 2505 -1121
rect 2471 -1155 2505 -1123
rect 2471 -1225 2505 -1193
rect 2471 -1227 2505 -1225
rect 2665 -1123 2699 -1121
rect 2665 -1155 2699 -1123
rect 2665 -1225 2699 -1193
rect 2665 -1227 2699 -1225
rect 2923 -1123 2957 -1121
rect 2923 -1155 2957 -1123
rect 2923 -1225 2957 -1193
rect 2923 -1227 2957 -1225
rect 3181 -1123 3215 -1121
rect 3181 -1155 3215 -1123
rect 3181 -1225 3215 -1193
rect 3181 -1227 3215 -1225
rect 3439 -1123 3473 -1121
rect 3439 -1155 3473 -1123
rect 3439 -1225 3473 -1193
rect 3439 -1227 3473 -1225
rect 3633 -1123 3667 -1121
rect 3633 -1155 3667 -1123
rect 3633 -1225 3667 -1193
rect 3633 -1227 3667 -1225
rect 3891 -1123 3925 -1121
rect 3891 -1155 3925 -1123
rect 3891 -1225 3925 -1193
rect 3891 -1227 3925 -1225
rect 4149 -1123 4183 -1121
rect 4149 -1155 4183 -1123
rect 4149 -1225 4183 -1193
rect 4149 -1227 4183 -1225
rect 4407 -1123 4441 -1121
rect 4407 -1155 4441 -1123
rect 4407 -1225 4441 -1193
rect 4407 -1227 4441 -1225
rect 4665 -1123 4699 -1121
rect 4665 -1155 4699 -1123
rect 4665 -1225 4699 -1193
rect 4665 -1227 4699 -1225
rect 4859 -1123 4893 -1121
rect 4859 -1155 4893 -1123
rect 4859 -1225 4893 -1193
rect 4859 -1227 4893 -1225
rect 5117 -1123 5151 -1121
rect 5117 -1155 5151 -1123
rect 5117 -1225 5151 -1193
rect 5117 -1227 5151 -1225
rect 5231 -1089 5265 -1057
rect 5231 -1091 5265 -1089
rect 5231 -1157 5265 -1129
rect 5231 -1163 5265 -1157
rect 5231 -1225 5265 -1201
rect 5231 -1235 5265 -1225
rect 872 -1307 906 -1293
rect 872 -1361 906 -1345
rect 872 -1379 906 -1361
rect 872 -1429 906 -1417
rect 872 -1451 906 -1429
rect 872 -1497 906 -1489
rect 872 -1523 906 -1497
rect 872 -1595 906 -1561
rect 5231 -1293 5265 -1273
rect 5345 -1123 5379 -1121
rect 5345 -1155 5379 -1123
rect 5345 -1225 5379 -1193
rect 5345 -1227 5379 -1225
rect 5603 -1123 5637 -1121
rect 5603 -1155 5637 -1123
rect 5603 -1225 5637 -1193
rect 5603 -1227 5637 -1225
rect 5796 -1123 5830 -1121
rect 5796 -1155 5830 -1123
rect 5796 -1225 5830 -1193
rect 5796 -1227 5830 -1225
rect 6054 -1123 6088 -1121
rect 6054 -1155 6088 -1123
rect 6054 -1225 6088 -1193
rect 6054 -1227 6088 -1225
rect 6312 -1123 6346 -1121
rect 6312 -1155 6346 -1123
rect 6312 -1225 6346 -1193
rect 6312 -1227 6346 -1225
rect 6570 -1123 6604 -1121
rect 6570 -1155 6604 -1123
rect 6570 -1225 6604 -1193
rect 6570 -1227 6604 -1225
rect 6828 -1123 6862 -1121
rect 6828 -1155 6862 -1123
rect 6828 -1225 6862 -1193
rect 6828 -1227 6862 -1225
rect 7022 -1123 7056 -1121
rect 7022 -1155 7056 -1123
rect 7022 -1225 7056 -1193
rect 7022 -1227 7056 -1225
rect 7280 -1123 7314 -1121
rect 7280 -1155 7314 -1123
rect 7280 -1225 7314 -1193
rect 7280 -1227 7314 -1225
rect 7538 -1123 7572 -1121
rect 7538 -1155 7572 -1123
rect 7538 -1225 7572 -1193
rect 7538 -1227 7572 -1225
rect 7796 -1123 7830 -1121
rect 7796 -1155 7830 -1123
rect 7796 -1225 7830 -1193
rect 7796 -1227 7830 -1225
rect 7990 -1123 8024 -1121
rect 7990 -1155 8024 -1123
rect 7990 -1225 8024 -1193
rect 7990 -1227 8024 -1225
rect 8248 -1123 8282 -1121
rect 8248 -1155 8282 -1123
rect 8248 -1225 8282 -1193
rect 8248 -1227 8282 -1225
rect 8506 -1123 8540 -1121
rect 8506 -1155 8540 -1123
rect 8506 -1225 8540 -1193
rect 8506 -1227 8540 -1225
rect 8764 -1123 8798 -1121
rect 8764 -1155 8798 -1123
rect 8764 -1225 8798 -1193
rect 8764 -1227 8798 -1225
rect 9022 -1123 9056 -1121
rect 9022 -1155 9056 -1123
rect 9022 -1225 9056 -1193
rect 9022 -1227 9056 -1225
rect 9216 -1123 9250 -1121
rect 9216 -1155 9250 -1123
rect 9216 -1225 9250 -1193
rect 9216 -1227 9250 -1225
rect 9474 -1123 9508 -1121
rect 9474 -1155 9508 -1123
rect 9474 -1225 9508 -1193
rect 9474 -1227 9508 -1225
rect 9589 -1089 9623 -1057
rect 9589 -1091 9623 -1089
rect 9589 -1157 9623 -1129
rect 9589 -1163 9623 -1157
rect 9589 -1225 9623 -1201
rect 9589 -1235 9623 -1225
rect 5231 -1307 5265 -1293
rect 5231 -1361 5265 -1345
rect 5231 -1379 5265 -1361
rect 5231 -1429 5265 -1417
rect 5231 -1451 5265 -1429
rect 5231 -1497 5265 -1489
rect 5231 -1523 5265 -1497
rect 5231 -1595 5265 -1561
rect 9589 -1293 9623 -1273
rect 9589 -1307 9623 -1293
rect 9589 -1361 9623 -1345
rect 9589 -1379 9623 -1361
rect 9589 -1429 9623 -1417
rect 9589 -1451 9623 -1429
rect 9589 -1497 9623 -1489
rect 9589 -1523 9623 -1497
rect 9589 -1595 9623 -1561
rect 872 -1667 906 -1633
rect 5231 -1667 5265 -1633
rect 9589 -1667 9623 -1633
rect 872 -1739 906 -1705
rect 872 -1803 906 -1777
rect 872 -1811 906 -1803
rect 872 -1871 906 -1849
rect 872 -1883 906 -1871
rect 872 -1939 906 -1921
rect 872 -1955 906 -1939
rect 872 -2007 906 -1993
rect 872 -2027 906 -2007
rect 5231 -1739 5265 -1705
rect 5231 -1803 5265 -1777
rect 5231 -1811 5265 -1803
rect 5231 -1871 5265 -1849
rect 5231 -1883 5265 -1871
rect 5231 -1939 5265 -1921
rect 5231 -1955 5265 -1939
rect 872 -2075 906 -2065
rect 872 -2099 906 -2075
rect 872 -2143 906 -2137
rect 872 -2171 906 -2143
rect 872 -2211 906 -2209
rect 872 -2243 906 -2211
rect 987 -2079 1021 -2077
rect 987 -2111 1021 -2079
rect 987 -2181 1021 -2149
rect 987 -2183 1021 -2181
rect 1245 -2079 1279 -2077
rect 1245 -2111 1279 -2079
rect 1245 -2181 1279 -2149
rect 1245 -2183 1279 -2181
rect 1439 -2079 1473 -2077
rect 1439 -2111 1473 -2079
rect 1439 -2181 1473 -2149
rect 1439 -2183 1473 -2181
rect 1697 -2079 1731 -2077
rect 1697 -2111 1731 -2079
rect 1697 -2181 1731 -2149
rect 1697 -2183 1731 -2181
rect 1955 -2079 1989 -2077
rect 1955 -2111 1989 -2079
rect 1955 -2181 1989 -2149
rect 1955 -2183 1989 -2181
rect 2213 -2079 2247 -2077
rect 2213 -2111 2247 -2079
rect 2213 -2181 2247 -2149
rect 2213 -2183 2247 -2181
rect 2471 -2079 2505 -2077
rect 2471 -2111 2505 -2079
rect 2471 -2181 2505 -2149
rect 2471 -2183 2505 -2181
rect 2665 -2079 2699 -2077
rect 2665 -2111 2699 -2079
rect 2665 -2181 2699 -2149
rect 2665 -2183 2699 -2181
rect 2923 -2079 2957 -2077
rect 2923 -2111 2957 -2079
rect 2923 -2181 2957 -2149
rect 2923 -2183 2957 -2181
rect 3181 -2079 3215 -2077
rect 3181 -2111 3215 -2079
rect 3181 -2181 3215 -2149
rect 3181 -2183 3215 -2181
rect 3439 -2079 3473 -2077
rect 3439 -2111 3473 -2079
rect 3439 -2181 3473 -2149
rect 3439 -2183 3473 -2181
rect 3633 -2079 3667 -2077
rect 3633 -2111 3667 -2079
rect 3633 -2181 3667 -2149
rect 3633 -2183 3667 -2181
rect 3891 -2079 3925 -2077
rect 3891 -2111 3925 -2079
rect 3891 -2181 3925 -2149
rect 3891 -2183 3925 -2181
rect 4149 -2079 4183 -2077
rect 4149 -2111 4183 -2079
rect 4149 -2181 4183 -2149
rect 4149 -2183 4183 -2181
rect 4407 -2079 4441 -2077
rect 4407 -2111 4441 -2079
rect 4407 -2181 4441 -2149
rect 4407 -2183 4441 -2181
rect 4665 -2079 4699 -2077
rect 4665 -2111 4699 -2079
rect 4665 -2181 4699 -2149
rect 4665 -2183 4699 -2181
rect 4859 -2079 4893 -2077
rect 4859 -2111 4893 -2079
rect 4859 -2181 4893 -2149
rect 4859 -2183 4893 -2181
rect 5117 -2079 5151 -2077
rect 5117 -2111 5151 -2079
rect 5117 -2181 5151 -2149
rect 5117 -2183 5151 -2181
rect 5231 -2007 5265 -1993
rect 5231 -2027 5265 -2007
rect 9589 -1739 9623 -1705
rect 9589 -1803 9623 -1777
rect 9589 -1811 9623 -1803
rect 9589 -1871 9623 -1849
rect 9589 -1883 9623 -1871
rect 9589 -1939 9623 -1921
rect 9589 -1955 9623 -1939
rect 9589 -2007 9623 -1993
rect 5231 -2075 5265 -2065
rect 5231 -2099 5265 -2075
rect 5231 -2143 5265 -2137
rect 5231 -2171 5265 -2143
rect 5231 -2211 5265 -2209
rect 5231 -2243 5265 -2211
rect 5345 -2079 5379 -2077
rect 5345 -2111 5379 -2079
rect 5345 -2181 5379 -2149
rect 5345 -2183 5379 -2181
rect 5603 -2079 5637 -2077
rect 5603 -2111 5637 -2079
rect 5603 -2181 5637 -2149
rect 5603 -2183 5637 -2181
rect 5796 -2079 5830 -2077
rect 5796 -2111 5830 -2079
rect 5796 -2181 5830 -2149
rect 5796 -2183 5830 -2181
rect 6054 -2079 6088 -2077
rect 6054 -2111 6088 -2079
rect 6054 -2181 6088 -2149
rect 6054 -2183 6088 -2181
rect 6312 -2079 6346 -2077
rect 6312 -2111 6346 -2079
rect 6312 -2181 6346 -2149
rect 6312 -2183 6346 -2181
rect 6570 -2079 6604 -2077
rect 6570 -2111 6604 -2079
rect 6570 -2181 6604 -2149
rect 6570 -2183 6604 -2181
rect 6828 -2079 6862 -2077
rect 6828 -2111 6862 -2079
rect 6828 -2181 6862 -2149
rect 6828 -2183 6862 -2181
rect 7022 -2079 7056 -2077
rect 7022 -2111 7056 -2079
rect 7022 -2181 7056 -2149
rect 7022 -2183 7056 -2181
rect 7280 -2079 7314 -2077
rect 7280 -2111 7314 -2079
rect 7280 -2181 7314 -2149
rect 7280 -2183 7314 -2181
rect 7538 -2079 7572 -2077
rect 7538 -2111 7572 -2079
rect 7538 -2181 7572 -2149
rect 7538 -2183 7572 -2181
rect 7796 -2079 7830 -2077
rect 7796 -2111 7830 -2079
rect 7796 -2181 7830 -2149
rect 7796 -2183 7830 -2181
rect 7990 -2079 8024 -2077
rect 7990 -2111 8024 -2079
rect 7990 -2181 8024 -2149
rect 7990 -2183 8024 -2181
rect 8248 -2079 8282 -2077
rect 8248 -2111 8282 -2079
rect 8248 -2181 8282 -2149
rect 8248 -2183 8282 -2181
rect 8506 -2079 8540 -2077
rect 8506 -2111 8540 -2079
rect 8506 -2181 8540 -2149
rect 8506 -2183 8540 -2181
rect 8764 -2079 8798 -2077
rect 8764 -2111 8798 -2079
rect 8764 -2181 8798 -2149
rect 8764 -2183 8798 -2181
rect 9022 -2079 9056 -2077
rect 9022 -2111 9056 -2079
rect 9022 -2181 9056 -2149
rect 9022 -2183 9056 -2181
rect 9216 -2079 9250 -2077
rect 9216 -2111 9250 -2079
rect 9216 -2181 9250 -2149
rect 9216 -2183 9250 -2181
rect 9474 -2079 9508 -2077
rect 9474 -2111 9508 -2079
rect 9474 -2181 9508 -2149
rect 9474 -2183 9508 -2181
rect 9589 -2027 9623 -2007
rect 9589 -2075 9623 -2065
rect 9589 -2099 9623 -2075
rect 9589 -2143 9623 -2137
rect 9589 -2171 9623 -2143
rect 9589 -2211 9623 -2209
rect 872 -2313 906 -2281
rect 1080 -2311 1082 -2277
rect 1082 -2311 1114 -2277
rect 1152 -2311 1184 -2277
rect 1184 -2311 1186 -2277
rect 1532 -2311 1534 -2277
rect 1534 -2311 1566 -2277
rect 1604 -2311 1636 -2277
rect 1636 -2311 1638 -2277
rect 1790 -2311 1792 -2277
rect 1792 -2311 1824 -2277
rect 1862 -2311 1894 -2277
rect 1894 -2311 1896 -2277
rect 2048 -2311 2050 -2277
rect 2050 -2311 2082 -2277
rect 2120 -2311 2152 -2277
rect 2152 -2311 2154 -2277
rect 2306 -2311 2308 -2277
rect 2308 -2311 2340 -2277
rect 2378 -2311 2410 -2277
rect 2410 -2311 2412 -2277
rect 2758 -2311 2760 -2277
rect 2760 -2311 2792 -2277
rect 2830 -2311 2862 -2277
rect 2862 -2311 2864 -2277
rect 3016 -2311 3018 -2277
rect 3018 -2311 3050 -2277
rect 3088 -2311 3120 -2277
rect 3120 -2311 3122 -2277
rect 3274 -2311 3276 -2277
rect 3276 -2311 3308 -2277
rect 3346 -2311 3378 -2277
rect 3378 -2311 3380 -2277
rect 3726 -2311 3728 -2277
rect 3728 -2311 3760 -2277
rect 3798 -2311 3830 -2277
rect 3830 -2311 3832 -2277
rect 3984 -2311 3986 -2277
rect 3986 -2311 4018 -2277
rect 4056 -2311 4088 -2277
rect 4088 -2311 4090 -2277
rect 4242 -2311 4244 -2277
rect 4244 -2311 4276 -2277
rect 4314 -2311 4346 -2277
rect 4346 -2311 4348 -2277
rect 4500 -2311 4502 -2277
rect 4502 -2311 4534 -2277
rect 4572 -2311 4604 -2277
rect 4604 -2311 4606 -2277
rect 4952 -2311 4954 -2277
rect 4954 -2311 4986 -2277
rect 5024 -2311 5056 -2277
rect 5056 -2311 5058 -2277
rect 9589 -2243 9623 -2211
rect 872 -2315 906 -2313
rect 872 -2381 906 -2353
rect 872 -2387 906 -2381
rect 872 -2449 906 -2425
rect 872 -2459 906 -2449
rect 872 -2517 906 -2497
rect 872 -2531 906 -2517
rect 872 -2585 906 -2569
rect 872 -2603 906 -2585
rect 5231 -2313 5265 -2281
rect 5438 -2311 5440 -2277
rect 5440 -2311 5472 -2277
rect 5510 -2311 5542 -2277
rect 5542 -2311 5544 -2277
rect 5889 -2311 5891 -2277
rect 5891 -2311 5923 -2277
rect 5961 -2311 5993 -2277
rect 5993 -2311 5995 -2277
rect 6147 -2311 6149 -2277
rect 6149 -2311 6181 -2277
rect 6219 -2311 6251 -2277
rect 6251 -2311 6253 -2277
rect 6405 -2311 6407 -2277
rect 6407 -2311 6439 -2277
rect 6477 -2311 6509 -2277
rect 6509 -2311 6511 -2277
rect 6663 -2311 6665 -2277
rect 6665 -2311 6697 -2277
rect 6735 -2311 6767 -2277
rect 6767 -2311 6769 -2277
rect 7115 -2311 7117 -2277
rect 7117 -2311 7149 -2277
rect 7187 -2311 7219 -2277
rect 7219 -2311 7221 -2277
rect 7373 -2311 7375 -2277
rect 7375 -2311 7407 -2277
rect 7445 -2311 7477 -2277
rect 7477 -2311 7479 -2277
rect 7631 -2311 7633 -2277
rect 7633 -2311 7665 -2277
rect 7703 -2311 7735 -2277
rect 7735 -2311 7737 -2277
rect 8083 -2311 8085 -2277
rect 8085 -2311 8117 -2277
rect 8155 -2311 8187 -2277
rect 8187 -2311 8189 -2277
rect 8341 -2311 8343 -2277
rect 8343 -2311 8375 -2277
rect 8413 -2311 8445 -2277
rect 8445 -2311 8447 -2277
rect 8599 -2311 8601 -2277
rect 8601 -2311 8633 -2277
rect 8671 -2311 8703 -2277
rect 8703 -2311 8705 -2277
rect 8857 -2311 8859 -2277
rect 8859 -2311 8891 -2277
rect 8929 -2311 8961 -2277
rect 8961 -2311 8963 -2277
rect 9309 -2311 9311 -2277
rect 9311 -2311 9343 -2277
rect 9381 -2311 9413 -2277
rect 9413 -2311 9415 -2277
rect 5231 -2315 5265 -2313
rect 5231 -2381 5265 -2353
rect 5231 -2387 5265 -2381
rect 5231 -2449 5265 -2425
rect 5231 -2459 5265 -2449
rect 5231 -2517 5265 -2497
rect 5231 -2531 5265 -2517
rect 5231 -2585 5265 -2569
rect 5231 -2603 5265 -2585
rect 872 -2653 906 -2641
rect 872 -2675 906 -2653
rect 1080 -2674 1082 -2640
rect 1082 -2674 1114 -2640
rect 1152 -2674 1184 -2640
rect 1184 -2674 1186 -2640
rect 1532 -2674 1534 -2640
rect 1534 -2674 1566 -2640
rect 1604 -2674 1636 -2640
rect 1636 -2674 1638 -2640
rect 1790 -2674 1792 -2640
rect 1792 -2674 1824 -2640
rect 1862 -2674 1894 -2640
rect 1894 -2674 1896 -2640
rect 2048 -2674 2050 -2640
rect 2050 -2674 2082 -2640
rect 2120 -2674 2152 -2640
rect 2152 -2674 2154 -2640
rect 2306 -2674 2308 -2640
rect 2308 -2674 2340 -2640
rect 2378 -2674 2410 -2640
rect 2410 -2674 2412 -2640
rect 2758 -2674 2760 -2640
rect 2760 -2674 2792 -2640
rect 2830 -2674 2862 -2640
rect 2862 -2674 2864 -2640
rect 3016 -2674 3018 -2640
rect 3018 -2674 3050 -2640
rect 3088 -2674 3120 -2640
rect 3120 -2674 3122 -2640
rect 3274 -2674 3276 -2640
rect 3276 -2674 3308 -2640
rect 3346 -2674 3378 -2640
rect 3378 -2674 3380 -2640
rect 3726 -2674 3728 -2640
rect 3728 -2674 3760 -2640
rect 3798 -2674 3830 -2640
rect 3830 -2674 3832 -2640
rect 3984 -2674 3986 -2640
rect 3986 -2674 4018 -2640
rect 4056 -2674 4088 -2640
rect 4088 -2674 4090 -2640
rect 4242 -2674 4244 -2640
rect 4244 -2674 4276 -2640
rect 4314 -2674 4346 -2640
rect 4346 -2674 4348 -2640
rect 4500 -2674 4502 -2640
rect 4502 -2674 4534 -2640
rect 4572 -2674 4604 -2640
rect 4604 -2674 4606 -2640
rect 4952 -2674 4954 -2640
rect 4954 -2674 4986 -2640
rect 5024 -2674 5056 -2640
rect 5056 -2674 5058 -2640
rect 9589 -2313 9623 -2281
rect 9589 -2315 9623 -2313
rect 9589 -2381 9623 -2353
rect 9589 -2387 9623 -2381
rect 9589 -2449 9623 -2425
rect 9589 -2459 9623 -2449
rect 9589 -2517 9623 -2497
rect 9589 -2531 9623 -2517
rect 9589 -2585 9623 -2569
rect 9589 -2603 9623 -2585
rect 872 -2721 906 -2713
rect 5231 -2653 5265 -2641
rect 5231 -2675 5265 -2653
rect 5438 -2674 5440 -2640
rect 5440 -2674 5472 -2640
rect 5510 -2674 5542 -2640
rect 5542 -2674 5544 -2640
rect 5889 -2674 5891 -2640
rect 5891 -2674 5923 -2640
rect 5961 -2674 5993 -2640
rect 5993 -2674 5995 -2640
rect 6147 -2674 6149 -2640
rect 6149 -2674 6181 -2640
rect 6219 -2674 6251 -2640
rect 6251 -2674 6253 -2640
rect 6405 -2674 6407 -2640
rect 6407 -2674 6439 -2640
rect 6477 -2674 6509 -2640
rect 6509 -2674 6511 -2640
rect 6663 -2674 6665 -2640
rect 6665 -2674 6697 -2640
rect 6735 -2674 6767 -2640
rect 6767 -2674 6769 -2640
rect 7115 -2674 7117 -2640
rect 7117 -2674 7149 -2640
rect 7187 -2674 7219 -2640
rect 7219 -2674 7221 -2640
rect 7373 -2674 7375 -2640
rect 7375 -2674 7407 -2640
rect 7445 -2674 7477 -2640
rect 7477 -2674 7479 -2640
rect 7631 -2674 7633 -2640
rect 7633 -2674 7665 -2640
rect 7703 -2674 7735 -2640
rect 7735 -2674 7737 -2640
rect 8083 -2674 8085 -2640
rect 8085 -2674 8117 -2640
rect 8155 -2674 8187 -2640
rect 8187 -2674 8189 -2640
rect 8341 -2674 8343 -2640
rect 8343 -2674 8375 -2640
rect 8413 -2674 8445 -2640
rect 8445 -2674 8447 -2640
rect 8599 -2674 8601 -2640
rect 8601 -2674 8633 -2640
rect 8671 -2674 8703 -2640
rect 8703 -2674 8705 -2640
rect 8857 -2674 8859 -2640
rect 8859 -2674 8891 -2640
rect 8929 -2674 8961 -2640
rect 8961 -2674 8963 -2640
rect 9309 -2674 9311 -2640
rect 9311 -2674 9343 -2640
rect 9381 -2674 9413 -2640
rect 9413 -2674 9415 -2640
rect 9589 -2653 9623 -2641
rect 872 -2747 906 -2721
rect 872 -2789 906 -2785
rect 872 -2819 906 -2789
rect 872 -2891 906 -2857
rect 987 -2770 1021 -2768
rect 987 -2802 1021 -2770
rect 987 -2872 1021 -2840
rect 987 -2874 1021 -2872
rect 1245 -2770 1279 -2768
rect 1245 -2802 1279 -2770
rect 1245 -2872 1279 -2840
rect 1245 -2874 1279 -2872
rect 1439 -2770 1473 -2768
rect 1439 -2802 1473 -2770
rect 1439 -2872 1473 -2840
rect 1439 -2874 1473 -2872
rect 1697 -2770 1731 -2768
rect 1697 -2802 1731 -2770
rect 1697 -2872 1731 -2840
rect 1697 -2874 1731 -2872
rect 1955 -2770 1989 -2768
rect 1955 -2802 1989 -2770
rect 1955 -2872 1989 -2840
rect 1955 -2874 1989 -2872
rect 2213 -2770 2247 -2768
rect 2213 -2802 2247 -2770
rect 2213 -2872 2247 -2840
rect 2213 -2874 2247 -2872
rect 2471 -2770 2505 -2768
rect 2471 -2802 2505 -2770
rect 2471 -2872 2505 -2840
rect 2471 -2874 2505 -2872
rect 2665 -2770 2699 -2768
rect 2665 -2802 2699 -2770
rect 2665 -2872 2699 -2840
rect 2665 -2874 2699 -2872
rect 2923 -2770 2957 -2768
rect 2923 -2802 2957 -2770
rect 2923 -2872 2957 -2840
rect 2923 -2874 2957 -2872
rect 3181 -2770 3215 -2768
rect 3181 -2802 3215 -2770
rect 3181 -2872 3215 -2840
rect 3181 -2874 3215 -2872
rect 3439 -2770 3473 -2768
rect 3439 -2802 3473 -2770
rect 3439 -2872 3473 -2840
rect 3439 -2874 3473 -2872
rect 3633 -2770 3667 -2768
rect 3633 -2802 3667 -2770
rect 3633 -2872 3667 -2840
rect 3633 -2874 3667 -2872
rect 3891 -2770 3925 -2768
rect 3891 -2802 3925 -2770
rect 3891 -2872 3925 -2840
rect 3891 -2874 3925 -2872
rect 4149 -2770 4183 -2768
rect 4149 -2802 4183 -2770
rect 4149 -2872 4183 -2840
rect 4149 -2874 4183 -2872
rect 4407 -2770 4441 -2768
rect 4407 -2802 4441 -2770
rect 4407 -2872 4441 -2840
rect 4407 -2874 4441 -2872
rect 4665 -2770 4699 -2768
rect 4665 -2802 4699 -2770
rect 4665 -2872 4699 -2840
rect 4665 -2874 4699 -2872
rect 4859 -2770 4893 -2768
rect 4859 -2802 4893 -2770
rect 4859 -2872 4893 -2840
rect 4859 -2874 4893 -2872
rect 5117 -2770 5151 -2768
rect 5117 -2802 5151 -2770
rect 5117 -2872 5151 -2840
rect 5117 -2874 5151 -2872
rect 5231 -2721 5265 -2713
rect 9589 -2675 9623 -2653
rect 5231 -2747 5265 -2721
rect 5231 -2789 5265 -2785
rect 5231 -2819 5265 -2789
rect 5231 -2891 5265 -2857
rect 5345 -2770 5379 -2768
rect 5345 -2802 5379 -2770
rect 5345 -2872 5379 -2840
rect 5345 -2874 5379 -2872
rect 5603 -2770 5637 -2768
rect 5603 -2802 5637 -2770
rect 5603 -2872 5637 -2840
rect 5603 -2874 5637 -2872
rect 5796 -2770 5830 -2768
rect 5796 -2802 5830 -2770
rect 5796 -2872 5830 -2840
rect 5796 -2874 5830 -2872
rect 6054 -2770 6088 -2768
rect 6054 -2802 6088 -2770
rect 6054 -2872 6088 -2840
rect 6054 -2874 6088 -2872
rect 6312 -2770 6346 -2768
rect 6312 -2802 6346 -2770
rect 6312 -2872 6346 -2840
rect 6312 -2874 6346 -2872
rect 6570 -2770 6604 -2768
rect 6570 -2802 6604 -2770
rect 6570 -2872 6604 -2840
rect 6570 -2874 6604 -2872
rect 6828 -2770 6862 -2768
rect 6828 -2802 6862 -2770
rect 6828 -2872 6862 -2840
rect 6828 -2874 6862 -2872
rect 7022 -2770 7056 -2768
rect 7022 -2802 7056 -2770
rect 7022 -2872 7056 -2840
rect 7022 -2874 7056 -2872
rect 7280 -2770 7314 -2768
rect 7280 -2802 7314 -2770
rect 7280 -2872 7314 -2840
rect 7280 -2874 7314 -2872
rect 7538 -2770 7572 -2768
rect 7538 -2802 7572 -2770
rect 7538 -2872 7572 -2840
rect 7538 -2874 7572 -2872
rect 7796 -2770 7830 -2768
rect 7796 -2802 7830 -2770
rect 7796 -2872 7830 -2840
rect 7796 -2874 7830 -2872
rect 7990 -2770 8024 -2768
rect 7990 -2802 8024 -2770
rect 7990 -2872 8024 -2840
rect 7990 -2874 8024 -2872
rect 8248 -2770 8282 -2768
rect 8248 -2802 8282 -2770
rect 8248 -2872 8282 -2840
rect 8248 -2874 8282 -2872
rect 8506 -2770 8540 -2768
rect 8506 -2802 8540 -2770
rect 8506 -2872 8540 -2840
rect 8506 -2874 8540 -2872
rect 8764 -2770 8798 -2768
rect 8764 -2802 8798 -2770
rect 8764 -2872 8798 -2840
rect 8764 -2874 8798 -2872
rect 9022 -2770 9056 -2768
rect 9022 -2802 9056 -2770
rect 9022 -2872 9056 -2840
rect 9022 -2874 9056 -2872
rect 9216 -2770 9250 -2768
rect 9216 -2802 9250 -2770
rect 9216 -2872 9250 -2840
rect 9216 -2874 9250 -2872
rect 9474 -2770 9508 -2768
rect 9474 -2802 9508 -2770
rect 9474 -2872 9508 -2840
rect 9474 -2874 9508 -2872
rect 9589 -2721 9623 -2713
rect 9589 -2747 9623 -2721
rect 9589 -2789 9623 -2785
rect 9589 -2819 9623 -2789
rect 9589 -2891 9623 -2857
rect 872 -2959 906 -2929
rect 872 -2963 906 -2959
rect 872 -3027 906 -3001
rect 872 -3035 906 -3027
rect 872 -3095 906 -3073
rect 872 -3107 906 -3095
rect 872 -3163 906 -3145
rect 872 -3179 906 -3163
rect 872 -3231 906 -3217
rect 872 -3251 906 -3231
rect 872 -3299 906 -3289
rect 5231 -2959 5265 -2929
rect 5231 -2963 5265 -2959
rect 5231 -3027 5265 -3001
rect 5231 -3035 5265 -3027
rect 5231 -3095 5265 -3073
rect 5231 -3107 5265 -3095
rect 5231 -3163 5265 -3145
rect 5231 -3179 5265 -3163
rect 5231 -3231 5265 -3217
rect 5231 -3251 5265 -3231
rect 5231 -3299 5265 -3289
rect 9589 -2959 9623 -2929
rect 9589 -2963 9623 -2959
rect 9589 -3027 9623 -3001
rect 9589 -3035 9623 -3027
rect 9589 -3095 9623 -3073
rect 9589 -3107 9623 -3095
rect 9589 -3163 9623 -3145
rect 9589 -3179 9623 -3163
rect 9589 -3231 9623 -3217
rect 9589 -3251 9623 -3231
rect 9589 -3299 9623 -3289
rect 872 -3323 906 -3299
rect 5231 -3323 5265 -3299
rect 9589 -3323 9623 -3299
rect 872 -3367 906 -3361
rect 872 -3395 906 -3367
rect 872 -3435 906 -3433
rect 872 -3467 906 -3435
rect 872 -3537 906 -3505
rect 872 -3539 906 -3537
rect 872 -3605 906 -3577
rect 872 -3611 906 -3605
rect 872 -3673 906 -3649
rect 872 -3683 906 -3673
rect 5231 -3367 5265 -3361
rect 5231 -3395 5265 -3367
rect 5231 -3435 5265 -3433
rect 5231 -3467 5265 -3435
rect 5231 -3537 5265 -3505
rect 5231 -3539 5265 -3537
rect 5231 -3605 5265 -3577
rect 5231 -3611 5265 -3605
rect 5231 -3673 5265 -3649
rect 5231 -3683 5265 -3673
rect 9589 -3367 9623 -3361
rect 9589 -3395 9623 -3367
rect 9589 -3435 9623 -3433
rect 9589 -3467 9623 -3435
rect 9589 -3537 9623 -3505
rect 9589 -3539 9623 -3537
rect 9589 -3605 9623 -3577
rect 9589 -3611 9623 -3605
rect 9589 -3673 9623 -3649
rect 9589 -3683 9623 -3673
rect 872 -3741 906 -3721
rect 872 -3755 906 -3741
rect 872 -3809 906 -3793
rect 872 -3827 906 -3809
rect 872 -3899 906 -3865
rect 987 -3760 1021 -3758
rect 987 -3792 1021 -3760
rect 987 -3862 1021 -3830
rect 987 -3864 1021 -3862
rect 1245 -3760 1279 -3758
rect 1245 -3792 1279 -3760
rect 1245 -3862 1279 -3830
rect 1245 -3864 1279 -3862
rect 1439 -3760 1473 -3758
rect 1439 -3792 1473 -3760
rect 1439 -3862 1473 -3830
rect 1439 -3864 1473 -3862
rect 1697 -3760 1731 -3758
rect 1697 -3792 1731 -3760
rect 1697 -3862 1731 -3830
rect 1697 -3864 1731 -3862
rect 1955 -3760 1989 -3758
rect 1955 -3792 1989 -3760
rect 1955 -3862 1989 -3830
rect 1955 -3864 1989 -3862
rect 2213 -3760 2247 -3758
rect 2213 -3792 2247 -3760
rect 2213 -3862 2247 -3830
rect 2213 -3864 2247 -3862
rect 2471 -3760 2505 -3758
rect 2471 -3792 2505 -3760
rect 2471 -3862 2505 -3830
rect 2471 -3864 2505 -3862
rect 2665 -3760 2699 -3758
rect 2665 -3792 2699 -3760
rect 2665 -3862 2699 -3830
rect 2665 -3864 2699 -3862
rect 2923 -3760 2957 -3758
rect 2923 -3792 2957 -3760
rect 2923 -3862 2957 -3830
rect 2923 -3864 2957 -3862
rect 3181 -3760 3215 -3758
rect 3181 -3792 3215 -3760
rect 3181 -3862 3215 -3830
rect 3181 -3864 3215 -3862
rect 3439 -3760 3473 -3758
rect 3439 -3792 3473 -3760
rect 3439 -3862 3473 -3830
rect 3439 -3864 3473 -3862
rect 3633 -3760 3667 -3758
rect 3633 -3792 3667 -3760
rect 3633 -3862 3667 -3830
rect 3633 -3864 3667 -3862
rect 3891 -3760 3925 -3758
rect 3891 -3792 3925 -3760
rect 3891 -3862 3925 -3830
rect 3891 -3864 3925 -3862
rect 4149 -3760 4183 -3758
rect 4149 -3792 4183 -3760
rect 4149 -3862 4183 -3830
rect 4149 -3864 4183 -3862
rect 4407 -3760 4441 -3758
rect 4407 -3792 4441 -3760
rect 4407 -3862 4441 -3830
rect 4407 -3864 4441 -3862
rect 4665 -3760 4699 -3758
rect 4665 -3792 4699 -3760
rect 4665 -3862 4699 -3830
rect 4665 -3864 4699 -3862
rect 4859 -3760 4893 -3758
rect 4859 -3792 4893 -3760
rect 4859 -3862 4893 -3830
rect 4859 -3864 4893 -3862
rect 5117 -3760 5151 -3758
rect 5117 -3792 5151 -3760
rect 5117 -3862 5151 -3830
rect 5117 -3864 5151 -3862
rect 5231 -3741 5265 -3721
rect 5231 -3755 5265 -3741
rect 5231 -3809 5265 -3793
rect 5231 -3827 5265 -3809
rect 5231 -3899 5265 -3865
rect 872 -3971 906 -3937
rect 5345 -3760 5379 -3758
rect 5345 -3792 5379 -3760
rect 5345 -3862 5379 -3830
rect 5345 -3864 5379 -3862
rect 5603 -3760 5637 -3758
rect 5603 -3792 5637 -3760
rect 5603 -3862 5637 -3830
rect 5603 -3864 5637 -3862
rect 5796 -3760 5830 -3758
rect 5796 -3792 5830 -3760
rect 5796 -3862 5830 -3830
rect 5796 -3864 5830 -3862
rect 6054 -3760 6088 -3758
rect 6054 -3792 6088 -3760
rect 6054 -3862 6088 -3830
rect 6054 -3864 6088 -3862
rect 6312 -3760 6346 -3758
rect 6312 -3792 6346 -3760
rect 6312 -3862 6346 -3830
rect 6312 -3864 6346 -3862
rect 6570 -3760 6604 -3758
rect 6570 -3792 6604 -3760
rect 6570 -3862 6604 -3830
rect 6570 -3864 6604 -3862
rect 6828 -3760 6862 -3758
rect 6828 -3792 6862 -3760
rect 6828 -3862 6862 -3830
rect 6828 -3864 6862 -3862
rect 7022 -3760 7056 -3758
rect 7022 -3792 7056 -3760
rect 7022 -3862 7056 -3830
rect 7022 -3864 7056 -3862
rect 7280 -3760 7314 -3758
rect 7280 -3792 7314 -3760
rect 7280 -3862 7314 -3830
rect 7280 -3864 7314 -3862
rect 7538 -3760 7572 -3758
rect 7538 -3792 7572 -3760
rect 7538 -3862 7572 -3830
rect 7538 -3864 7572 -3862
rect 7796 -3760 7830 -3758
rect 7796 -3792 7830 -3760
rect 7796 -3862 7830 -3830
rect 7796 -3864 7830 -3862
rect 7990 -3760 8024 -3758
rect 7990 -3792 8024 -3760
rect 7990 -3862 8024 -3830
rect 7990 -3864 8024 -3862
rect 8248 -3760 8282 -3758
rect 8248 -3792 8282 -3760
rect 8248 -3862 8282 -3830
rect 8248 -3864 8282 -3862
rect 8506 -3760 8540 -3758
rect 8506 -3792 8540 -3760
rect 8506 -3862 8540 -3830
rect 8506 -3864 8540 -3862
rect 8764 -3760 8798 -3758
rect 8764 -3792 8798 -3760
rect 8764 -3862 8798 -3830
rect 8764 -3864 8798 -3862
rect 9022 -3760 9056 -3758
rect 9022 -3792 9056 -3760
rect 9022 -3862 9056 -3830
rect 9022 -3864 9056 -3862
rect 9216 -3760 9250 -3758
rect 9216 -3792 9250 -3760
rect 9216 -3862 9250 -3830
rect 9216 -3864 9250 -3862
rect 9474 -3760 9508 -3758
rect 9474 -3792 9508 -3760
rect 9474 -3862 9508 -3830
rect 9474 -3864 9508 -3862
rect 9589 -3741 9623 -3721
rect 9589 -3755 9623 -3741
rect 9589 -3809 9623 -3793
rect 9589 -3827 9623 -3809
rect 9589 -3899 9623 -3865
rect 1080 -3992 1082 -3958
rect 1082 -3992 1114 -3958
rect 1152 -3992 1184 -3958
rect 1184 -3992 1186 -3958
rect 1532 -3992 1534 -3958
rect 1534 -3992 1566 -3958
rect 1604 -3992 1636 -3958
rect 1636 -3992 1638 -3958
rect 1790 -3992 1792 -3958
rect 1792 -3992 1824 -3958
rect 1862 -3992 1894 -3958
rect 1894 -3992 1896 -3958
rect 2048 -3992 2050 -3958
rect 2050 -3992 2082 -3958
rect 2120 -3992 2152 -3958
rect 2152 -3992 2154 -3958
rect 2306 -3992 2308 -3958
rect 2308 -3992 2340 -3958
rect 2378 -3992 2410 -3958
rect 2410 -3992 2412 -3958
rect 2758 -3992 2760 -3958
rect 2760 -3992 2792 -3958
rect 2830 -3992 2862 -3958
rect 2862 -3992 2864 -3958
rect 3016 -3992 3018 -3958
rect 3018 -3992 3050 -3958
rect 3088 -3992 3120 -3958
rect 3120 -3992 3122 -3958
rect 3274 -3992 3276 -3958
rect 3276 -3992 3308 -3958
rect 3346 -3992 3378 -3958
rect 3378 -3992 3380 -3958
rect 3726 -3992 3728 -3958
rect 3728 -3992 3760 -3958
rect 3798 -3992 3830 -3958
rect 3830 -3992 3832 -3958
rect 3984 -3992 3986 -3958
rect 3986 -3992 4018 -3958
rect 4056 -3992 4088 -3958
rect 4088 -3992 4090 -3958
rect 4242 -3992 4244 -3958
rect 4244 -3992 4276 -3958
rect 4314 -3992 4346 -3958
rect 4346 -3992 4348 -3958
rect 4500 -3992 4502 -3958
rect 4502 -3992 4534 -3958
rect 4572 -3992 4604 -3958
rect 4604 -3992 4606 -3958
rect 4952 -3992 4954 -3958
rect 4954 -3992 4986 -3958
rect 5024 -3992 5056 -3958
rect 5056 -3992 5058 -3958
rect 5231 -3971 5265 -3937
rect 872 -4043 906 -4009
rect 5438 -3992 5440 -3958
rect 5440 -3992 5472 -3958
rect 5510 -3992 5542 -3958
rect 5542 -3992 5544 -3958
rect 5889 -3992 5891 -3958
rect 5891 -3992 5923 -3958
rect 5961 -3992 5993 -3958
rect 5993 -3992 5995 -3958
rect 6147 -3992 6149 -3958
rect 6149 -3992 6181 -3958
rect 6219 -3992 6251 -3958
rect 6251 -3992 6253 -3958
rect 6405 -3992 6407 -3958
rect 6407 -3992 6439 -3958
rect 6477 -3992 6509 -3958
rect 6509 -3992 6511 -3958
rect 6663 -3992 6665 -3958
rect 6665 -3992 6697 -3958
rect 6735 -3992 6767 -3958
rect 6767 -3992 6769 -3958
rect 7115 -3992 7117 -3958
rect 7117 -3992 7149 -3958
rect 7187 -3992 7219 -3958
rect 7219 -3992 7221 -3958
rect 7373 -3992 7375 -3958
rect 7375 -3992 7407 -3958
rect 7445 -3992 7477 -3958
rect 7477 -3992 7479 -3958
rect 7631 -3992 7633 -3958
rect 7633 -3992 7665 -3958
rect 7703 -3992 7735 -3958
rect 7735 -3992 7737 -3958
rect 8083 -3992 8085 -3958
rect 8085 -3992 8117 -3958
rect 8155 -3992 8187 -3958
rect 8187 -3992 8189 -3958
rect 8341 -3992 8343 -3958
rect 8343 -3992 8375 -3958
rect 8413 -3992 8445 -3958
rect 8445 -3992 8447 -3958
rect 8599 -3992 8601 -3958
rect 8601 -3992 8633 -3958
rect 8671 -3992 8703 -3958
rect 8703 -3992 8705 -3958
rect 8857 -3992 8859 -3958
rect 8859 -3992 8891 -3958
rect 8929 -3992 8961 -3958
rect 8961 -3992 8963 -3958
rect 9309 -3992 9311 -3958
rect 9311 -3992 9343 -3958
rect 9381 -3992 9413 -3958
rect 9413 -3992 9415 -3958
rect 9589 -3971 9623 -3937
rect 5231 -4043 5265 -4009
rect 9589 -4043 9623 -4009
rect 946 -4106 980 -4072
rect 1018 -4106 1027 -4072
rect 1027 -4106 1052 -4072
rect 1090 -4106 1095 -4072
rect 1095 -4106 1124 -4072
rect 1162 -4106 1163 -4072
rect 1163 -4106 1196 -4072
rect 1234 -4106 1265 -4072
rect 1265 -4106 1268 -4072
rect 1306 -4106 1333 -4072
rect 1333 -4106 1340 -4072
rect 1378 -4106 1401 -4072
rect 1401 -4106 1412 -4072
rect 1450 -4106 1469 -4072
rect 1469 -4106 1484 -4072
rect 1522 -4106 1537 -4072
rect 1537 -4106 1556 -4072
rect 1594 -4106 1605 -4072
rect 1605 -4106 1628 -4072
rect 1666 -4106 1673 -4072
rect 1673 -4106 1700 -4072
rect 1738 -4106 1741 -4072
rect 1741 -4106 1772 -4072
rect 1810 -4106 1843 -4072
rect 1843 -4106 1844 -4072
rect 1882 -4106 1911 -4072
rect 1911 -4106 1916 -4072
rect 1954 -4106 1979 -4072
rect 1979 -4106 1988 -4072
rect 2026 -4106 2047 -4072
rect 2047 -4106 2060 -4072
rect 2098 -4106 2115 -4072
rect 2115 -4106 2132 -4072
rect 2170 -4106 2183 -4072
rect 2183 -4106 2204 -4072
rect 2242 -4106 2251 -4072
rect 2251 -4106 2276 -4072
rect 2314 -4106 2319 -4072
rect 2319 -4106 2348 -4072
rect 2386 -4106 2387 -4072
rect 2387 -4106 2420 -4072
rect 2458 -4106 2489 -4072
rect 2489 -4106 2492 -4072
rect 2530 -4106 2557 -4072
rect 2557 -4106 2564 -4072
rect 2602 -4106 2625 -4072
rect 2625 -4106 2636 -4072
rect 2674 -4106 2693 -4072
rect 2693 -4106 2708 -4072
rect 2746 -4106 2761 -4072
rect 2761 -4106 2780 -4072
rect 2818 -4106 2829 -4072
rect 2829 -4106 2852 -4072
rect 2890 -4106 2897 -4072
rect 2897 -4106 2924 -4072
rect 2962 -4106 2965 -4072
rect 2965 -4106 2996 -4072
rect 3034 -4106 3067 -4072
rect 3067 -4106 3068 -4072
rect 3106 -4106 3135 -4072
rect 3135 -4106 3140 -4072
rect 3178 -4106 3203 -4072
rect 3203 -4106 3212 -4072
rect 3250 -4106 3271 -4072
rect 3271 -4106 3284 -4072
rect 3322 -4106 3339 -4072
rect 3339 -4106 3356 -4072
rect 3394 -4106 3407 -4072
rect 3407 -4106 3428 -4072
rect 3466 -4106 3475 -4072
rect 3475 -4106 3500 -4072
rect 3538 -4106 3543 -4072
rect 3543 -4106 3572 -4072
rect 3610 -4106 3611 -4072
rect 3611 -4106 3644 -4072
rect 3682 -4106 3713 -4072
rect 3713 -4106 3716 -4072
rect 3754 -4106 3781 -4072
rect 3781 -4106 3788 -4072
rect 3826 -4106 3849 -4072
rect 3849 -4106 3860 -4072
rect 3898 -4106 3917 -4072
rect 3917 -4106 3932 -4072
rect 3970 -4106 3985 -4072
rect 3985 -4106 4004 -4072
rect 4042 -4106 4053 -4072
rect 4053 -4106 4076 -4072
rect 4114 -4106 4121 -4072
rect 4121 -4106 4148 -4072
rect 4186 -4106 4189 -4072
rect 4189 -4106 4220 -4072
rect 4258 -4106 4291 -4072
rect 4291 -4106 4292 -4072
rect 4330 -4106 4359 -4072
rect 4359 -4106 4364 -4072
rect 4402 -4106 4427 -4072
rect 4427 -4106 4436 -4072
rect 4474 -4106 4495 -4072
rect 4495 -4106 4508 -4072
rect 4546 -4106 4563 -4072
rect 4563 -4106 4580 -4072
rect 4618 -4106 4631 -4072
rect 4631 -4106 4652 -4072
rect 4690 -4106 4699 -4072
rect 4699 -4106 4724 -4072
rect 4762 -4106 4767 -4072
rect 4767 -4106 4796 -4072
rect 4834 -4106 4835 -4072
rect 4835 -4106 4868 -4072
rect 4906 -4106 4937 -4072
rect 4937 -4106 4940 -4072
rect 4978 -4106 5005 -4072
rect 5005 -4106 5012 -4072
rect 5050 -4106 5073 -4072
rect 5073 -4106 5084 -4072
rect 5122 -4106 5156 -4072
rect 5339 -4106 5373 -4072
rect 5411 -4106 5422 -4072
rect 5422 -4106 5445 -4072
rect 5483 -4106 5490 -4072
rect 5490 -4106 5517 -4072
rect 5555 -4106 5558 -4072
rect 5558 -4106 5589 -4072
rect 5627 -4106 5660 -4072
rect 5660 -4106 5661 -4072
rect 5699 -4106 5728 -4072
rect 5728 -4106 5733 -4072
rect 5771 -4106 5796 -4072
rect 5796 -4106 5805 -4072
rect 5843 -4106 5864 -4072
rect 5864 -4106 5877 -4072
rect 5915 -4106 5932 -4072
rect 5932 -4106 5949 -4072
rect 5987 -4106 6000 -4072
rect 6000 -4106 6021 -4072
rect 6059 -4106 6068 -4072
rect 6068 -4106 6093 -4072
rect 6131 -4106 6136 -4072
rect 6136 -4106 6165 -4072
rect 6203 -4106 6204 -4072
rect 6204 -4106 6237 -4072
rect 6275 -4106 6306 -4072
rect 6306 -4106 6309 -4072
rect 6347 -4106 6374 -4072
rect 6374 -4106 6381 -4072
rect 6419 -4106 6442 -4072
rect 6442 -4106 6453 -4072
rect 6491 -4106 6510 -4072
rect 6510 -4106 6525 -4072
rect 6563 -4106 6578 -4072
rect 6578 -4106 6597 -4072
rect 6635 -4106 6646 -4072
rect 6646 -4106 6669 -4072
rect 6707 -4106 6714 -4072
rect 6714 -4106 6741 -4072
rect 6779 -4106 6782 -4072
rect 6782 -4106 6813 -4072
rect 6851 -4106 6884 -4072
rect 6884 -4106 6885 -4072
rect 6923 -4106 6952 -4072
rect 6952 -4106 6957 -4072
rect 6995 -4106 7020 -4072
rect 7020 -4106 7029 -4072
rect 7067 -4106 7088 -4072
rect 7088 -4106 7101 -4072
rect 7139 -4106 7156 -4072
rect 7156 -4106 7173 -4072
rect 7211 -4106 7224 -4072
rect 7224 -4106 7245 -4072
rect 7283 -4106 7292 -4072
rect 7292 -4106 7317 -4072
rect 7355 -4106 7360 -4072
rect 7360 -4106 7389 -4072
rect 7427 -4106 7428 -4072
rect 7428 -4106 7461 -4072
rect 7499 -4106 7530 -4072
rect 7530 -4106 7533 -4072
rect 7571 -4106 7598 -4072
rect 7598 -4106 7605 -4072
rect 7643 -4106 7666 -4072
rect 7666 -4106 7677 -4072
rect 7715 -4106 7734 -4072
rect 7734 -4106 7749 -4072
rect 7787 -4106 7802 -4072
rect 7802 -4106 7821 -4072
rect 7859 -4106 7870 -4072
rect 7870 -4106 7893 -4072
rect 7931 -4106 7938 -4072
rect 7938 -4106 7965 -4072
rect 8003 -4106 8006 -4072
rect 8006 -4106 8037 -4072
rect 8075 -4106 8108 -4072
rect 8108 -4106 8109 -4072
rect 8147 -4106 8176 -4072
rect 8176 -4106 8181 -4072
rect 8219 -4106 8244 -4072
rect 8244 -4106 8253 -4072
rect 8291 -4106 8312 -4072
rect 8312 -4106 8325 -4072
rect 8363 -4106 8380 -4072
rect 8380 -4106 8397 -4072
rect 8435 -4106 8448 -4072
rect 8448 -4106 8469 -4072
rect 8507 -4106 8516 -4072
rect 8516 -4106 8541 -4072
rect 8579 -4106 8584 -4072
rect 8584 -4106 8613 -4072
rect 8651 -4106 8652 -4072
rect 8652 -4106 8685 -4072
rect 8723 -4106 8754 -4072
rect 8754 -4106 8757 -4072
rect 8795 -4106 8822 -4072
rect 8822 -4106 8829 -4072
rect 8867 -4106 8890 -4072
rect 8890 -4106 8901 -4072
rect 8939 -4106 8958 -4072
rect 8958 -4106 8973 -4072
rect 9011 -4106 9026 -4072
rect 9026 -4106 9045 -4072
rect 9083 -4106 9094 -4072
rect 9094 -4106 9117 -4072
rect 9155 -4106 9162 -4072
rect 9162 -4106 9189 -4072
rect 9227 -4106 9230 -4072
rect 9230 -4106 9261 -4072
rect 9299 -4106 9332 -4072
rect 9332 -4106 9333 -4072
rect 9371 -4106 9400 -4072
rect 9400 -4106 9405 -4072
rect 9443 -4106 9468 -4072
rect 9468 -4106 9477 -4072
rect 9515 -4106 9549 -4072
rect 872 -4169 906 -4135
rect 5231 -4169 5265 -4135
rect 872 -4241 906 -4207
rect 1080 -4220 1082 -4186
rect 1082 -4220 1114 -4186
rect 1152 -4220 1184 -4186
rect 1184 -4220 1186 -4186
rect 1532 -4220 1534 -4186
rect 1534 -4220 1566 -4186
rect 1604 -4220 1636 -4186
rect 1636 -4220 1638 -4186
rect 1790 -4220 1792 -4186
rect 1792 -4220 1824 -4186
rect 1862 -4220 1894 -4186
rect 1894 -4220 1896 -4186
rect 2048 -4220 2050 -4186
rect 2050 -4220 2082 -4186
rect 2120 -4220 2152 -4186
rect 2152 -4220 2154 -4186
rect 2306 -4220 2308 -4186
rect 2308 -4220 2340 -4186
rect 2378 -4220 2410 -4186
rect 2410 -4220 2412 -4186
rect 2758 -4220 2760 -4186
rect 2760 -4220 2792 -4186
rect 2830 -4220 2862 -4186
rect 2862 -4220 2864 -4186
rect 3016 -4220 3018 -4186
rect 3018 -4220 3050 -4186
rect 3088 -4220 3120 -4186
rect 3120 -4220 3122 -4186
rect 3274 -4220 3276 -4186
rect 3276 -4220 3308 -4186
rect 3346 -4220 3378 -4186
rect 3378 -4220 3380 -4186
rect 3726 -4220 3728 -4186
rect 3728 -4220 3760 -4186
rect 3798 -4220 3830 -4186
rect 3830 -4220 3832 -4186
rect 3984 -4220 3986 -4186
rect 3986 -4220 4018 -4186
rect 4056 -4220 4088 -4186
rect 4088 -4220 4090 -4186
rect 4242 -4220 4244 -4186
rect 4244 -4220 4276 -4186
rect 4314 -4220 4346 -4186
rect 4346 -4220 4348 -4186
rect 4500 -4220 4502 -4186
rect 4502 -4220 4534 -4186
rect 4572 -4220 4604 -4186
rect 4604 -4220 4606 -4186
rect 4952 -4220 4954 -4186
rect 4954 -4220 4986 -4186
rect 5024 -4220 5056 -4186
rect 5056 -4220 5058 -4186
rect 9589 -4169 9623 -4135
rect 5231 -4241 5265 -4207
rect 5438 -4220 5440 -4186
rect 5440 -4220 5472 -4186
rect 5510 -4220 5542 -4186
rect 5542 -4220 5544 -4186
rect 5889 -4220 5891 -4186
rect 5891 -4220 5923 -4186
rect 5961 -4220 5993 -4186
rect 5993 -4220 5995 -4186
rect 6147 -4220 6149 -4186
rect 6149 -4220 6181 -4186
rect 6219 -4220 6251 -4186
rect 6251 -4220 6253 -4186
rect 6405 -4220 6407 -4186
rect 6407 -4220 6439 -4186
rect 6477 -4220 6509 -4186
rect 6509 -4220 6511 -4186
rect 6663 -4220 6665 -4186
rect 6665 -4220 6697 -4186
rect 6735 -4220 6767 -4186
rect 6767 -4220 6769 -4186
rect 7115 -4220 7117 -4186
rect 7117 -4220 7149 -4186
rect 7187 -4220 7219 -4186
rect 7219 -4220 7221 -4186
rect 7373 -4220 7375 -4186
rect 7375 -4220 7407 -4186
rect 7445 -4220 7477 -4186
rect 7477 -4220 7479 -4186
rect 7631 -4220 7633 -4186
rect 7633 -4220 7665 -4186
rect 7703 -4220 7735 -4186
rect 7735 -4220 7737 -4186
rect 8083 -4220 8085 -4186
rect 8085 -4220 8117 -4186
rect 8155 -4220 8187 -4186
rect 8187 -4220 8189 -4186
rect 8341 -4220 8343 -4186
rect 8343 -4220 8375 -4186
rect 8413 -4220 8445 -4186
rect 8445 -4220 8447 -4186
rect 8599 -4220 8601 -4186
rect 8601 -4220 8633 -4186
rect 8671 -4220 8703 -4186
rect 8703 -4220 8705 -4186
rect 8857 -4220 8859 -4186
rect 8859 -4220 8891 -4186
rect 8929 -4220 8961 -4186
rect 8961 -4220 8963 -4186
rect 9309 -4220 9311 -4186
rect 9311 -4220 9343 -4186
rect 9381 -4220 9413 -4186
rect 9413 -4220 9415 -4186
rect 872 -4313 906 -4279
rect 872 -4369 906 -4351
rect 872 -4385 906 -4369
rect 872 -4437 906 -4423
rect 872 -4457 906 -4437
rect 987 -4316 1021 -4314
rect 987 -4348 1021 -4316
rect 987 -4418 1021 -4386
rect 987 -4420 1021 -4418
rect 1245 -4316 1279 -4314
rect 1245 -4348 1279 -4316
rect 1245 -4418 1279 -4386
rect 1245 -4420 1279 -4418
rect 1439 -4316 1473 -4314
rect 1439 -4348 1473 -4316
rect 1439 -4418 1473 -4386
rect 1439 -4420 1473 -4418
rect 1697 -4316 1731 -4314
rect 1697 -4348 1731 -4316
rect 1697 -4418 1731 -4386
rect 1697 -4420 1731 -4418
rect 1955 -4316 1989 -4314
rect 1955 -4348 1989 -4316
rect 1955 -4418 1989 -4386
rect 1955 -4420 1989 -4418
rect 2213 -4316 2247 -4314
rect 2213 -4348 2247 -4316
rect 2213 -4418 2247 -4386
rect 2213 -4420 2247 -4418
rect 2471 -4316 2505 -4314
rect 2471 -4348 2505 -4316
rect 2471 -4418 2505 -4386
rect 2471 -4420 2505 -4418
rect 2665 -4316 2699 -4314
rect 2665 -4348 2699 -4316
rect 2665 -4418 2699 -4386
rect 2665 -4420 2699 -4418
rect 2923 -4316 2957 -4314
rect 2923 -4348 2957 -4316
rect 2923 -4418 2957 -4386
rect 2923 -4420 2957 -4418
rect 3181 -4316 3215 -4314
rect 3181 -4348 3215 -4316
rect 3181 -4418 3215 -4386
rect 3181 -4420 3215 -4418
rect 3439 -4316 3473 -4314
rect 3439 -4348 3473 -4316
rect 3439 -4418 3473 -4386
rect 3439 -4420 3473 -4418
rect 3633 -4316 3667 -4314
rect 3633 -4348 3667 -4316
rect 3633 -4418 3667 -4386
rect 3633 -4420 3667 -4418
rect 3891 -4316 3925 -4314
rect 3891 -4348 3925 -4316
rect 3891 -4418 3925 -4386
rect 3891 -4420 3925 -4418
rect 4149 -4316 4183 -4314
rect 4149 -4348 4183 -4316
rect 4149 -4418 4183 -4386
rect 4149 -4420 4183 -4418
rect 4407 -4316 4441 -4314
rect 4407 -4348 4441 -4316
rect 4407 -4418 4441 -4386
rect 4407 -4420 4441 -4418
rect 4665 -4316 4699 -4314
rect 4665 -4348 4699 -4316
rect 4665 -4418 4699 -4386
rect 4665 -4420 4699 -4418
rect 4859 -4316 4893 -4314
rect 4859 -4348 4893 -4316
rect 4859 -4418 4893 -4386
rect 4859 -4420 4893 -4418
rect 5117 -4316 5151 -4314
rect 5117 -4348 5151 -4316
rect 5117 -4418 5151 -4386
rect 5117 -4420 5151 -4418
rect 9589 -4241 9623 -4207
rect 5231 -4313 5265 -4279
rect 5231 -4369 5265 -4351
rect 5231 -4385 5265 -4369
rect 5231 -4437 5265 -4423
rect 5231 -4457 5265 -4437
rect 5345 -4316 5379 -4314
rect 5345 -4348 5379 -4316
rect 5345 -4418 5379 -4386
rect 5345 -4420 5379 -4418
rect 5603 -4316 5637 -4314
rect 5603 -4348 5637 -4316
rect 5603 -4418 5637 -4386
rect 5603 -4420 5637 -4418
rect 5796 -4316 5830 -4314
rect 5796 -4348 5830 -4316
rect 5796 -4418 5830 -4386
rect 5796 -4420 5830 -4418
rect 6054 -4316 6088 -4314
rect 6054 -4348 6088 -4316
rect 6054 -4418 6088 -4386
rect 6054 -4420 6088 -4418
rect 6312 -4316 6346 -4314
rect 6312 -4348 6346 -4316
rect 6312 -4418 6346 -4386
rect 6312 -4420 6346 -4418
rect 6570 -4316 6604 -4314
rect 6570 -4348 6604 -4316
rect 6570 -4418 6604 -4386
rect 6570 -4420 6604 -4418
rect 6828 -4316 6862 -4314
rect 6828 -4348 6862 -4316
rect 6828 -4418 6862 -4386
rect 6828 -4420 6862 -4418
rect 7022 -4316 7056 -4314
rect 7022 -4348 7056 -4316
rect 7022 -4418 7056 -4386
rect 7022 -4420 7056 -4418
rect 7280 -4316 7314 -4314
rect 7280 -4348 7314 -4316
rect 7280 -4418 7314 -4386
rect 7280 -4420 7314 -4418
rect 7538 -4316 7572 -4314
rect 7538 -4348 7572 -4316
rect 7538 -4418 7572 -4386
rect 7538 -4420 7572 -4418
rect 7796 -4316 7830 -4314
rect 7796 -4348 7830 -4316
rect 7796 -4418 7830 -4386
rect 7796 -4420 7830 -4418
rect 7990 -4316 8024 -4314
rect 7990 -4348 8024 -4316
rect 7990 -4418 8024 -4386
rect 7990 -4420 8024 -4418
rect 8248 -4316 8282 -4314
rect 8248 -4348 8282 -4316
rect 8248 -4418 8282 -4386
rect 8248 -4420 8282 -4418
rect 8506 -4316 8540 -4314
rect 8506 -4348 8540 -4316
rect 8506 -4418 8540 -4386
rect 8506 -4420 8540 -4418
rect 8764 -4316 8798 -4314
rect 8764 -4348 8798 -4316
rect 8764 -4418 8798 -4386
rect 8764 -4420 8798 -4418
rect 9022 -4316 9056 -4314
rect 9022 -4348 9056 -4316
rect 9022 -4418 9056 -4386
rect 9022 -4420 9056 -4418
rect 9216 -4316 9250 -4314
rect 9216 -4348 9250 -4316
rect 9216 -4418 9250 -4386
rect 9216 -4420 9250 -4418
rect 9474 -4316 9508 -4314
rect 9474 -4348 9508 -4316
rect 9474 -4418 9508 -4386
rect 9474 -4420 9508 -4418
rect 9589 -4313 9623 -4279
rect 9589 -4369 9623 -4351
rect 9589 -4385 9623 -4369
rect 9589 -4437 9623 -4423
rect 9589 -4457 9623 -4437
rect 872 -4505 906 -4495
rect 872 -4529 906 -4505
rect 872 -4573 906 -4567
rect 872 -4601 906 -4573
rect 872 -4641 906 -4639
rect 872 -4673 906 -4641
rect 872 -4743 906 -4711
rect 872 -4745 906 -4743
rect 872 -4811 906 -4783
rect 872 -4817 906 -4811
rect 5231 -4505 5265 -4495
rect 5231 -4529 5265 -4505
rect 5231 -4573 5265 -4567
rect 5231 -4601 5265 -4573
rect 5231 -4641 5265 -4639
rect 5231 -4673 5265 -4641
rect 5231 -4743 5265 -4711
rect 5231 -4745 5265 -4743
rect 5231 -4811 5265 -4783
rect 5231 -4817 5265 -4811
rect 9589 -4505 9623 -4495
rect 9589 -4529 9623 -4505
rect 9589 -4573 9623 -4567
rect 9589 -4601 9623 -4573
rect 9589 -4641 9623 -4639
rect 9589 -4673 9623 -4641
rect 9589 -4743 9623 -4711
rect 9589 -4745 9623 -4743
rect 9589 -4811 9623 -4783
rect 9589 -4817 9623 -4811
rect 872 -4879 906 -4855
rect 5231 -4879 5265 -4855
rect 9589 -4879 9623 -4855
rect 872 -4889 906 -4879
rect 872 -4947 906 -4927
rect 872 -4961 906 -4947
rect 872 -5015 906 -4999
rect 872 -5033 906 -5015
rect 872 -5083 906 -5071
rect 872 -5105 906 -5083
rect 872 -5151 906 -5143
rect 872 -5177 906 -5151
rect 872 -5219 906 -5215
rect 872 -5249 906 -5219
rect 5231 -4889 5265 -4879
rect 5231 -4947 5265 -4927
rect 5231 -4961 5265 -4947
rect 5231 -5015 5265 -4999
rect 5231 -5033 5265 -5015
rect 5231 -5083 5265 -5071
rect 5231 -5105 5265 -5083
rect 5231 -5151 5265 -5143
rect 5231 -5177 5265 -5151
rect 5231 -5219 5265 -5215
rect 5231 -5249 5265 -5219
rect 9589 -4889 9623 -4879
rect 9589 -4947 9623 -4927
rect 9589 -4961 9623 -4947
rect 9589 -5015 9623 -4999
rect 9589 -5033 9623 -5015
rect 9589 -5083 9623 -5071
rect 9589 -5105 9623 -5083
rect 9589 -5151 9623 -5143
rect 9589 -5177 9623 -5151
rect 9589 -5219 9623 -5215
rect 9589 -5249 9623 -5219
rect 872 -5321 906 -5287
rect 872 -5389 906 -5359
rect 872 -5393 906 -5389
rect 872 -5457 906 -5431
rect 872 -5465 906 -5457
rect 987 -5306 1021 -5304
rect 987 -5338 1021 -5306
rect 987 -5408 1021 -5376
rect 987 -5410 1021 -5408
rect 1245 -5306 1279 -5304
rect 1245 -5338 1279 -5306
rect 1245 -5408 1279 -5376
rect 1245 -5410 1279 -5408
rect 1439 -5306 1473 -5304
rect 1439 -5338 1473 -5306
rect 1439 -5408 1473 -5376
rect 1439 -5410 1473 -5408
rect 1697 -5306 1731 -5304
rect 1697 -5338 1731 -5306
rect 1697 -5408 1731 -5376
rect 1697 -5410 1731 -5408
rect 1955 -5306 1989 -5304
rect 1955 -5338 1989 -5306
rect 1955 -5408 1989 -5376
rect 1955 -5410 1989 -5408
rect 2213 -5306 2247 -5304
rect 2213 -5338 2247 -5306
rect 2213 -5408 2247 -5376
rect 2213 -5410 2247 -5408
rect 2471 -5306 2505 -5304
rect 2471 -5338 2505 -5306
rect 2471 -5408 2505 -5376
rect 2471 -5410 2505 -5408
rect 2665 -5306 2699 -5304
rect 2665 -5338 2699 -5306
rect 2665 -5408 2699 -5376
rect 2665 -5410 2699 -5408
rect 2923 -5306 2957 -5304
rect 2923 -5338 2957 -5306
rect 2923 -5408 2957 -5376
rect 2923 -5410 2957 -5408
rect 3181 -5306 3215 -5304
rect 3181 -5338 3215 -5306
rect 3181 -5408 3215 -5376
rect 3181 -5410 3215 -5408
rect 3439 -5306 3473 -5304
rect 3439 -5338 3473 -5306
rect 3439 -5408 3473 -5376
rect 3439 -5410 3473 -5408
rect 3633 -5306 3667 -5304
rect 3633 -5338 3667 -5306
rect 3633 -5408 3667 -5376
rect 3633 -5410 3667 -5408
rect 3891 -5306 3925 -5304
rect 3891 -5338 3925 -5306
rect 3891 -5408 3925 -5376
rect 3891 -5410 3925 -5408
rect 4149 -5306 4183 -5304
rect 4149 -5338 4183 -5306
rect 4149 -5408 4183 -5376
rect 4149 -5410 4183 -5408
rect 4407 -5306 4441 -5304
rect 4407 -5338 4441 -5306
rect 4407 -5408 4441 -5376
rect 4407 -5410 4441 -5408
rect 4665 -5306 4699 -5304
rect 4665 -5338 4699 -5306
rect 4665 -5408 4699 -5376
rect 4665 -5410 4699 -5408
rect 4859 -5306 4893 -5304
rect 4859 -5338 4893 -5306
rect 4859 -5408 4893 -5376
rect 4859 -5410 4893 -5408
rect 5117 -5306 5151 -5304
rect 5117 -5338 5151 -5306
rect 5117 -5408 5151 -5376
rect 5117 -5410 5151 -5408
rect 5231 -5321 5265 -5287
rect 5231 -5389 5265 -5359
rect 5231 -5393 5265 -5389
rect 872 -5525 906 -5503
rect 5231 -5457 5265 -5431
rect 5231 -5465 5265 -5457
rect 5345 -5306 5379 -5304
rect 5345 -5338 5379 -5306
rect 5345 -5408 5379 -5376
rect 5345 -5410 5379 -5408
rect 5603 -5306 5637 -5304
rect 5603 -5338 5637 -5306
rect 5603 -5408 5637 -5376
rect 5603 -5410 5637 -5408
rect 5796 -5306 5830 -5304
rect 5796 -5338 5830 -5306
rect 5796 -5408 5830 -5376
rect 5796 -5410 5830 -5408
rect 6054 -5306 6088 -5304
rect 6054 -5338 6088 -5306
rect 6054 -5408 6088 -5376
rect 6054 -5410 6088 -5408
rect 6312 -5306 6346 -5304
rect 6312 -5338 6346 -5306
rect 6312 -5408 6346 -5376
rect 6312 -5410 6346 -5408
rect 6570 -5306 6604 -5304
rect 6570 -5338 6604 -5306
rect 6570 -5408 6604 -5376
rect 6570 -5410 6604 -5408
rect 6828 -5306 6862 -5304
rect 6828 -5338 6862 -5306
rect 6828 -5408 6862 -5376
rect 6828 -5410 6862 -5408
rect 7022 -5306 7056 -5304
rect 7022 -5338 7056 -5306
rect 7022 -5408 7056 -5376
rect 7022 -5410 7056 -5408
rect 7280 -5306 7314 -5304
rect 7280 -5338 7314 -5306
rect 7280 -5408 7314 -5376
rect 7280 -5410 7314 -5408
rect 7538 -5306 7572 -5304
rect 7538 -5338 7572 -5306
rect 7538 -5408 7572 -5376
rect 7538 -5410 7572 -5408
rect 7796 -5306 7830 -5304
rect 7796 -5338 7830 -5306
rect 7796 -5408 7830 -5376
rect 7796 -5410 7830 -5408
rect 7990 -5306 8024 -5304
rect 7990 -5338 8024 -5306
rect 7990 -5408 8024 -5376
rect 7990 -5410 8024 -5408
rect 8248 -5306 8282 -5304
rect 8248 -5338 8282 -5306
rect 8248 -5408 8282 -5376
rect 8248 -5410 8282 -5408
rect 8506 -5306 8540 -5304
rect 8506 -5338 8540 -5306
rect 8506 -5408 8540 -5376
rect 8506 -5410 8540 -5408
rect 8764 -5306 8798 -5304
rect 8764 -5338 8798 -5306
rect 8764 -5408 8798 -5376
rect 8764 -5410 8798 -5408
rect 9022 -5306 9056 -5304
rect 9022 -5338 9056 -5306
rect 9022 -5408 9056 -5376
rect 9022 -5410 9056 -5408
rect 9216 -5306 9250 -5304
rect 9216 -5338 9250 -5306
rect 9216 -5408 9250 -5376
rect 9216 -5410 9250 -5408
rect 9474 -5306 9508 -5304
rect 9474 -5338 9508 -5306
rect 9474 -5408 9508 -5376
rect 9474 -5410 9508 -5408
rect 9589 -5321 9623 -5287
rect 9589 -5389 9623 -5359
rect 9589 -5393 9623 -5389
rect 9589 -5457 9623 -5431
rect 872 -5537 906 -5525
rect 1080 -5538 1082 -5504
rect 1082 -5538 1114 -5504
rect 1152 -5538 1184 -5504
rect 1184 -5538 1186 -5504
rect 1532 -5538 1534 -5504
rect 1534 -5538 1566 -5504
rect 1604 -5538 1636 -5504
rect 1636 -5538 1638 -5504
rect 1790 -5538 1792 -5504
rect 1792 -5538 1824 -5504
rect 1862 -5538 1894 -5504
rect 1894 -5538 1896 -5504
rect 2048 -5538 2050 -5504
rect 2050 -5538 2082 -5504
rect 2120 -5538 2152 -5504
rect 2152 -5538 2154 -5504
rect 2306 -5538 2308 -5504
rect 2308 -5538 2340 -5504
rect 2378 -5538 2410 -5504
rect 2410 -5538 2412 -5504
rect 2758 -5538 2760 -5504
rect 2760 -5538 2792 -5504
rect 2830 -5538 2862 -5504
rect 2862 -5538 2864 -5504
rect 3016 -5538 3018 -5504
rect 3018 -5538 3050 -5504
rect 3088 -5538 3120 -5504
rect 3120 -5538 3122 -5504
rect 3274 -5538 3276 -5504
rect 3276 -5538 3308 -5504
rect 3346 -5538 3378 -5504
rect 3378 -5538 3380 -5504
rect 3726 -5538 3728 -5504
rect 3728 -5538 3760 -5504
rect 3798 -5538 3830 -5504
rect 3830 -5538 3832 -5504
rect 3984 -5538 3986 -5504
rect 3986 -5538 4018 -5504
rect 4056 -5538 4088 -5504
rect 4088 -5538 4090 -5504
rect 4242 -5538 4244 -5504
rect 4244 -5538 4276 -5504
rect 4314 -5538 4346 -5504
rect 4346 -5538 4348 -5504
rect 4500 -5538 4502 -5504
rect 4502 -5538 4534 -5504
rect 4572 -5538 4604 -5504
rect 4604 -5538 4606 -5504
rect 4952 -5538 4954 -5504
rect 4954 -5538 4986 -5504
rect 5024 -5538 5056 -5504
rect 5056 -5538 5058 -5504
rect 5231 -5525 5265 -5503
rect 9589 -5465 9623 -5457
rect 5231 -5537 5265 -5525
rect 872 -5593 906 -5575
rect 872 -5609 906 -5593
rect 872 -5661 906 -5647
rect 872 -5681 906 -5661
rect 872 -5729 906 -5719
rect 872 -5753 906 -5729
rect 872 -5797 906 -5791
rect 872 -5825 906 -5797
rect 872 -5865 906 -5863
rect 872 -5897 906 -5865
rect 5438 -5538 5440 -5504
rect 5440 -5538 5472 -5504
rect 5510 -5538 5542 -5504
rect 5542 -5538 5544 -5504
rect 5889 -5538 5891 -5504
rect 5891 -5538 5923 -5504
rect 5961 -5538 5993 -5504
rect 5993 -5538 5995 -5504
rect 6147 -5538 6149 -5504
rect 6149 -5538 6181 -5504
rect 6219 -5538 6251 -5504
rect 6251 -5538 6253 -5504
rect 6405 -5538 6407 -5504
rect 6407 -5538 6439 -5504
rect 6477 -5538 6509 -5504
rect 6509 -5538 6511 -5504
rect 6663 -5538 6665 -5504
rect 6665 -5538 6697 -5504
rect 6735 -5538 6767 -5504
rect 6767 -5538 6769 -5504
rect 7115 -5538 7117 -5504
rect 7117 -5538 7149 -5504
rect 7187 -5538 7219 -5504
rect 7219 -5538 7221 -5504
rect 7373 -5538 7375 -5504
rect 7375 -5538 7407 -5504
rect 7445 -5538 7477 -5504
rect 7477 -5538 7479 -5504
rect 7631 -5538 7633 -5504
rect 7633 -5538 7665 -5504
rect 7703 -5538 7735 -5504
rect 7735 -5538 7737 -5504
rect 8083 -5538 8085 -5504
rect 8085 -5538 8117 -5504
rect 8155 -5538 8187 -5504
rect 8187 -5538 8189 -5504
rect 8341 -5538 8343 -5504
rect 8343 -5538 8375 -5504
rect 8413 -5538 8445 -5504
rect 8445 -5538 8447 -5504
rect 8599 -5538 8601 -5504
rect 8601 -5538 8633 -5504
rect 8671 -5538 8703 -5504
rect 8703 -5538 8705 -5504
rect 8857 -5538 8859 -5504
rect 8859 -5538 8891 -5504
rect 8929 -5538 8961 -5504
rect 8961 -5538 8963 -5504
rect 9309 -5538 9311 -5504
rect 9311 -5538 9343 -5504
rect 9381 -5538 9413 -5504
rect 9413 -5538 9415 -5504
rect 9589 -5525 9623 -5503
rect 9589 -5537 9623 -5525
rect 5231 -5593 5265 -5575
rect 5231 -5609 5265 -5593
rect 5231 -5661 5265 -5647
rect 5231 -5681 5265 -5661
rect 5231 -5729 5265 -5719
rect 5231 -5753 5265 -5729
rect 5231 -5797 5265 -5791
rect 5231 -5825 5265 -5797
rect 1080 -5900 1082 -5866
rect 1082 -5900 1114 -5866
rect 1152 -5900 1184 -5866
rect 1184 -5900 1186 -5866
rect 1532 -5900 1534 -5866
rect 1534 -5900 1566 -5866
rect 1604 -5900 1636 -5866
rect 1636 -5900 1638 -5866
rect 1790 -5900 1792 -5866
rect 1792 -5900 1824 -5866
rect 1862 -5900 1894 -5866
rect 1894 -5900 1896 -5866
rect 2048 -5900 2050 -5866
rect 2050 -5900 2082 -5866
rect 2120 -5900 2152 -5866
rect 2152 -5900 2154 -5866
rect 2306 -5900 2308 -5866
rect 2308 -5900 2340 -5866
rect 2378 -5900 2410 -5866
rect 2410 -5900 2412 -5866
rect 2758 -5900 2760 -5866
rect 2760 -5900 2792 -5866
rect 2830 -5900 2862 -5866
rect 2862 -5900 2864 -5866
rect 3016 -5900 3018 -5866
rect 3018 -5900 3050 -5866
rect 3088 -5900 3120 -5866
rect 3120 -5900 3122 -5866
rect 3274 -5900 3276 -5866
rect 3276 -5900 3308 -5866
rect 3346 -5900 3378 -5866
rect 3378 -5900 3380 -5866
rect 3726 -5900 3728 -5866
rect 3728 -5900 3760 -5866
rect 3798 -5900 3830 -5866
rect 3830 -5900 3832 -5866
rect 3984 -5900 3986 -5866
rect 3986 -5900 4018 -5866
rect 4056 -5900 4088 -5866
rect 4088 -5900 4090 -5866
rect 4242 -5900 4244 -5866
rect 4244 -5900 4276 -5866
rect 4314 -5900 4346 -5866
rect 4346 -5900 4348 -5866
rect 4500 -5900 4502 -5866
rect 4502 -5900 4534 -5866
rect 4572 -5900 4604 -5866
rect 4604 -5900 4606 -5866
rect 4952 -5900 4954 -5866
rect 4954 -5900 4986 -5866
rect 5024 -5900 5056 -5866
rect 5056 -5900 5058 -5866
rect 5231 -5865 5265 -5863
rect 5231 -5897 5265 -5865
rect 9589 -5593 9623 -5575
rect 9589 -5609 9623 -5593
rect 9589 -5661 9623 -5647
rect 9589 -5681 9623 -5661
rect 9589 -5729 9623 -5719
rect 9589 -5753 9623 -5729
rect 9589 -5797 9623 -5791
rect 9589 -5825 9623 -5797
rect 9589 -5865 9623 -5863
rect 872 -5967 906 -5935
rect 5438 -5900 5440 -5866
rect 5440 -5900 5472 -5866
rect 5510 -5900 5542 -5866
rect 5542 -5900 5544 -5866
rect 5889 -5900 5891 -5866
rect 5891 -5900 5923 -5866
rect 5961 -5900 5993 -5866
rect 5993 -5900 5995 -5866
rect 6147 -5900 6149 -5866
rect 6149 -5900 6181 -5866
rect 6219 -5900 6251 -5866
rect 6251 -5900 6253 -5866
rect 6405 -5900 6407 -5866
rect 6407 -5900 6439 -5866
rect 6477 -5900 6509 -5866
rect 6509 -5900 6511 -5866
rect 6663 -5900 6665 -5866
rect 6665 -5900 6697 -5866
rect 6735 -5900 6767 -5866
rect 6767 -5900 6769 -5866
rect 7115 -5900 7117 -5866
rect 7117 -5900 7149 -5866
rect 7187 -5900 7219 -5866
rect 7219 -5900 7221 -5866
rect 7373 -5900 7375 -5866
rect 7375 -5900 7407 -5866
rect 7445 -5900 7477 -5866
rect 7477 -5900 7479 -5866
rect 7631 -5900 7633 -5866
rect 7633 -5900 7665 -5866
rect 7703 -5900 7735 -5866
rect 7735 -5900 7737 -5866
rect 8083 -5900 8085 -5866
rect 8085 -5900 8117 -5866
rect 8155 -5900 8187 -5866
rect 8187 -5900 8189 -5866
rect 8341 -5900 8343 -5866
rect 8343 -5900 8375 -5866
rect 8413 -5900 8445 -5866
rect 8445 -5900 8447 -5866
rect 8599 -5900 8601 -5866
rect 8601 -5900 8633 -5866
rect 8671 -5900 8703 -5866
rect 8703 -5900 8705 -5866
rect 8857 -5900 8859 -5866
rect 8859 -5900 8891 -5866
rect 8929 -5900 8961 -5866
rect 8961 -5900 8963 -5866
rect 9309 -5900 9311 -5866
rect 9311 -5900 9343 -5866
rect 9381 -5900 9413 -5866
rect 9413 -5900 9415 -5866
rect 9589 -5897 9623 -5865
rect 872 -5969 906 -5967
rect 872 -6035 906 -6007
rect 872 -6041 906 -6035
rect 872 -6103 906 -6079
rect 872 -6113 906 -6103
rect 987 -5996 1021 -5994
rect 987 -6028 1021 -5996
rect 987 -6098 1021 -6066
rect 987 -6100 1021 -6098
rect 1245 -5996 1279 -5994
rect 1245 -6028 1279 -5996
rect 1245 -6098 1279 -6066
rect 1245 -6100 1279 -6098
rect 1439 -5996 1473 -5994
rect 1439 -6028 1473 -5996
rect 1439 -6098 1473 -6066
rect 1439 -6100 1473 -6098
rect 1697 -5996 1731 -5994
rect 1697 -6028 1731 -5996
rect 1697 -6098 1731 -6066
rect 1697 -6100 1731 -6098
rect 1955 -5996 1989 -5994
rect 1955 -6028 1989 -5996
rect 1955 -6098 1989 -6066
rect 1955 -6100 1989 -6098
rect 2213 -5996 2247 -5994
rect 2213 -6028 2247 -5996
rect 2213 -6098 2247 -6066
rect 2213 -6100 2247 -6098
rect 2471 -5996 2505 -5994
rect 2471 -6028 2505 -5996
rect 2471 -6098 2505 -6066
rect 2471 -6100 2505 -6098
rect 2665 -5996 2699 -5994
rect 2665 -6028 2699 -5996
rect 2665 -6098 2699 -6066
rect 2665 -6100 2699 -6098
rect 2923 -5996 2957 -5994
rect 2923 -6028 2957 -5996
rect 2923 -6098 2957 -6066
rect 2923 -6100 2957 -6098
rect 3181 -5996 3215 -5994
rect 3181 -6028 3215 -5996
rect 3181 -6098 3215 -6066
rect 3181 -6100 3215 -6098
rect 3439 -5996 3473 -5994
rect 3439 -6028 3473 -5996
rect 3439 -6098 3473 -6066
rect 3439 -6100 3473 -6098
rect 3633 -5996 3667 -5994
rect 3633 -6028 3667 -5996
rect 3633 -6098 3667 -6066
rect 3633 -6100 3667 -6098
rect 3891 -5996 3925 -5994
rect 3891 -6028 3925 -5996
rect 3891 -6098 3925 -6066
rect 3891 -6100 3925 -6098
rect 4149 -5996 4183 -5994
rect 4149 -6028 4183 -5996
rect 4149 -6098 4183 -6066
rect 4149 -6100 4183 -6098
rect 4407 -5996 4441 -5994
rect 4407 -6028 4441 -5996
rect 4407 -6098 4441 -6066
rect 4407 -6100 4441 -6098
rect 4665 -5996 4699 -5994
rect 4665 -6028 4699 -5996
rect 4665 -6098 4699 -6066
rect 4665 -6100 4699 -6098
rect 4859 -5996 4893 -5994
rect 4859 -6028 4893 -5996
rect 4859 -6098 4893 -6066
rect 4859 -6100 4893 -6098
rect 5117 -5996 5151 -5994
rect 5117 -6028 5151 -5996
rect 5117 -6098 5151 -6066
rect 5117 -6100 5151 -6098
rect 5231 -5967 5265 -5935
rect 5231 -5969 5265 -5967
rect 5231 -6035 5265 -6007
rect 5231 -6041 5265 -6035
rect 5231 -6103 5265 -6079
rect 5231 -6113 5265 -6103
rect 5345 -5996 5379 -5994
rect 5345 -6028 5379 -5996
rect 5345 -6098 5379 -6066
rect 5345 -6100 5379 -6098
rect 5603 -5996 5637 -5994
rect 5603 -6028 5637 -5996
rect 5603 -6098 5637 -6066
rect 5603 -6100 5637 -6098
rect 5796 -5996 5830 -5994
rect 5796 -6028 5830 -5996
rect 5796 -6098 5830 -6066
rect 5796 -6100 5830 -6098
rect 6054 -5996 6088 -5994
rect 6054 -6028 6088 -5996
rect 6054 -6098 6088 -6066
rect 6054 -6100 6088 -6098
rect 6312 -5996 6346 -5994
rect 6312 -6028 6346 -5996
rect 6312 -6098 6346 -6066
rect 6312 -6100 6346 -6098
rect 6570 -5996 6604 -5994
rect 6570 -6028 6604 -5996
rect 6570 -6098 6604 -6066
rect 6570 -6100 6604 -6098
rect 6828 -5996 6862 -5994
rect 6828 -6028 6862 -5996
rect 6828 -6098 6862 -6066
rect 6828 -6100 6862 -6098
rect 7022 -5996 7056 -5994
rect 7022 -6028 7056 -5996
rect 7022 -6098 7056 -6066
rect 7022 -6100 7056 -6098
rect 7280 -5996 7314 -5994
rect 7280 -6028 7314 -5996
rect 7280 -6098 7314 -6066
rect 7280 -6100 7314 -6098
rect 7538 -5996 7572 -5994
rect 7538 -6028 7572 -5996
rect 7538 -6098 7572 -6066
rect 7538 -6100 7572 -6098
rect 7796 -5996 7830 -5994
rect 7796 -6028 7830 -5996
rect 7796 -6098 7830 -6066
rect 7796 -6100 7830 -6098
rect 7990 -5996 8024 -5994
rect 7990 -6028 8024 -5996
rect 7990 -6098 8024 -6066
rect 7990 -6100 8024 -6098
rect 8248 -5996 8282 -5994
rect 8248 -6028 8282 -5996
rect 8248 -6098 8282 -6066
rect 8248 -6100 8282 -6098
rect 8506 -5996 8540 -5994
rect 8506 -6028 8540 -5996
rect 8506 -6098 8540 -6066
rect 8506 -6100 8540 -6098
rect 8764 -5996 8798 -5994
rect 8764 -6028 8798 -5996
rect 8764 -6098 8798 -6066
rect 8764 -6100 8798 -6098
rect 9022 -5996 9056 -5994
rect 9022 -6028 9056 -5996
rect 9022 -6098 9056 -6066
rect 9022 -6100 9056 -6098
rect 9216 -5996 9250 -5994
rect 9216 -6028 9250 -5996
rect 9216 -6098 9250 -6066
rect 9216 -6100 9250 -6098
rect 9474 -5996 9508 -5994
rect 9474 -6028 9508 -5996
rect 9474 -6098 9508 -6066
rect 9474 -6100 9508 -6098
rect 9589 -5967 9623 -5935
rect 9589 -5969 9623 -5967
rect 9589 -6035 9623 -6007
rect 9589 -6041 9623 -6035
rect 9589 -6103 9623 -6079
rect 9589 -6113 9623 -6103
rect 872 -6171 906 -6151
rect 872 -6185 906 -6171
rect 872 -6239 906 -6223
rect 872 -6257 906 -6239
rect 872 -6307 906 -6295
rect 872 -6329 906 -6307
rect 872 -6375 906 -6367
rect 872 -6401 906 -6375
rect 872 -6473 906 -6439
rect 5231 -6171 5265 -6151
rect 5231 -6185 5265 -6171
rect 5231 -6239 5265 -6223
rect 5231 -6257 5265 -6239
rect 5231 -6307 5265 -6295
rect 5231 -6329 5265 -6307
rect 5231 -6375 5265 -6367
rect 5231 -6401 5265 -6375
rect 5231 -6473 5265 -6439
rect 9589 -6171 9623 -6151
rect 9589 -6185 9623 -6171
rect 9589 -6239 9623 -6223
rect 9589 -6257 9623 -6239
rect 9589 -6307 9623 -6295
rect 9589 -6329 9623 -6307
rect 9589 -6375 9623 -6367
rect 9589 -6401 9623 -6375
rect 9589 -6473 9623 -6439
rect 872 -6545 906 -6511
rect 5231 -6545 5265 -6511
rect 9589 -6545 9623 -6511
rect 872 -6617 906 -6583
rect 872 -6681 906 -6655
rect 872 -6689 906 -6681
rect 872 -6749 906 -6727
rect 872 -6761 906 -6749
rect 872 -6817 906 -6799
rect 872 -6833 906 -6817
rect 872 -6885 906 -6871
rect 872 -6905 906 -6885
rect 5231 -6617 5265 -6583
rect 5231 -6681 5265 -6655
rect 5231 -6689 5265 -6681
rect 5231 -6749 5265 -6727
rect 5231 -6761 5265 -6749
rect 5231 -6817 5265 -6799
rect 5231 -6833 5265 -6817
rect 872 -6953 906 -6943
rect 872 -6977 906 -6953
rect 872 -7021 906 -7015
rect 872 -7049 906 -7021
rect 872 -7089 906 -7087
rect 872 -7121 906 -7089
rect 987 -6953 1021 -6951
rect 987 -6985 1021 -6953
rect 987 -7055 1021 -7023
rect 987 -7057 1021 -7055
rect 1245 -6953 1279 -6951
rect 1245 -6985 1279 -6953
rect 1245 -7055 1279 -7023
rect 1245 -7057 1279 -7055
rect 1439 -6953 1473 -6951
rect 1439 -6985 1473 -6953
rect 1439 -7055 1473 -7023
rect 1439 -7057 1473 -7055
rect 1697 -6953 1731 -6951
rect 1697 -6985 1731 -6953
rect 1697 -7055 1731 -7023
rect 1697 -7057 1731 -7055
rect 1955 -6953 1989 -6951
rect 1955 -6985 1989 -6953
rect 1955 -7055 1989 -7023
rect 1955 -7057 1989 -7055
rect 2213 -6953 2247 -6951
rect 2213 -6985 2247 -6953
rect 2213 -7055 2247 -7023
rect 2213 -7057 2247 -7055
rect 2471 -6953 2505 -6951
rect 2471 -6985 2505 -6953
rect 2471 -7055 2505 -7023
rect 2471 -7057 2505 -7055
rect 2665 -6953 2699 -6951
rect 2665 -6985 2699 -6953
rect 2665 -7055 2699 -7023
rect 2665 -7057 2699 -7055
rect 2923 -6953 2957 -6951
rect 2923 -6985 2957 -6953
rect 2923 -7055 2957 -7023
rect 2923 -7057 2957 -7055
rect 3181 -6953 3215 -6951
rect 3181 -6985 3215 -6953
rect 3181 -7055 3215 -7023
rect 3181 -7057 3215 -7055
rect 3439 -6953 3473 -6951
rect 3439 -6985 3473 -6953
rect 3439 -7055 3473 -7023
rect 3439 -7057 3473 -7055
rect 3633 -6953 3667 -6951
rect 3633 -6985 3667 -6953
rect 3633 -7055 3667 -7023
rect 3633 -7057 3667 -7055
rect 3891 -6953 3925 -6951
rect 3891 -6985 3925 -6953
rect 3891 -7055 3925 -7023
rect 3891 -7057 3925 -7055
rect 4149 -6953 4183 -6951
rect 4149 -6985 4183 -6953
rect 4149 -7055 4183 -7023
rect 4149 -7057 4183 -7055
rect 4407 -6953 4441 -6951
rect 4407 -6985 4441 -6953
rect 4407 -7055 4441 -7023
rect 4407 -7057 4441 -7055
rect 4665 -6953 4699 -6951
rect 4665 -6985 4699 -6953
rect 4665 -7055 4699 -7023
rect 4665 -7057 4699 -7055
rect 4859 -6953 4893 -6951
rect 4859 -6985 4893 -6953
rect 4859 -7055 4893 -7023
rect 4859 -7057 4893 -7055
rect 5117 -6953 5151 -6951
rect 5117 -6985 5151 -6953
rect 5117 -7055 5151 -7023
rect 5117 -7057 5151 -7055
rect 5231 -6885 5265 -6871
rect 5231 -6905 5265 -6885
rect 9589 -6617 9623 -6583
rect 9589 -6681 9623 -6655
rect 9589 -6689 9623 -6681
rect 9589 -6749 9623 -6727
rect 9589 -6761 9623 -6749
rect 9589 -6817 9623 -6799
rect 9589 -6833 9623 -6817
rect 9589 -6885 9623 -6871
rect 5231 -6953 5265 -6943
rect 5231 -6977 5265 -6953
rect 5231 -7021 5265 -7015
rect 5231 -7049 5265 -7021
rect 5231 -7089 5265 -7087
rect 5231 -7121 5265 -7089
rect 5345 -6953 5379 -6951
rect 5345 -6985 5379 -6953
rect 5345 -7055 5379 -7023
rect 5345 -7057 5379 -7055
rect 5603 -6953 5637 -6951
rect 5603 -6985 5637 -6953
rect 5603 -7055 5637 -7023
rect 5603 -7057 5637 -7055
rect 5796 -6953 5830 -6951
rect 5796 -6985 5830 -6953
rect 5796 -7055 5830 -7023
rect 5796 -7057 5830 -7055
rect 6054 -6953 6088 -6951
rect 6054 -6985 6088 -6953
rect 6054 -7055 6088 -7023
rect 6054 -7057 6088 -7055
rect 6312 -6953 6346 -6951
rect 6312 -6985 6346 -6953
rect 6312 -7055 6346 -7023
rect 6312 -7057 6346 -7055
rect 6570 -6953 6604 -6951
rect 6570 -6985 6604 -6953
rect 6570 -7055 6604 -7023
rect 6570 -7057 6604 -7055
rect 6828 -6953 6862 -6951
rect 6828 -6985 6862 -6953
rect 6828 -7055 6862 -7023
rect 6828 -7057 6862 -7055
rect 7022 -6953 7056 -6951
rect 7022 -6985 7056 -6953
rect 7022 -7055 7056 -7023
rect 7022 -7057 7056 -7055
rect 7280 -6953 7314 -6951
rect 7280 -6985 7314 -6953
rect 7280 -7055 7314 -7023
rect 7280 -7057 7314 -7055
rect 7538 -6953 7572 -6951
rect 7538 -6985 7572 -6953
rect 7538 -7055 7572 -7023
rect 7538 -7057 7572 -7055
rect 7796 -6953 7830 -6951
rect 7796 -6985 7830 -6953
rect 7796 -7055 7830 -7023
rect 7796 -7057 7830 -7055
rect 7990 -6953 8024 -6951
rect 7990 -6985 8024 -6953
rect 7990 -7055 8024 -7023
rect 7990 -7057 8024 -7055
rect 8248 -6953 8282 -6951
rect 8248 -6985 8282 -6953
rect 8248 -7055 8282 -7023
rect 8248 -7057 8282 -7055
rect 8506 -6953 8540 -6951
rect 8506 -6985 8540 -6953
rect 8506 -7055 8540 -7023
rect 8506 -7057 8540 -7055
rect 8764 -6953 8798 -6951
rect 8764 -6985 8798 -6953
rect 8764 -7055 8798 -7023
rect 8764 -7057 8798 -7055
rect 9022 -6953 9056 -6951
rect 9022 -6985 9056 -6953
rect 9022 -7055 9056 -7023
rect 9022 -7057 9056 -7055
rect 9216 -6953 9250 -6951
rect 9216 -6985 9250 -6953
rect 9216 -7055 9250 -7023
rect 9216 -7057 9250 -7055
rect 9474 -6953 9508 -6951
rect 9474 -6985 9508 -6953
rect 9474 -7055 9508 -7023
rect 9474 -7057 9508 -7055
rect 9589 -6905 9623 -6885
rect 9589 -6953 9623 -6943
rect 9589 -6977 9623 -6953
rect 9589 -7021 9623 -7015
rect 9589 -7049 9623 -7021
rect 9589 -7089 9623 -7087
rect 872 -7191 906 -7159
rect 1080 -7185 1082 -7151
rect 1082 -7185 1114 -7151
rect 1152 -7185 1184 -7151
rect 1184 -7185 1186 -7151
rect 1532 -7185 1534 -7151
rect 1534 -7185 1566 -7151
rect 1604 -7185 1636 -7151
rect 1636 -7185 1638 -7151
rect 1790 -7185 1792 -7151
rect 1792 -7185 1824 -7151
rect 1862 -7185 1894 -7151
rect 1894 -7185 1896 -7151
rect 2048 -7185 2050 -7151
rect 2050 -7185 2082 -7151
rect 2120 -7185 2152 -7151
rect 2152 -7185 2154 -7151
rect 2306 -7185 2308 -7151
rect 2308 -7185 2340 -7151
rect 2378 -7185 2410 -7151
rect 2410 -7185 2412 -7151
rect 2758 -7185 2760 -7151
rect 2760 -7185 2792 -7151
rect 2830 -7185 2862 -7151
rect 2862 -7185 2864 -7151
rect 3016 -7185 3018 -7151
rect 3018 -7185 3050 -7151
rect 3088 -7185 3120 -7151
rect 3120 -7185 3122 -7151
rect 3274 -7185 3276 -7151
rect 3276 -7185 3308 -7151
rect 3346 -7185 3378 -7151
rect 3378 -7185 3380 -7151
rect 3726 -7185 3728 -7151
rect 3728 -7185 3760 -7151
rect 3798 -7185 3830 -7151
rect 3830 -7185 3832 -7151
rect 3984 -7185 3986 -7151
rect 3986 -7185 4018 -7151
rect 4056 -7185 4088 -7151
rect 4088 -7185 4090 -7151
rect 4242 -7185 4244 -7151
rect 4244 -7185 4276 -7151
rect 4314 -7185 4346 -7151
rect 4346 -7185 4348 -7151
rect 4500 -7185 4502 -7151
rect 4502 -7185 4534 -7151
rect 4572 -7185 4604 -7151
rect 4604 -7185 4606 -7151
rect 4952 -7185 4954 -7151
rect 4954 -7185 4986 -7151
rect 5024 -7185 5056 -7151
rect 5056 -7185 5058 -7151
rect 9589 -7121 9623 -7089
rect 872 -7193 906 -7191
rect 872 -7259 906 -7231
rect 872 -7265 906 -7259
rect 872 -7327 906 -7303
rect 872 -7337 906 -7327
rect 872 -7395 906 -7375
rect 872 -7409 906 -7395
rect 872 -7463 906 -7447
rect 872 -7481 906 -7463
rect 5231 -7191 5265 -7159
rect 5438 -7185 5440 -7151
rect 5440 -7185 5472 -7151
rect 5510 -7185 5542 -7151
rect 5542 -7185 5544 -7151
rect 5889 -7185 5891 -7151
rect 5891 -7185 5923 -7151
rect 5961 -7185 5993 -7151
rect 5993 -7185 5995 -7151
rect 6147 -7185 6149 -7151
rect 6149 -7185 6181 -7151
rect 6219 -7185 6251 -7151
rect 6251 -7185 6253 -7151
rect 6405 -7185 6407 -7151
rect 6407 -7185 6439 -7151
rect 6477 -7185 6509 -7151
rect 6509 -7185 6511 -7151
rect 6663 -7185 6665 -7151
rect 6665 -7185 6697 -7151
rect 6735 -7185 6767 -7151
rect 6767 -7185 6769 -7151
rect 7115 -7185 7117 -7151
rect 7117 -7185 7149 -7151
rect 7187 -7185 7219 -7151
rect 7219 -7185 7221 -7151
rect 7373 -7185 7375 -7151
rect 7375 -7185 7407 -7151
rect 7445 -7185 7477 -7151
rect 7477 -7185 7479 -7151
rect 7631 -7185 7633 -7151
rect 7633 -7185 7665 -7151
rect 7703 -7185 7735 -7151
rect 7735 -7185 7737 -7151
rect 8083 -7185 8085 -7151
rect 8085 -7185 8117 -7151
rect 8155 -7185 8187 -7151
rect 8187 -7185 8189 -7151
rect 8341 -7185 8343 -7151
rect 8343 -7185 8375 -7151
rect 8413 -7185 8445 -7151
rect 8445 -7185 8447 -7151
rect 8599 -7185 8601 -7151
rect 8601 -7185 8633 -7151
rect 8671 -7185 8703 -7151
rect 8703 -7185 8705 -7151
rect 8857 -7185 8859 -7151
rect 8859 -7185 8891 -7151
rect 8929 -7185 8961 -7151
rect 8961 -7185 8963 -7151
rect 9309 -7185 9311 -7151
rect 9311 -7185 9343 -7151
rect 9381 -7185 9413 -7151
rect 9413 -7185 9415 -7151
rect 5231 -7193 5265 -7191
rect 5231 -7259 5265 -7231
rect 5231 -7265 5265 -7259
rect 5231 -7327 5265 -7303
rect 5231 -7337 5265 -7327
rect 5231 -7395 5265 -7375
rect 5231 -7409 5265 -7395
rect 5231 -7463 5265 -7447
rect 5231 -7481 5265 -7463
rect 872 -7531 906 -7519
rect 872 -7553 906 -7531
rect 1080 -7547 1082 -7513
rect 1082 -7547 1114 -7513
rect 1152 -7547 1184 -7513
rect 1184 -7547 1186 -7513
rect 1532 -7547 1534 -7513
rect 1534 -7547 1566 -7513
rect 1604 -7547 1636 -7513
rect 1636 -7547 1638 -7513
rect 1790 -7547 1792 -7513
rect 1792 -7547 1824 -7513
rect 1862 -7547 1894 -7513
rect 1894 -7547 1896 -7513
rect 2048 -7547 2050 -7513
rect 2050 -7547 2082 -7513
rect 2120 -7547 2152 -7513
rect 2152 -7547 2154 -7513
rect 2306 -7547 2308 -7513
rect 2308 -7547 2340 -7513
rect 2378 -7547 2410 -7513
rect 2410 -7547 2412 -7513
rect 2758 -7547 2760 -7513
rect 2760 -7547 2792 -7513
rect 2830 -7547 2862 -7513
rect 2862 -7547 2864 -7513
rect 3016 -7547 3018 -7513
rect 3018 -7547 3050 -7513
rect 3088 -7547 3120 -7513
rect 3120 -7547 3122 -7513
rect 3274 -7547 3276 -7513
rect 3276 -7547 3308 -7513
rect 3346 -7547 3378 -7513
rect 3378 -7547 3380 -7513
rect 3726 -7547 3728 -7513
rect 3728 -7547 3760 -7513
rect 3798 -7547 3830 -7513
rect 3830 -7547 3832 -7513
rect 3984 -7547 3986 -7513
rect 3986 -7547 4018 -7513
rect 4056 -7547 4088 -7513
rect 4088 -7547 4090 -7513
rect 4242 -7547 4244 -7513
rect 4244 -7547 4276 -7513
rect 4314 -7547 4346 -7513
rect 4346 -7547 4348 -7513
rect 4500 -7547 4502 -7513
rect 4502 -7547 4534 -7513
rect 4572 -7547 4604 -7513
rect 4604 -7547 4606 -7513
rect 4952 -7547 4954 -7513
rect 4954 -7547 4986 -7513
rect 5024 -7547 5056 -7513
rect 5056 -7547 5058 -7513
rect 9589 -7191 9623 -7159
rect 9589 -7193 9623 -7191
rect 9589 -7259 9623 -7231
rect 9589 -7265 9623 -7259
rect 9589 -7327 9623 -7303
rect 9589 -7337 9623 -7327
rect 9589 -7395 9623 -7375
rect 9589 -7409 9623 -7395
rect 9589 -7463 9623 -7447
rect 9589 -7481 9623 -7463
rect 5231 -7531 5265 -7519
rect 5231 -7553 5265 -7531
rect 5438 -7547 5440 -7513
rect 5440 -7547 5472 -7513
rect 5510 -7547 5542 -7513
rect 5542 -7547 5544 -7513
rect 5889 -7547 5891 -7513
rect 5891 -7547 5923 -7513
rect 5961 -7547 5993 -7513
rect 5993 -7547 5995 -7513
rect 6147 -7547 6149 -7513
rect 6149 -7547 6181 -7513
rect 6219 -7547 6251 -7513
rect 6251 -7547 6253 -7513
rect 6405 -7547 6407 -7513
rect 6407 -7547 6439 -7513
rect 6477 -7547 6509 -7513
rect 6509 -7547 6511 -7513
rect 6663 -7547 6665 -7513
rect 6665 -7547 6697 -7513
rect 6735 -7547 6767 -7513
rect 6767 -7547 6769 -7513
rect 7115 -7547 7117 -7513
rect 7117 -7547 7149 -7513
rect 7187 -7547 7219 -7513
rect 7219 -7547 7221 -7513
rect 7373 -7547 7375 -7513
rect 7375 -7547 7407 -7513
rect 7445 -7547 7477 -7513
rect 7477 -7547 7479 -7513
rect 7631 -7547 7633 -7513
rect 7633 -7547 7665 -7513
rect 7703 -7547 7735 -7513
rect 7735 -7547 7737 -7513
rect 8083 -7547 8085 -7513
rect 8085 -7547 8117 -7513
rect 8155 -7547 8187 -7513
rect 8187 -7547 8189 -7513
rect 8341 -7547 8343 -7513
rect 8343 -7547 8375 -7513
rect 8413 -7547 8445 -7513
rect 8445 -7547 8447 -7513
rect 8599 -7547 8601 -7513
rect 8601 -7547 8633 -7513
rect 8671 -7547 8703 -7513
rect 8703 -7547 8705 -7513
rect 8857 -7547 8859 -7513
rect 8859 -7547 8891 -7513
rect 8929 -7547 8961 -7513
rect 8961 -7547 8963 -7513
rect 9309 -7547 9311 -7513
rect 9311 -7547 9343 -7513
rect 9381 -7547 9413 -7513
rect 9413 -7547 9415 -7513
rect 9589 -7531 9623 -7519
rect 872 -7599 906 -7591
rect 872 -7625 906 -7599
rect 872 -7667 906 -7663
rect 872 -7697 906 -7667
rect 872 -7769 906 -7735
rect 987 -7643 1021 -7641
rect 987 -7675 1021 -7643
rect 987 -7745 1021 -7713
rect 987 -7747 1021 -7745
rect 1245 -7643 1279 -7641
rect 1245 -7675 1279 -7643
rect 1245 -7745 1279 -7713
rect 1245 -7747 1279 -7745
rect 1439 -7643 1473 -7641
rect 1439 -7675 1473 -7643
rect 1439 -7745 1473 -7713
rect 1439 -7747 1473 -7745
rect 1697 -7643 1731 -7641
rect 1697 -7675 1731 -7643
rect 1697 -7745 1731 -7713
rect 1697 -7747 1731 -7745
rect 1955 -7643 1989 -7641
rect 1955 -7675 1989 -7643
rect 1955 -7745 1989 -7713
rect 1955 -7747 1989 -7745
rect 2213 -7643 2247 -7641
rect 2213 -7675 2247 -7643
rect 2213 -7745 2247 -7713
rect 2213 -7747 2247 -7745
rect 2471 -7643 2505 -7641
rect 2471 -7675 2505 -7643
rect 2471 -7745 2505 -7713
rect 2471 -7747 2505 -7745
rect 2665 -7643 2699 -7641
rect 2665 -7675 2699 -7643
rect 2665 -7745 2699 -7713
rect 2665 -7747 2699 -7745
rect 2923 -7643 2957 -7641
rect 2923 -7675 2957 -7643
rect 2923 -7745 2957 -7713
rect 2923 -7747 2957 -7745
rect 3181 -7643 3215 -7641
rect 3181 -7675 3215 -7643
rect 3181 -7745 3215 -7713
rect 3181 -7747 3215 -7745
rect 3439 -7643 3473 -7641
rect 3439 -7675 3473 -7643
rect 3439 -7745 3473 -7713
rect 3439 -7747 3473 -7745
rect 3633 -7643 3667 -7641
rect 3633 -7675 3667 -7643
rect 3633 -7745 3667 -7713
rect 3633 -7747 3667 -7745
rect 3891 -7643 3925 -7641
rect 3891 -7675 3925 -7643
rect 3891 -7745 3925 -7713
rect 3891 -7747 3925 -7745
rect 4149 -7643 4183 -7641
rect 4149 -7675 4183 -7643
rect 4149 -7745 4183 -7713
rect 4149 -7747 4183 -7745
rect 4407 -7643 4441 -7641
rect 4407 -7675 4441 -7643
rect 4407 -7745 4441 -7713
rect 4407 -7747 4441 -7745
rect 4665 -7643 4699 -7641
rect 4665 -7675 4699 -7643
rect 4665 -7745 4699 -7713
rect 4665 -7747 4699 -7745
rect 4859 -7643 4893 -7641
rect 4859 -7675 4893 -7643
rect 4859 -7745 4893 -7713
rect 4859 -7747 4893 -7745
rect 5117 -7643 5151 -7641
rect 5117 -7675 5151 -7643
rect 5117 -7745 5151 -7713
rect 5117 -7747 5151 -7745
rect 9589 -7553 9623 -7531
rect 5231 -7599 5265 -7591
rect 5231 -7625 5265 -7599
rect 5231 -7667 5265 -7663
rect 5231 -7697 5265 -7667
rect 5231 -7769 5265 -7735
rect 872 -7837 906 -7807
rect 872 -7841 906 -7837
rect 872 -7905 906 -7879
rect 872 -7913 906 -7905
rect 872 -7973 906 -7951
rect 872 -7985 906 -7973
rect 872 -8041 906 -8023
rect 872 -8057 906 -8041
rect 872 -8109 906 -8095
rect 5345 -7643 5379 -7641
rect 5345 -7675 5379 -7643
rect 5345 -7745 5379 -7713
rect 5345 -7747 5379 -7745
rect 5603 -7643 5637 -7641
rect 5603 -7675 5637 -7643
rect 5603 -7745 5637 -7713
rect 5603 -7747 5637 -7745
rect 5796 -7643 5830 -7641
rect 5796 -7675 5830 -7643
rect 5796 -7745 5830 -7713
rect 5796 -7747 5830 -7745
rect 6054 -7643 6088 -7641
rect 6054 -7675 6088 -7643
rect 6054 -7745 6088 -7713
rect 6054 -7747 6088 -7745
rect 6312 -7643 6346 -7641
rect 6312 -7675 6346 -7643
rect 6312 -7745 6346 -7713
rect 6312 -7747 6346 -7745
rect 6570 -7643 6604 -7641
rect 6570 -7675 6604 -7643
rect 6570 -7745 6604 -7713
rect 6570 -7747 6604 -7745
rect 6828 -7643 6862 -7641
rect 6828 -7675 6862 -7643
rect 6828 -7745 6862 -7713
rect 6828 -7747 6862 -7745
rect 7022 -7643 7056 -7641
rect 7022 -7675 7056 -7643
rect 7022 -7745 7056 -7713
rect 7022 -7747 7056 -7745
rect 7280 -7643 7314 -7641
rect 7280 -7675 7314 -7643
rect 7280 -7745 7314 -7713
rect 7280 -7747 7314 -7745
rect 7538 -7643 7572 -7641
rect 7538 -7675 7572 -7643
rect 7538 -7745 7572 -7713
rect 7538 -7747 7572 -7745
rect 7796 -7643 7830 -7641
rect 7796 -7675 7830 -7643
rect 7796 -7745 7830 -7713
rect 7796 -7747 7830 -7745
rect 7990 -7643 8024 -7641
rect 7990 -7675 8024 -7643
rect 7990 -7745 8024 -7713
rect 7990 -7747 8024 -7745
rect 8248 -7643 8282 -7641
rect 8248 -7675 8282 -7643
rect 8248 -7745 8282 -7713
rect 8248 -7747 8282 -7745
rect 8506 -7643 8540 -7641
rect 8506 -7675 8540 -7643
rect 8506 -7745 8540 -7713
rect 8506 -7747 8540 -7745
rect 8764 -7643 8798 -7641
rect 8764 -7675 8798 -7643
rect 8764 -7745 8798 -7713
rect 8764 -7747 8798 -7745
rect 9022 -7643 9056 -7641
rect 9022 -7675 9056 -7643
rect 9022 -7745 9056 -7713
rect 9022 -7747 9056 -7745
rect 9216 -7643 9250 -7641
rect 9216 -7675 9250 -7643
rect 9216 -7745 9250 -7713
rect 9216 -7747 9250 -7745
rect 9474 -7643 9508 -7641
rect 9474 -7675 9508 -7643
rect 9474 -7745 9508 -7713
rect 9474 -7747 9508 -7745
rect 9589 -7599 9623 -7591
rect 9589 -7625 9623 -7599
rect 9589 -7667 9623 -7663
rect 9589 -7697 9623 -7667
rect 9589 -7769 9623 -7735
rect 5231 -7837 5265 -7807
rect 5231 -7841 5265 -7837
rect 5231 -7905 5265 -7879
rect 5231 -7913 5265 -7905
rect 5231 -7973 5265 -7951
rect 5231 -7985 5265 -7973
rect 5231 -8041 5265 -8023
rect 5231 -8057 5265 -8041
rect 5231 -8109 5265 -8095
rect 9589 -7837 9623 -7807
rect 9589 -7841 9623 -7837
rect 9589 -7905 9623 -7879
rect 9589 -7913 9623 -7905
rect 9589 -7973 9623 -7951
rect 9589 -7985 9623 -7973
rect 9589 -8041 9623 -8023
rect 9589 -8057 9623 -8041
rect 9589 -8109 9623 -8095
rect 872 -8129 906 -8109
rect 5231 -8129 5265 -8109
rect 9589 -8129 9623 -8109
rect 872 -8177 906 -8167
rect 872 -8201 906 -8177
rect 872 -8245 906 -8239
rect 872 -8273 906 -8245
rect 872 -8313 906 -8311
rect 872 -8345 906 -8313
rect 872 -8415 906 -8383
rect 872 -8417 906 -8415
rect 872 -8483 906 -8455
rect 872 -8489 906 -8483
rect 872 -8551 906 -8527
rect 5231 -8177 5265 -8167
rect 5231 -8201 5265 -8177
rect 5231 -8245 5265 -8239
rect 5231 -8273 5265 -8245
rect 5231 -8313 5265 -8311
rect 5231 -8345 5265 -8313
rect 5231 -8415 5265 -8383
rect 5231 -8417 5265 -8415
rect 5231 -8483 5265 -8455
rect 5231 -8489 5265 -8483
rect 872 -8561 906 -8551
rect 872 -8619 906 -8599
rect 872 -8633 906 -8619
rect 872 -8687 906 -8671
rect 872 -8705 906 -8687
rect 987 -8587 1021 -8585
rect 987 -8619 1021 -8587
rect 987 -8689 1021 -8657
rect 987 -8691 1021 -8689
rect 1245 -8587 1279 -8585
rect 1245 -8619 1279 -8587
rect 1245 -8689 1279 -8657
rect 1245 -8691 1279 -8689
rect 1439 -8587 1473 -8585
rect 1439 -8619 1473 -8587
rect 1439 -8689 1473 -8657
rect 1439 -8691 1473 -8689
rect 1697 -8587 1731 -8585
rect 1697 -8619 1731 -8587
rect 1697 -8689 1731 -8657
rect 1697 -8691 1731 -8689
rect 1955 -8587 1989 -8585
rect 1955 -8619 1989 -8587
rect 1955 -8689 1989 -8657
rect 1955 -8691 1989 -8689
rect 2213 -8587 2247 -8585
rect 2213 -8619 2247 -8587
rect 2213 -8689 2247 -8657
rect 2213 -8691 2247 -8689
rect 2471 -8587 2505 -8585
rect 2471 -8619 2505 -8587
rect 2471 -8689 2505 -8657
rect 2471 -8691 2505 -8689
rect 2665 -8587 2699 -8585
rect 2665 -8619 2699 -8587
rect 2665 -8689 2699 -8657
rect 2665 -8691 2699 -8689
rect 2923 -8587 2957 -8585
rect 2923 -8619 2957 -8587
rect 2923 -8689 2957 -8657
rect 2923 -8691 2957 -8689
rect 3181 -8587 3215 -8585
rect 3181 -8619 3215 -8587
rect 3181 -8689 3215 -8657
rect 3181 -8691 3215 -8689
rect 3439 -8587 3473 -8585
rect 3439 -8619 3473 -8587
rect 3439 -8689 3473 -8657
rect 3439 -8691 3473 -8689
rect 3633 -8587 3667 -8585
rect 3633 -8619 3667 -8587
rect 3633 -8689 3667 -8657
rect 3633 -8691 3667 -8689
rect 3891 -8587 3925 -8585
rect 3891 -8619 3925 -8587
rect 3891 -8689 3925 -8657
rect 3891 -8691 3925 -8689
rect 4149 -8587 4183 -8585
rect 4149 -8619 4183 -8587
rect 4149 -8689 4183 -8657
rect 4149 -8691 4183 -8689
rect 4407 -8587 4441 -8585
rect 4407 -8619 4441 -8587
rect 4407 -8689 4441 -8657
rect 4407 -8691 4441 -8689
rect 4665 -8587 4699 -8585
rect 4665 -8619 4699 -8587
rect 4665 -8689 4699 -8657
rect 4665 -8691 4699 -8689
rect 4859 -8587 4893 -8585
rect 4859 -8619 4893 -8587
rect 4859 -8689 4893 -8657
rect 4859 -8691 4893 -8689
rect 5117 -8587 5151 -8585
rect 5117 -8619 5151 -8587
rect 5117 -8689 5151 -8657
rect 5117 -8691 5151 -8689
rect 5231 -8551 5265 -8527
rect 9589 -8177 9623 -8167
rect 9589 -8201 9623 -8177
rect 9589 -8245 9623 -8239
rect 9589 -8273 9623 -8245
rect 9589 -8313 9623 -8311
rect 9589 -8345 9623 -8313
rect 9589 -8415 9623 -8383
rect 9589 -8417 9623 -8415
rect 9589 -8483 9623 -8455
rect 9589 -8489 9623 -8483
rect 5231 -8561 5265 -8551
rect 5231 -8619 5265 -8599
rect 5231 -8633 5265 -8619
rect 5231 -8687 5265 -8671
rect 5231 -8705 5265 -8687
rect 872 -8777 906 -8743
rect 5345 -8587 5379 -8585
rect 5345 -8619 5379 -8587
rect 5345 -8689 5379 -8657
rect 5345 -8691 5379 -8689
rect 5603 -8587 5637 -8585
rect 5603 -8619 5637 -8587
rect 5603 -8689 5637 -8657
rect 5603 -8691 5637 -8689
rect 5796 -8587 5830 -8585
rect 5796 -8619 5830 -8587
rect 5796 -8689 5830 -8657
rect 5796 -8691 5830 -8689
rect 6054 -8587 6088 -8585
rect 6054 -8619 6088 -8587
rect 6054 -8689 6088 -8657
rect 6054 -8691 6088 -8689
rect 6312 -8587 6346 -8585
rect 6312 -8619 6346 -8587
rect 6312 -8689 6346 -8657
rect 6312 -8691 6346 -8689
rect 6570 -8587 6604 -8585
rect 6570 -8619 6604 -8587
rect 6570 -8689 6604 -8657
rect 6570 -8691 6604 -8689
rect 6828 -8587 6862 -8585
rect 6828 -8619 6862 -8587
rect 6828 -8689 6862 -8657
rect 6828 -8691 6862 -8689
rect 7022 -8587 7056 -8585
rect 7022 -8619 7056 -8587
rect 7022 -8689 7056 -8657
rect 7022 -8691 7056 -8689
rect 7280 -8587 7314 -8585
rect 7280 -8619 7314 -8587
rect 7280 -8689 7314 -8657
rect 7280 -8691 7314 -8689
rect 7538 -8587 7572 -8585
rect 7538 -8619 7572 -8587
rect 7538 -8689 7572 -8657
rect 7538 -8691 7572 -8689
rect 7796 -8587 7830 -8585
rect 7796 -8619 7830 -8587
rect 7796 -8689 7830 -8657
rect 7796 -8691 7830 -8689
rect 7990 -8587 8024 -8585
rect 7990 -8619 8024 -8587
rect 7990 -8689 8024 -8657
rect 7990 -8691 8024 -8689
rect 8248 -8587 8282 -8585
rect 8248 -8619 8282 -8587
rect 8248 -8689 8282 -8657
rect 8248 -8691 8282 -8689
rect 8506 -8587 8540 -8585
rect 8506 -8619 8540 -8587
rect 8506 -8689 8540 -8657
rect 8506 -8691 8540 -8689
rect 8764 -8587 8798 -8585
rect 8764 -8619 8798 -8587
rect 8764 -8689 8798 -8657
rect 8764 -8691 8798 -8689
rect 9022 -8587 9056 -8585
rect 9022 -8619 9056 -8587
rect 9022 -8689 9056 -8657
rect 9022 -8691 9056 -8689
rect 9216 -8587 9250 -8585
rect 9216 -8619 9250 -8587
rect 9216 -8689 9250 -8657
rect 9216 -8691 9250 -8689
rect 9474 -8587 9508 -8585
rect 9474 -8619 9508 -8587
rect 9474 -8689 9508 -8657
rect 9474 -8691 9508 -8689
rect 9589 -8551 9623 -8527
rect 9589 -8561 9623 -8551
rect 9589 -8619 9623 -8599
rect 9589 -8633 9623 -8619
rect 9589 -8687 9623 -8671
rect 9589 -8705 9623 -8687
rect 5231 -8777 5265 -8743
rect 1080 -8819 1082 -8785
rect 1082 -8819 1114 -8785
rect 1152 -8819 1184 -8785
rect 1184 -8819 1186 -8785
rect 1532 -8819 1534 -8785
rect 1534 -8819 1566 -8785
rect 1604 -8819 1636 -8785
rect 1636 -8819 1638 -8785
rect 1790 -8819 1792 -8785
rect 1792 -8819 1824 -8785
rect 1862 -8819 1894 -8785
rect 1894 -8819 1896 -8785
rect 2048 -8819 2050 -8785
rect 2050 -8819 2082 -8785
rect 2120 -8819 2152 -8785
rect 2152 -8819 2154 -8785
rect 2306 -8819 2308 -8785
rect 2308 -8819 2340 -8785
rect 2378 -8819 2410 -8785
rect 2410 -8819 2412 -8785
rect 2758 -8819 2760 -8785
rect 2760 -8819 2792 -8785
rect 2830 -8819 2862 -8785
rect 2862 -8819 2864 -8785
rect 3016 -8819 3018 -8785
rect 3018 -8819 3050 -8785
rect 3088 -8819 3120 -8785
rect 3120 -8819 3122 -8785
rect 3274 -8819 3276 -8785
rect 3276 -8819 3308 -8785
rect 3346 -8819 3378 -8785
rect 3378 -8819 3380 -8785
rect 3726 -8819 3728 -8785
rect 3728 -8819 3760 -8785
rect 3798 -8819 3830 -8785
rect 3830 -8819 3832 -8785
rect 3984 -8819 3986 -8785
rect 3986 -8819 4018 -8785
rect 4056 -8819 4088 -8785
rect 4088 -8819 4090 -8785
rect 4242 -8819 4244 -8785
rect 4244 -8819 4276 -8785
rect 4314 -8819 4346 -8785
rect 4346 -8819 4348 -8785
rect 4500 -8819 4502 -8785
rect 4502 -8819 4534 -8785
rect 4572 -8819 4604 -8785
rect 4604 -8819 4606 -8785
rect 4952 -8819 4954 -8785
rect 4954 -8819 4986 -8785
rect 5024 -8819 5056 -8785
rect 5056 -8819 5058 -8785
rect 9589 -8777 9623 -8743
rect 5438 -8819 5440 -8785
rect 5440 -8819 5472 -8785
rect 5510 -8819 5542 -8785
rect 5542 -8819 5544 -8785
rect 5889 -8819 5891 -8785
rect 5891 -8819 5923 -8785
rect 5961 -8819 5993 -8785
rect 5993 -8819 5995 -8785
rect 6147 -8819 6149 -8785
rect 6149 -8819 6181 -8785
rect 6219 -8819 6251 -8785
rect 6251 -8819 6253 -8785
rect 6405 -8819 6407 -8785
rect 6407 -8819 6439 -8785
rect 6477 -8819 6509 -8785
rect 6509 -8819 6511 -8785
rect 6663 -8819 6665 -8785
rect 6665 -8819 6697 -8785
rect 6735 -8819 6767 -8785
rect 6767 -8819 6769 -8785
rect 7115 -8819 7117 -8785
rect 7117 -8819 7149 -8785
rect 7187 -8819 7219 -8785
rect 7219 -8819 7221 -8785
rect 7373 -8819 7375 -8785
rect 7375 -8819 7407 -8785
rect 7445 -8819 7477 -8785
rect 7477 -8819 7479 -8785
rect 7631 -8819 7633 -8785
rect 7633 -8819 7665 -8785
rect 7703 -8819 7735 -8785
rect 7735 -8819 7737 -8785
rect 8083 -8819 8085 -8785
rect 8085 -8819 8117 -8785
rect 8155 -8819 8187 -8785
rect 8187 -8819 8189 -8785
rect 8341 -8819 8343 -8785
rect 8343 -8819 8375 -8785
rect 8413 -8819 8445 -8785
rect 8445 -8819 8447 -8785
rect 8599 -8819 8601 -8785
rect 8601 -8819 8633 -8785
rect 8671 -8819 8703 -8785
rect 8703 -8819 8705 -8785
rect 8857 -8819 8859 -8785
rect 8859 -8819 8891 -8785
rect 8929 -8819 8961 -8785
rect 8961 -8819 8963 -8785
rect 9309 -8819 9311 -8785
rect 9311 -8819 9343 -8785
rect 9381 -8819 9413 -8785
rect 9413 -8819 9415 -8785
rect 946 -8933 980 -8899
rect 1018 -8933 1027 -8899
rect 1027 -8933 1052 -8899
rect 1090 -8933 1095 -8899
rect 1095 -8933 1124 -8899
rect 1162 -8933 1163 -8899
rect 1163 -8933 1196 -8899
rect 1234 -8933 1265 -8899
rect 1265 -8933 1268 -8899
rect 1306 -8933 1333 -8899
rect 1333 -8933 1340 -8899
rect 1378 -8933 1401 -8899
rect 1401 -8933 1412 -8899
rect 1450 -8933 1469 -8899
rect 1469 -8933 1484 -8899
rect 1522 -8933 1537 -8899
rect 1537 -8933 1556 -8899
rect 1594 -8933 1605 -8899
rect 1605 -8933 1628 -8899
rect 1666 -8933 1673 -8899
rect 1673 -8933 1700 -8899
rect 1738 -8933 1741 -8899
rect 1741 -8933 1772 -8899
rect 1810 -8933 1843 -8899
rect 1843 -8933 1844 -8899
rect 1882 -8933 1911 -8899
rect 1911 -8933 1916 -8899
rect 1954 -8933 1979 -8899
rect 1979 -8933 1988 -8899
rect 2026 -8933 2047 -8899
rect 2047 -8933 2060 -8899
rect 2098 -8933 2115 -8899
rect 2115 -8933 2132 -8899
rect 2170 -8933 2183 -8899
rect 2183 -8933 2204 -8899
rect 2242 -8933 2251 -8899
rect 2251 -8933 2276 -8899
rect 2314 -8933 2319 -8899
rect 2319 -8933 2348 -8899
rect 2386 -8933 2387 -8899
rect 2387 -8933 2420 -8899
rect 2458 -8933 2489 -8899
rect 2489 -8933 2492 -8899
rect 2530 -8933 2557 -8899
rect 2557 -8933 2564 -8899
rect 2602 -8933 2625 -8899
rect 2625 -8933 2636 -8899
rect 2674 -8933 2693 -8899
rect 2693 -8933 2708 -8899
rect 2746 -8933 2761 -8899
rect 2761 -8933 2780 -8899
rect 2818 -8933 2829 -8899
rect 2829 -8933 2852 -8899
rect 2890 -8933 2897 -8899
rect 2897 -8933 2924 -8899
rect 2962 -8933 2965 -8899
rect 2965 -8933 2996 -8899
rect 3034 -8933 3067 -8899
rect 3067 -8933 3068 -8899
rect 3106 -8933 3135 -8899
rect 3135 -8933 3140 -8899
rect 3178 -8933 3203 -8899
rect 3203 -8933 3212 -8899
rect 3250 -8933 3271 -8899
rect 3271 -8933 3284 -8899
rect 3322 -8933 3339 -8899
rect 3339 -8933 3356 -8899
rect 3394 -8933 3407 -8899
rect 3407 -8933 3428 -8899
rect 3466 -8933 3475 -8899
rect 3475 -8933 3500 -8899
rect 3538 -8933 3543 -8899
rect 3543 -8933 3572 -8899
rect 3610 -8933 3611 -8899
rect 3611 -8933 3644 -8899
rect 3682 -8933 3713 -8899
rect 3713 -8933 3716 -8899
rect 3754 -8933 3781 -8899
rect 3781 -8933 3788 -8899
rect 3826 -8933 3849 -8899
rect 3849 -8933 3860 -8899
rect 3898 -8933 3917 -8899
rect 3917 -8933 3932 -8899
rect 3970 -8933 3985 -8899
rect 3985 -8933 4004 -8899
rect 4042 -8933 4053 -8899
rect 4053 -8933 4076 -8899
rect 4114 -8933 4121 -8899
rect 4121 -8933 4148 -8899
rect 4186 -8933 4189 -8899
rect 4189 -8933 4220 -8899
rect 4258 -8933 4291 -8899
rect 4291 -8933 4292 -8899
rect 4330 -8933 4359 -8899
rect 4359 -8933 4364 -8899
rect 4402 -8933 4427 -8899
rect 4427 -8933 4436 -8899
rect 4474 -8933 4495 -8899
rect 4495 -8933 4508 -8899
rect 4546 -8933 4563 -8899
rect 4563 -8933 4580 -8899
rect 4618 -8933 4631 -8899
rect 4631 -8933 4652 -8899
rect 4690 -8933 4699 -8899
rect 4699 -8933 4724 -8899
rect 4762 -8933 4767 -8899
rect 4767 -8933 4796 -8899
rect 4834 -8933 4835 -8899
rect 4835 -8933 4868 -8899
rect 4906 -8933 4937 -8899
rect 4937 -8933 4940 -8899
rect 4978 -8933 5005 -8899
rect 5005 -8933 5012 -8899
rect 5050 -8933 5073 -8899
rect 5073 -8933 5084 -8899
rect 5122 -8933 5156 -8899
rect 5339 -8933 5373 -8899
rect 5411 -8933 5422 -8899
rect 5422 -8933 5445 -8899
rect 5483 -8933 5490 -8899
rect 5490 -8933 5517 -8899
rect 5555 -8933 5558 -8899
rect 5558 -8933 5589 -8899
rect 5627 -8933 5660 -8899
rect 5660 -8933 5661 -8899
rect 5699 -8933 5728 -8899
rect 5728 -8933 5733 -8899
rect 5771 -8933 5796 -8899
rect 5796 -8933 5805 -8899
rect 5843 -8933 5864 -8899
rect 5864 -8933 5877 -8899
rect 5915 -8933 5932 -8899
rect 5932 -8933 5949 -8899
rect 5987 -8933 6000 -8899
rect 6000 -8933 6021 -8899
rect 6059 -8933 6068 -8899
rect 6068 -8933 6093 -8899
rect 6131 -8933 6136 -8899
rect 6136 -8933 6165 -8899
rect 6203 -8933 6204 -8899
rect 6204 -8933 6237 -8899
rect 6275 -8933 6306 -8899
rect 6306 -8933 6309 -8899
rect 6347 -8933 6374 -8899
rect 6374 -8933 6381 -8899
rect 6419 -8933 6442 -8899
rect 6442 -8933 6453 -8899
rect 6491 -8933 6510 -8899
rect 6510 -8933 6525 -8899
rect 6563 -8933 6578 -8899
rect 6578 -8933 6597 -8899
rect 6635 -8933 6646 -8899
rect 6646 -8933 6669 -8899
rect 6707 -8933 6714 -8899
rect 6714 -8933 6741 -8899
rect 6779 -8933 6782 -8899
rect 6782 -8933 6813 -8899
rect 6851 -8933 6884 -8899
rect 6884 -8933 6885 -8899
rect 6923 -8933 6952 -8899
rect 6952 -8933 6957 -8899
rect 6995 -8933 7020 -8899
rect 7020 -8933 7029 -8899
rect 7067 -8933 7088 -8899
rect 7088 -8933 7101 -8899
rect 7139 -8933 7156 -8899
rect 7156 -8933 7173 -8899
rect 7211 -8933 7224 -8899
rect 7224 -8933 7245 -8899
rect 7283 -8933 7292 -8899
rect 7292 -8933 7317 -8899
rect 7355 -8933 7360 -8899
rect 7360 -8933 7389 -8899
rect 7427 -8933 7428 -8899
rect 7428 -8933 7461 -8899
rect 7499 -8933 7530 -8899
rect 7530 -8933 7533 -8899
rect 7571 -8933 7598 -8899
rect 7598 -8933 7605 -8899
rect 7643 -8933 7666 -8899
rect 7666 -8933 7677 -8899
rect 7715 -8933 7734 -8899
rect 7734 -8933 7749 -8899
rect 7787 -8933 7802 -8899
rect 7802 -8933 7821 -8899
rect 7859 -8933 7870 -8899
rect 7870 -8933 7893 -8899
rect 7931 -8933 7938 -8899
rect 7938 -8933 7965 -8899
rect 8003 -8933 8006 -8899
rect 8006 -8933 8037 -8899
rect 8075 -8933 8108 -8899
rect 8108 -8933 8109 -8899
rect 8147 -8933 8176 -8899
rect 8176 -8933 8181 -8899
rect 8219 -8933 8244 -8899
rect 8244 -8933 8253 -8899
rect 8291 -8933 8312 -8899
rect 8312 -8933 8325 -8899
rect 8363 -8933 8380 -8899
rect 8380 -8933 8397 -8899
rect 8435 -8933 8448 -8899
rect 8448 -8933 8469 -8899
rect 8507 -8933 8516 -8899
rect 8516 -8933 8541 -8899
rect 8579 -8933 8584 -8899
rect 8584 -8933 8613 -8899
rect 8651 -8933 8652 -8899
rect 8652 -8933 8685 -8899
rect 8723 -8933 8754 -8899
rect 8754 -8933 8757 -8899
rect 8795 -8933 8822 -8899
rect 8822 -8933 8829 -8899
rect 8867 -8933 8890 -8899
rect 8890 -8933 8901 -8899
rect 8939 -8933 8958 -8899
rect 8958 -8933 8973 -8899
rect 9011 -8933 9026 -8899
rect 9026 -8933 9045 -8899
rect 9083 -8933 9094 -8899
rect 9094 -8933 9117 -8899
rect 9155 -8933 9162 -8899
rect 9162 -8933 9189 -8899
rect 9227 -8933 9230 -8899
rect 9230 -8933 9261 -8899
rect 9299 -8933 9332 -8899
rect 9332 -8933 9333 -8899
rect 9371 -8933 9400 -8899
rect 9400 -8933 9405 -8899
rect 9443 -8933 9468 -8899
rect 9468 -8933 9477 -8899
rect 9515 -8933 9549 -8899
<< metal1 >>
rect 847 756 9648 781
rect 847 722 946 756
rect 980 722 1018 756
rect 1052 722 1090 756
rect 1124 722 1162 756
rect 1196 722 1234 756
rect 1268 722 1306 756
rect 1340 722 1378 756
rect 1412 722 1450 756
rect 1484 722 1522 756
rect 1556 722 1594 756
rect 1628 722 1666 756
rect 1700 722 1738 756
rect 1772 722 1810 756
rect 1844 722 1882 756
rect 1916 722 1954 756
rect 1988 722 2026 756
rect 2060 722 2098 756
rect 2132 722 2170 756
rect 2204 722 2242 756
rect 2276 722 2314 756
rect 2348 722 2386 756
rect 2420 722 2458 756
rect 2492 722 2530 756
rect 2564 722 2602 756
rect 2636 722 2674 756
rect 2708 722 2746 756
rect 2780 722 2818 756
rect 2852 722 2890 756
rect 2924 722 2962 756
rect 2996 722 3034 756
rect 3068 722 3106 756
rect 3140 722 3178 756
rect 3212 722 3250 756
rect 3284 722 3322 756
rect 3356 722 3394 756
rect 3428 722 3466 756
rect 3500 722 3538 756
rect 3572 722 3610 756
rect 3644 722 3682 756
rect 3716 722 3754 756
rect 3788 722 3826 756
rect 3860 722 3898 756
rect 3932 722 3970 756
rect 4004 722 4042 756
rect 4076 722 4114 756
rect 4148 722 4186 756
rect 4220 722 4258 756
rect 4292 722 4330 756
rect 4364 722 4402 756
rect 4436 722 4474 756
rect 4508 722 4546 756
rect 4580 722 4618 756
rect 4652 722 4690 756
rect 4724 722 4762 756
rect 4796 722 4834 756
rect 4868 722 4906 756
rect 4940 722 4978 756
rect 5012 722 5050 756
rect 5084 722 5122 756
rect 5156 722 5339 756
rect 5373 722 5411 756
rect 5445 722 5483 756
rect 5517 722 5555 756
rect 5589 722 5627 756
rect 5661 722 5699 756
rect 5733 722 5771 756
rect 5805 722 5843 756
rect 5877 722 5915 756
rect 5949 722 5987 756
rect 6021 722 6059 756
rect 6093 722 6131 756
rect 6165 722 6203 756
rect 6237 722 6275 756
rect 6309 722 6347 756
rect 6381 722 6419 756
rect 6453 722 6491 756
rect 6525 722 6563 756
rect 6597 722 6635 756
rect 6669 722 6707 756
rect 6741 722 6779 756
rect 6813 722 6851 756
rect 6885 722 6923 756
rect 6957 722 6995 756
rect 7029 722 7067 756
rect 7101 722 7139 756
rect 7173 722 7211 756
rect 7245 722 7283 756
rect 7317 722 7355 756
rect 7389 722 7427 756
rect 7461 722 7499 756
rect 7533 722 7571 756
rect 7605 722 7643 756
rect 7677 722 7715 756
rect 7749 722 7787 756
rect 7821 722 7859 756
rect 7893 722 7931 756
rect 7965 722 8003 756
rect 8037 722 8075 756
rect 8109 722 8147 756
rect 8181 722 8219 756
rect 8253 722 8291 756
rect 8325 722 8363 756
rect 8397 722 8435 756
rect 8469 722 8507 756
rect 8541 722 8579 756
rect 8613 722 8651 756
rect 8685 722 8723 756
rect 8757 722 8795 756
rect 8829 722 8867 756
rect 8901 722 8939 756
rect 8973 722 9011 756
rect 9045 722 9083 756
rect 9117 722 9155 756
rect 9189 722 9227 756
rect 9261 722 9299 756
rect 9333 722 9371 756
rect 9405 722 9443 756
rect 9477 722 9515 756
rect 9549 722 9648 756
rect 847 642 9648 722
rect 847 608 1080 642
rect 1114 608 1152 642
rect 1186 608 1532 642
rect 1566 608 1604 642
rect 1638 608 1790 642
rect 1824 608 1862 642
rect 1896 608 2048 642
rect 2082 608 2120 642
rect 2154 608 2306 642
rect 2340 608 2378 642
rect 2412 608 2758 642
rect 2792 608 2830 642
rect 2864 608 3016 642
rect 3050 608 3088 642
rect 3122 608 3274 642
rect 3308 608 3346 642
rect 3380 608 3726 642
rect 3760 608 3798 642
rect 3832 608 3984 642
rect 4018 608 4056 642
rect 4090 608 4242 642
rect 4276 608 4314 642
rect 4348 608 4500 642
rect 4534 608 4572 642
rect 4606 608 4952 642
rect 4986 608 5024 642
rect 5058 608 5438 642
rect 5472 608 5510 642
rect 5544 608 5889 642
rect 5923 608 5961 642
rect 5995 608 6147 642
rect 6181 608 6219 642
rect 6253 608 6405 642
rect 6439 608 6477 642
rect 6511 608 6663 642
rect 6697 608 6735 642
rect 6769 608 7115 642
rect 7149 608 7187 642
rect 7221 608 7373 642
rect 7407 608 7445 642
rect 7479 608 7631 642
rect 7665 608 7703 642
rect 7737 608 8083 642
rect 8117 608 8155 642
rect 8189 608 8341 642
rect 8375 608 8413 642
rect 8447 608 8599 642
rect 8633 608 8671 642
rect 8705 608 8857 642
rect 8891 608 8929 642
rect 8963 608 9309 642
rect 9343 608 9381 642
rect 9415 608 9648 642
rect 847 602 9648 608
rect 849 599 1285 602
rect 849 565 872 599
rect 906 565 1285 599
rect 849 527 1285 565
rect 849 493 872 527
rect 906 514 1285 527
rect 906 493 987 514
rect 849 480 987 493
rect 1021 480 1245 514
rect 1279 480 1285 514
rect 849 455 1285 480
rect 849 421 872 455
rect 906 442 1285 455
rect 906 421 987 442
rect 849 408 987 421
rect 1021 408 1245 442
rect 1279 408 1285 442
rect 849 383 1285 408
rect 849 349 872 383
rect 906 349 1285 383
rect 1433 514 1479 602
rect 1433 480 1439 514
rect 1473 480 1479 514
rect 1433 442 1479 480
rect 1433 408 1439 442
rect 1473 408 1479 442
rect 1433 361 1479 408
rect 1691 514 1737 602
rect 1691 480 1697 514
rect 1731 480 1737 514
rect 1691 442 1737 480
rect 1691 408 1697 442
rect 1731 408 1737 442
rect 1691 361 1737 408
rect 1949 514 1995 602
rect 1949 480 1955 514
rect 1989 480 1995 514
rect 1949 442 1995 480
rect 1949 408 1955 442
rect 1989 408 1995 442
rect 1949 361 1995 408
rect 2207 514 2253 602
rect 2207 480 2213 514
rect 2247 480 2253 514
rect 2207 442 2253 480
rect 2207 408 2213 442
rect 2247 408 2253 442
rect 2207 361 2253 408
rect 2465 514 2511 602
rect 2465 480 2471 514
rect 2505 480 2511 514
rect 2465 442 2511 480
rect 2465 408 2471 442
rect 2505 408 2511 442
rect 2465 361 2511 408
rect 2659 514 2705 602
rect 2659 480 2665 514
rect 2699 480 2705 514
rect 2659 442 2705 480
rect 2659 408 2665 442
rect 2699 408 2705 442
rect 2659 361 2705 408
rect 2917 514 2963 602
rect 2917 480 2923 514
rect 2957 480 2963 514
rect 2917 442 2963 480
rect 2917 408 2923 442
rect 2957 408 2963 442
rect 2917 361 2963 408
rect 3175 514 3221 602
rect 3175 480 3181 514
rect 3215 480 3221 514
rect 3175 442 3221 480
rect 3175 408 3181 442
rect 3215 408 3221 442
rect 3175 361 3221 408
rect 3433 514 3479 602
rect 3433 480 3439 514
rect 3473 480 3479 514
rect 3433 442 3479 480
rect 3433 408 3439 442
rect 3473 408 3479 442
rect 3433 361 3479 408
rect 3627 514 3673 602
rect 3627 480 3633 514
rect 3667 480 3673 514
rect 3627 442 3673 480
rect 3627 408 3633 442
rect 3667 408 3673 442
rect 3627 361 3673 408
rect 3885 514 3931 602
rect 3885 480 3891 514
rect 3925 480 3931 514
rect 3885 442 3931 480
rect 3885 408 3891 442
rect 3925 408 3931 442
rect 3885 361 3931 408
rect 4143 514 4189 602
rect 4143 480 4149 514
rect 4183 480 4189 514
rect 4143 442 4189 480
rect 4143 408 4149 442
rect 4183 408 4189 442
rect 4143 361 4189 408
rect 4401 514 4447 602
rect 4401 480 4407 514
rect 4441 480 4447 514
rect 4401 442 4447 480
rect 4401 408 4407 442
rect 4441 408 4447 442
rect 4401 361 4447 408
rect 4659 514 4705 602
rect 4659 480 4665 514
rect 4699 480 4705 514
rect 4659 442 4705 480
rect 4659 408 4665 442
rect 4699 408 4705 442
rect 4659 361 4705 408
rect 4853 599 5643 602
rect 4853 565 5231 599
rect 5265 565 5643 599
rect 4853 527 5643 565
rect 4853 514 5231 527
rect 4853 480 4859 514
rect 4893 480 5117 514
rect 5151 493 5231 514
rect 5265 514 5643 527
rect 5265 493 5345 514
rect 5151 480 5345 493
rect 5379 480 5603 514
rect 5637 480 5643 514
rect 4853 455 5643 480
rect 4853 442 5231 455
rect 4853 408 4859 442
rect 4893 408 5117 442
rect 5151 421 5231 442
rect 5265 442 5643 455
rect 5265 421 5345 442
rect 5151 408 5345 421
rect 5379 408 5603 442
rect 5637 408 5643 442
rect 4853 383 5643 408
rect 849 311 1285 349
rect 849 277 872 311
rect 906 277 1285 311
rect 4853 349 5231 383
rect 5265 349 5643 383
rect 5790 514 5836 602
rect 5790 480 5796 514
rect 5830 480 5836 514
rect 5790 442 5836 480
rect 5790 408 5796 442
rect 5830 408 5836 442
rect 5790 361 5836 408
rect 6048 514 6094 602
rect 6048 480 6054 514
rect 6088 480 6094 514
rect 6048 442 6094 480
rect 6048 408 6054 442
rect 6088 408 6094 442
rect 6048 361 6094 408
rect 6306 514 6352 602
rect 6306 480 6312 514
rect 6346 480 6352 514
rect 6306 442 6352 480
rect 6306 408 6312 442
rect 6346 408 6352 442
rect 6306 361 6352 408
rect 6564 514 6610 602
rect 6564 480 6570 514
rect 6604 480 6610 514
rect 6564 442 6610 480
rect 6564 408 6570 442
rect 6604 408 6610 442
rect 6564 361 6610 408
rect 6822 514 6868 602
rect 6822 480 6828 514
rect 6862 480 6868 514
rect 6822 442 6868 480
rect 6822 408 6828 442
rect 6862 408 6868 442
rect 6822 361 6868 408
rect 7016 514 7062 602
rect 7016 480 7022 514
rect 7056 480 7062 514
rect 7016 442 7062 480
rect 7016 408 7022 442
rect 7056 408 7062 442
rect 7016 361 7062 408
rect 7274 514 7320 602
rect 7274 480 7280 514
rect 7314 480 7320 514
rect 7274 442 7320 480
rect 7274 408 7280 442
rect 7314 408 7320 442
rect 7274 361 7320 408
rect 7532 514 7578 602
rect 7532 480 7538 514
rect 7572 480 7578 514
rect 7532 442 7578 480
rect 7532 408 7538 442
rect 7572 408 7578 442
rect 7532 361 7578 408
rect 7790 514 7836 602
rect 7790 480 7796 514
rect 7830 480 7836 514
rect 7790 442 7836 480
rect 7790 408 7796 442
rect 7830 408 7836 442
rect 7790 361 7836 408
rect 7984 514 8030 602
rect 7984 480 7990 514
rect 8024 480 8030 514
rect 7984 442 8030 480
rect 7984 408 7990 442
rect 8024 408 8030 442
rect 7984 361 8030 408
rect 8242 514 8288 602
rect 8242 480 8248 514
rect 8282 480 8288 514
rect 8242 442 8288 480
rect 8242 408 8248 442
rect 8282 408 8288 442
rect 8242 361 8288 408
rect 8500 514 8546 602
rect 8500 480 8506 514
rect 8540 480 8546 514
rect 8500 442 8546 480
rect 8500 408 8506 442
rect 8540 408 8546 442
rect 8500 361 8546 408
rect 8758 514 8804 602
rect 8758 480 8764 514
rect 8798 480 8804 514
rect 8758 442 8804 480
rect 8758 408 8764 442
rect 8798 408 8804 442
rect 8758 361 8804 408
rect 9016 514 9062 602
rect 9016 480 9022 514
rect 9056 480 9062 514
rect 9016 442 9062 480
rect 9016 408 9022 442
rect 9056 408 9062 442
rect 9016 361 9062 408
rect 9210 599 9646 602
rect 9210 565 9589 599
rect 9623 565 9646 599
rect 9210 527 9646 565
rect 9210 514 9589 527
rect 9210 480 9216 514
rect 9250 480 9474 514
rect 9508 493 9589 514
rect 9623 493 9646 527
rect 9508 480 9646 493
rect 9210 455 9646 480
rect 9210 442 9589 455
rect 9210 408 9216 442
rect 9250 408 9474 442
rect 9508 421 9589 442
rect 9623 421 9646 455
rect 9508 408 9646 421
rect 9210 383 9646 408
rect 4853 311 5643 349
rect 849 239 1285 277
rect 849 205 872 239
rect 906 205 1285 239
rect 2843 281 3039 289
rect 2843 229 2850 281
rect 2902 229 2914 281
rect 2966 229 2978 281
rect 3030 229 3039 281
rect 2843 219 3039 229
rect 3361 281 3557 289
rect 3361 229 3368 281
rect 3420 229 3432 281
rect 3484 229 3496 281
rect 3548 229 3557 281
rect 3361 219 3557 229
rect 4853 277 5231 311
rect 5265 277 5643 311
rect 9210 349 9589 383
rect 9623 349 9646 383
rect 9210 311 9646 349
rect 4853 239 5643 277
rect 849 167 1285 205
rect 849 133 872 167
rect 906 133 1285 167
rect 849 95 1285 133
rect 849 61 872 95
rect 906 61 1285 95
rect 849 23 1285 61
rect 1355 112 1551 120
rect 1355 60 1364 112
rect 1416 60 1428 112
rect 1480 60 1492 112
rect 1544 60 1551 112
rect 1355 50 1551 60
rect 1873 112 2069 120
rect 1873 60 1882 112
rect 1934 60 1946 112
rect 1998 60 2010 112
rect 2062 60 2069 112
rect 1873 50 2069 60
rect 2389 112 2585 120
rect 2389 60 2398 112
rect 2450 60 2462 112
rect 2514 60 2526 112
rect 2578 60 2585 112
rect 2389 50 2585 60
rect 849 -11 872 23
rect 906 -11 1285 23
rect 849 -49 1285 -11
rect 849 -83 872 -49
rect 906 -83 1285 -49
rect 849 -121 1285 -83
rect 849 -155 872 -121
rect 906 -155 1285 -121
rect 849 -193 1285 -155
rect 849 -227 872 -193
rect 906 -227 1285 -193
rect 849 -265 1285 -227
rect 849 -299 872 -265
rect 906 -299 1285 -265
rect 849 -337 1285 -299
rect 849 -371 872 -337
rect 906 -371 1285 -337
rect 849 -409 1285 -371
rect 849 -443 872 -409
rect 906 -430 1285 -409
rect 906 -443 987 -430
rect 849 -464 987 -443
rect 1021 -464 1245 -430
rect 1279 -464 1285 -430
rect 849 -481 1285 -464
rect 849 -515 872 -481
rect 906 -502 1285 -481
rect 906 -515 987 -502
rect 849 -536 987 -515
rect 1021 -536 1245 -502
rect 1279 -536 1285 -502
rect 849 -553 1285 -536
rect 849 -587 872 -553
rect 906 -587 1285 -553
rect 1433 -430 1479 50
rect 1615 -219 1811 -211
rect 1615 -271 1624 -219
rect 1676 -271 1688 -219
rect 1740 -271 1752 -219
rect 1804 -271 1811 -219
rect 1615 -281 1811 -271
rect 1433 -464 1439 -430
rect 1473 -464 1479 -430
rect 1433 -502 1479 -464
rect 1433 -536 1439 -502
rect 1473 -536 1479 -502
rect 1433 -583 1479 -536
rect 1691 -430 1737 -281
rect 1691 -464 1697 -430
rect 1731 -464 1737 -430
rect 1691 -502 1737 -464
rect 1691 -536 1697 -502
rect 1731 -536 1737 -502
rect 1691 -583 1737 -536
rect 1949 -430 1995 50
rect 2132 -219 2328 -211
rect 2132 -271 2141 -219
rect 2193 -271 2205 -219
rect 2257 -271 2269 -219
rect 2321 -271 2328 -219
rect 2132 -281 2328 -271
rect 1949 -464 1955 -430
rect 1989 -464 1995 -430
rect 1949 -502 1995 -464
rect 1949 -536 1955 -502
rect 1989 -536 1995 -502
rect 1949 -583 1995 -536
rect 2207 -430 2253 -281
rect 2207 -464 2213 -430
rect 2247 -464 2253 -430
rect 2207 -502 2253 -464
rect 2207 -536 2213 -502
rect 2247 -536 2253 -502
rect 2207 -583 2253 -536
rect 2465 -430 2511 50
rect 2586 -51 2782 -43
rect 2586 -103 2593 -51
rect 2645 -103 2657 -51
rect 2709 -103 2721 -51
rect 2773 -103 2782 -51
rect 2586 -113 2782 -103
rect 2465 -464 2471 -430
rect 2505 -464 2511 -430
rect 2465 -502 2511 -464
rect 2465 -536 2471 -502
rect 2505 -536 2511 -502
rect 2465 -583 2511 -536
rect 2659 -430 2705 -113
rect 2659 -464 2665 -430
rect 2699 -464 2705 -430
rect 2659 -502 2705 -464
rect 2659 -536 2665 -502
rect 2699 -536 2705 -502
rect 2659 -583 2705 -536
rect 2917 -430 2963 219
rect 3103 -51 3299 -43
rect 3103 -103 3110 -51
rect 3162 -103 3174 -51
rect 3226 -103 3238 -51
rect 3290 -103 3299 -51
rect 3103 -113 3299 -103
rect 2917 -464 2923 -430
rect 2957 -464 2963 -430
rect 2917 -502 2963 -464
rect 2917 -536 2923 -502
rect 2957 -536 2963 -502
rect 2917 -583 2963 -536
rect 3175 -430 3221 -113
rect 3175 -464 3181 -430
rect 3215 -464 3221 -430
rect 3175 -502 3221 -464
rect 3175 -536 3181 -502
rect 3215 -536 3221 -502
rect 3175 -583 3221 -536
rect 3433 -430 3479 219
rect 4853 205 5231 239
rect 5265 205 5643 239
rect 6939 281 7135 289
rect 6939 229 6948 281
rect 7000 229 7012 281
rect 7064 229 7076 281
rect 7128 229 7135 281
rect 6939 219 7135 229
rect 7456 281 7652 289
rect 7456 229 7465 281
rect 7517 229 7529 281
rect 7581 229 7593 281
rect 7645 229 7652 281
rect 7456 219 7652 229
rect 9210 277 9589 311
rect 9623 277 9646 311
rect 9210 239 9646 277
rect 4853 167 5643 205
rect 4853 133 5231 167
rect 5265 133 5643 167
rect 3550 112 3746 120
rect 3550 60 3559 112
rect 3611 60 3623 112
rect 3675 60 3687 112
rect 3739 60 3746 112
rect 3550 50 3746 60
rect 4067 112 4263 120
rect 4067 60 4076 112
rect 4128 60 4140 112
rect 4192 60 4204 112
rect 4256 60 4263 112
rect 4067 50 4263 60
rect 4582 112 4778 120
rect 4582 60 4591 112
rect 4643 60 4655 112
rect 4707 60 4719 112
rect 4771 60 4778 112
rect 4582 50 4778 60
rect 4853 95 5643 133
rect 4853 61 5231 95
rect 5265 61 5643 95
rect 3433 -464 3439 -430
rect 3473 -464 3479 -430
rect 3433 -502 3479 -464
rect 3433 -536 3439 -502
rect 3473 -536 3479 -502
rect 3433 -583 3479 -536
rect 3627 -430 3673 50
rect 3809 -219 4005 -211
rect 3809 -271 3818 -219
rect 3870 -271 3882 -219
rect 3934 -271 3946 -219
rect 3998 -271 4005 -219
rect 3809 -281 4005 -271
rect 3627 -464 3633 -430
rect 3667 -464 3673 -430
rect 3627 -502 3673 -464
rect 3627 -536 3633 -502
rect 3667 -536 3673 -502
rect 3627 -583 3673 -536
rect 3885 -430 3931 -281
rect 3885 -464 3891 -430
rect 3925 -464 3931 -430
rect 3885 -502 3931 -464
rect 3885 -536 3891 -502
rect 3925 -536 3931 -502
rect 3885 -583 3931 -536
rect 4143 -430 4189 50
rect 4326 -219 4522 -211
rect 4326 -271 4335 -219
rect 4387 -271 4399 -219
rect 4451 -271 4463 -219
rect 4515 -271 4522 -219
rect 4326 -281 4522 -271
rect 4143 -464 4149 -430
rect 4183 -464 4189 -430
rect 4143 -502 4189 -464
rect 4143 -536 4149 -502
rect 4183 -536 4189 -502
rect 4143 -583 4189 -536
rect 4401 -430 4447 -281
rect 4401 -464 4407 -430
rect 4441 -464 4447 -430
rect 4401 -502 4447 -464
rect 4401 -536 4407 -502
rect 4441 -536 4447 -502
rect 4401 -583 4447 -536
rect 4659 -430 4705 50
rect 4659 -464 4665 -430
rect 4699 -464 4705 -430
rect 4659 -502 4705 -464
rect 4659 -536 4665 -502
rect 4699 -536 4705 -502
rect 4659 -583 4705 -536
rect 4853 23 5643 61
rect 5717 112 5913 120
rect 5717 60 5724 112
rect 5776 60 5788 112
rect 5840 60 5852 112
rect 5904 60 5913 112
rect 5717 50 5913 60
rect 6232 112 6428 120
rect 6232 60 6239 112
rect 6291 60 6303 112
rect 6355 60 6367 112
rect 6419 60 6428 112
rect 6232 50 6428 60
rect 6749 112 6945 120
rect 6749 60 6756 112
rect 6808 60 6820 112
rect 6872 60 6884 112
rect 6936 60 6945 112
rect 6749 50 6945 60
rect 4853 -11 5231 23
rect 5265 -11 5643 23
rect 4853 -49 5643 -11
rect 4853 -83 5231 -49
rect 5265 -83 5643 -49
rect 4853 -121 5643 -83
rect 4853 -155 5231 -121
rect 5265 -155 5643 -121
rect 4853 -193 5643 -155
rect 4853 -227 5231 -193
rect 5265 -227 5643 -193
rect 4853 -265 5643 -227
rect 4853 -299 5231 -265
rect 5265 -299 5643 -265
rect 4853 -337 5643 -299
rect 4853 -371 5231 -337
rect 5265 -371 5643 -337
rect 4853 -409 5643 -371
rect 4853 -430 5231 -409
rect 4853 -464 4859 -430
rect 4893 -464 5117 -430
rect 5151 -443 5231 -430
rect 5265 -430 5643 -409
rect 5265 -443 5345 -430
rect 5151 -464 5345 -443
rect 5379 -464 5603 -430
rect 5637 -464 5643 -430
rect 4853 -481 5643 -464
rect 4853 -502 5231 -481
rect 4853 -536 4859 -502
rect 4893 -536 5117 -502
rect 5151 -515 5231 -502
rect 5265 -502 5643 -481
rect 5265 -515 5345 -502
rect 5151 -536 5345 -515
rect 5379 -536 5603 -502
rect 5637 -536 5643 -502
rect 4853 -553 5643 -536
rect 849 -625 1285 -587
rect 4853 -587 5231 -553
rect 5265 -587 5643 -553
rect 5790 -430 5836 50
rect 5973 -219 6169 -211
rect 5973 -271 5980 -219
rect 6032 -271 6044 -219
rect 6096 -271 6108 -219
rect 6160 -271 6169 -219
rect 5973 -281 6169 -271
rect 5790 -464 5796 -430
rect 5830 -464 5836 -430
rect 5790 -502 5836 -464
rect 5790 -536 5796 -502
rect 5830 -536 5836 -502
rect 5790 -583 5836 -536
rect 6048 -430 6094 -281
rect 6048 -464 6054 -430
rect 6088 -464 6094 -430
rect 6048 -502 6094 -464
rect 6048 -536 6054 -502
rect 6088 -536 6094 -502
rect 6048 -583 6094 -536
rect 6306 -430 6352 50
rect 6490 -219 6686 -211
rect 6490 -271 6497 -219
rect 6549 -271 6561 -219
rect 6613 -271 6625 -219
rect 6677 -271 6686 -219
rect 6490 -281 6686 -271
rect 6306 -464 6312 -430
rect 6346 -464 6352 -430
rect 6306 -502 6352 -464
rect 6306 -536 6312 -502
rect 6346 -536 6352 -502
rect 6306 -583 6352 -536
rect 6564 -430 6610 -281
rect 6564 -464 6570 -430
rect 6604 -464 6610 -430
rect 6564 -502 6610 -464
rect 6564 -536 6570 -502
rect 6604 -536 6610 -502
rect 6564 -583 6610 -536
rect 6822 -430 6868 50
rect 6822 -464 6828 -430
rect 6862 -464 6868 -430
rect 6822 -502 6868 -464
rect 6822 -536 6828 -502
rect 6862 -536 6868 -502
rect 6822 -583 6868 -536
rect 7016 -430 7062 219
rect 7196 -51 7392 -43
rect 7196 -103 7205 -51
rect 7257 -103 7269 -51
rect 7321 -103 7333 -51
rect 7385 -103 7392 -51
rect 7196 -113 7392 -103
rect 7016 -464 7022 -430
rect 7056 -464 7062 -430
rect 7016 -502 7062 -464
rect 7016 -536 7022 -502
rect 7056 -536 7062 -502
rect 7016 -583 7062 -536
rect 7274 -430 7320 -113
rect 7274 -464 7280 -430
rect 7314 -464 7320 -430
rect 7274 -502 7320 -464
rect 7274 -536 7280 -502
rect 7314 -536 7320 -502
rect 7274 -583 7320 -536
rect 7532 -430 7578 219
rect 9210 205 9589 239
rect 9623 205 9646 239
rect 9210 167 9646 205
rect 9210 133 9589 167
rect 9623 133 9646 167
rect 7910 112 8106 120
rect 7910 60 7917 112
rect 7969 60 7981 112
rect 8033 60 8045 112
rect 8097 60 8106 112
rect 7910 50 8106 60
rect 8427 112 8623 120
rect 8427 60 8434 112
rect 8486 60 8498 112
rect 8550 60 8562 112
rect 8614 60 8623 112
rect 8427 50 8623 60
rect 8944 112 9140 120
rect 8944 60 8951 112
rect 9003 60 9015 112
rect 9067 60 9079 112
rect 9131 60 9140 112
rect 8944 50 9140 60
rect 9210 95 9646 133
rect 9210 61 9589 95
rect 9623 61 9646 95
rect 7713 -51 7909 -43
rect 7713 -103 7722 -51
rect 7774 -103 7786 -51
rect 7838 -103 7850 -51
rect 7902 -103 7909 -51
rect 7713 -113 7909 -103
rect 7532 -464 7538 -430
rect 7572 -464 7578 -430
rect 7532 -502 7578 -464
rect 7532 -536 7538 -502
rect 7572 -536 7578 -502
rect 7532 -583 7578 -536
rect 7790 -430 7836 -113
rect 7790 -464 7796 -430
rect 7830 -464 7836 -430
rect 7790 -502 7836 -464
rect 7790 -536 7796 -502
rect 7830 -536 7836 -502
rect 7790 -583 7836 -536
rect 7984 -430 8030 50
rect 8167 -219 8363 -211
rect 8167 -271 8174 -219
rect 8226 -271 8238 -219
rect 8290 -271 8302 -219
rect 8354 -271 8363 -219
rect 8167 -281 8363 -271
rect 7984 -464 7990 -430
rect 8024 -464 8030 -430
rect 7984 -502 8030 -464
rect 7984 -536 7990 -502
rect 8024 -536 8030 -502
rect 7984 -583 8030 -536
rect 8242 -430 8288 -281
rect 8242 -464 8248 -430
rect 8282 -464 8288 -430
rect 8242 -502 8288 -464
rect 8242 -536 8248 -502
rect 8282 -536 8288 -502
rect 8242 -583 8288 -536
rect 8500 -430 8546 50
rect 8685 -219 8881 -211
rect 8685 -271 8692 -219
rect 8744 -271 8756 -219
rect 8808 -271 8820 -219
rect 8872 -271 8881 -219
rect 8685 -281 8881 -271
rect 8500 -464 8506 -430
rect 8540 -464 8546 -430
rect 8500 -502 8546 -464
rect 8500 -536 8506 -502
rect 8540 -536 8546 -502
rect 8500 -583 8546 -536
rect 8758 -430 8804 -281
rect 8758 -464 8764 -430
rect 8798 -464 8804 -430
rect 8758 -502 8804 -464
rect 8758 -536 8764 -502
rect 8798 -536 8804 -502
rect 8758 -583 8804 -536
rect 9016 -430 9062 50
rect 9016 -464 9022 -430
rect 9056 -464 9062 -430
rect 9016 -502 9062 -464
rect 9016 -536 9022 -502
rect 9056 -536 9062 -502
rect 9016 -583 9062 -536
rect 9210 23 9646 61
rect 9210 -11 9589 23
rect 9623 -11 9646 23
rect 9210 -49 9646 -11
rect 9210 -83 9589 -49
rect 9623 -83 9646 -49
rect 9210 -121 9646 -83
rect 9210 -155 9589 -121
rect 9623 -155 9646 -121
rect 9210 -193 9646 -155
rect 9210 -227 9589 -193
rect 9623 -227 9646 -193
rect 9210 -265 9646 -227
rect 9210 -299 9589 -265
rect 9623 -299 9646 -265
rect 9210 -337 9646 -299
rect 9210 -371 9589 -337
rect 9623 -371 9646 -337
rect 9210 -409 9646 -371
rect 9210 -430 9589 -409
rect 9210 -464 9216 -430
rect 9250 -464 9474 -430
rect 9508 -443 9589 -430
rect 9623 -443 9646 -409
rect 9508 -464 9646 -443
rect 9210 -481 9646 -464
rect 9210 -502 9589 -481
rect 9210 -536 9216 -502
rect 9250 -536 9474 -502
rect 9508 -515 9589 -502
rect 9623 -515 9646 -481
rect 9508 -536 9646 -515
rect 9210 -553 9646 -536
rect 849 -659 872 -625
rect 906 -630 1285 -625
rect 906 -659 1080 -630
rect 849 -664 1080 -659
rect 1114 -664 1152 -630
rect 1186 -664 1285 -630
rect 849 -697 1285 -664
rect 849 -731 872 -697
rect 906 -731 1285 -697
rect 1489 -630 2593 -624
rect 1489 -664 1532 -630
rect 1566 -643 1604 -630
rect 1638 -643 1790 -630
rect 1824 -643 1862 -630
rect 1896 -643 2048 -630
rect 2082 -643 2120 -630
rect 2154 -643 2306 -630
rect 2340 -643 2378 -630
rect 1489 -695 1539 -664
rect 1591 -695 1603 -643
rect 1655 -695 1667 -643
rect 1719 -695 1735 -643
rect 1787 -664 1790 -643
rect 1851 -664 1862 -643
rect 1787 -695 1799 -664
rect 1851 -695 1863 -664
rect 1915 -695 2025 -643
rect 2082 -664 2089 -643
rect 2077 -695 2089 -664
rect 2141 -695 2153 -664
rect 2205 -695 2221 -643
rect 2273 -695 2285 -643
rect 2340 -664 2349 -643
rect 2412 -664 2593 -630
rect 2337 -695 2349 -664
rect 2401 -695 2593 -664
rect 1489 -713 2593 -695
rect 849 -769 1285 -731
rect 849 -803 872 -769
rect 906 -803 1285 -769
rect 849 -841 1285 -803
rect 849 -875 872 -841
rect 906 -875 1285 -841
rect 849 -913 1285 -875
rect 849 -947 872 -913
rect 906 -947 1285 -913
rect 849 -985 1285 -947
rect 849 -1019 872 -985
rect 906 -993 1285 -985
rect 906 -1019 1080 -993
rect 849 -1027 1080 -1019
rect 1114 -1027 1152 -993
rect 1186 -1027 1285 -993
rect 849 -1057 1285 -1027
rect 1489 -781 2455 -763
rect 1489 -833 1539 -781
rect 1591 -833 1603 -781
rect 1655 -833 1667 -781
rect 1719 -833 1735 -781
rect 1787 -833 1799 -781
rect 1851 -833 1863 -781
rect 1915 -833 2025 -781
rect 2077 -833 2089 -781
rect 2141 -833 2153 -781
rect 2205 -833 2221 -781
rect 2273 -833 2285 -781
rect 2337 -833 2349 -781
rect 2401 -833 2455 -781
rect 1489 -959 2455 -833
rect 1489 -993 1539 -959
rect 1489 -1027 1532 -993
rect 1591 -1011 1603 -959
rect 1655 -1011 1667 -959
rect 1719 -1011 1735 -959
rect 1787 -993 1799 -959
rect 1851 -993 1863 -959
rect 1787 -1011 1790 -993
rect 1851 -1011 1862 -993
rect 1915 -1011 2025 -959
rect 2077 -993 2089 -959
rect 2141 -993 2153 -959
rect 2082 -1011 2089 -993
rect 2205 -1011 2221 -959
rect 2273 -1011 2285 -959
rect 2337 -993 2349 -959
rect 2401 -993 2455 -959
rect 2340 -1011 2349 -993
rect 1566 -1027 1604 -1011
rect 1638 -1027 1790 -1011
rect 1824 -1027 1862 -1011
rect 1896 -1027 2048 -1011
rect 2082 -1027 2120 -1011
rect 2154 -1027 2306 -1011
rect 2340 -1027 2378 -1011
rect 2412 -1027 2455 -993
rect 1489 -1033 2455 -1027
rect 2532 -945 2593 -713
rect 2715 -630 3423 -624
rect 2715 -664 2758 -630
rect 2792 -664 2830 -630
rect 2864 -664 3016 -630
rect 3050 -664 3088 -630
rect 3122 -664 3274 -630
rect 3308 -664 3346 -630
rect 3380 -664 3423 -630
rect 2715 -781 3423 -664
rect 2715 -833 2749 -781
rect 2801 -833 2813 -781
rect 2865 -833 2877 -781
rect 2929 -833 2945 -781
rect 2997 -833 3009 -781
rect 3061 -833 3073 -781
rect 3125 -833 3137 -781
rect 3189 -833 3205 -781
rect 3257 -833 3269 -781
rect 3321 -833 3333 -781
rect 3385 -833 3423 -781
rect 2715 -851 3423 -833
rect 3545 -630 4649 -624
rect 3545 -664 3726 -630
rect 3760 -643 3798 -630
rect 3832 -643 3984 -630
rect 4018 -643 4056 -630
rect 4090 -643 4242 -630
rect 4276 -643 4314 -630
rect 4348 -643 4500 -630
rect 4534 -643 4572 -630
rect 3789 -664 3798 -643
rect 3545 -695 3737 -664
rect 3789 -695 3801 -664
rect 3853 -695 3865 -643
rect 3917 -695 3933 -643
rect 4049 -664 4056 -643
rect 3985 -695 3997 -664
rect 4049 -695 4061 -664
rect 4113 -695 4223 -643
rect 4276 -664 4287 -643
rect 4348 -664 4351 -643
rect 4275 -695 4287 -664
rect 4339 -695 4351 -664
rect 4403 -695 4419 -643
rect 4471 -695 4483 -643
rect 4535 -695 4547 -643
rect 4606 -664 4649 -630
rect 4599 -695 4649 -664
rect 3545 -713 4649 -695
rect 4853 -625 5643 -587
rect 9210 -587 9589 -553
rect 9623 -587 9646 -553
rect 4853 -630 5231 -625
rect 4853 -664 4952 -630
rect 4986 -664 5024 -630
rect 5058 -659 5231 -630
rect 5265 -630 5643 -625
rect 5265 -659 5438 -630
rect 5058 -664 5438 -659
rect 5472 -664 5510 -630
rect 5544 -664 5643 -630
rect 4853 -697 5643 -664
rect 3545 -945 3606 -713
rect 4853 -731 5231 -697
rect 5265 -731 5643 -697
rect 5846 -630 6950 -624
rect 5846 -664 5889 -630
rect 5923 -643 5961 -630
rect 5995 -643 6147 -630
rect 6181 -643 6219 -630
rect 6253 -643 6405 -630
rect 6439 -643 6477 -630
rect 6511 -643 6663 -630
rect 6697 -643 6735 -630
rect 5846 -695 5896 -664
rect 5948 -695 5960 -643
rect 6012 -695 6024 -643
rect 6076 -695 6092 -643
rect 6144 -664 6147 -643
rect 6208 -664 6219 -643
rect 6144 -695 6156 -664
rect 6208 -695 6220 -664
rect 6272 -695 6382 -643
rect 6439 -664 6446 -643
rect 6434 -695 6446 -664
rect 6498 -695 6510 -664
rect 6562 -695 6578 -643
rect 6630 -695 6642 -643
rect 6697 -664 6706 -643
rect 6769 -664 6950 -630
rect 6694 -695 6706 -664
rect 6758 -695 6950 -664
rect 5846 -713 6950 -695
rect 2532 -993 3606 -945
rect 2532 -1027 2758 -993
rect 2792 -1027 2830 -993
rect 2864 -1027 3016 -993
rect 3050 -1027 3088 -993
rect 3122 -1027 3274 -993
rect 3308 -1027 3346 -993
rect 3380 -1027 3606 -993
rect 2532 -1033 3606 -1027
rect 3683 -781 4649 -763
rect 3683 -833 3737 -781
rect 3789 -833 3801 -781
rect 3853 -833 3865 -781
rect 3917 -833 3933 -781
rect 3985 -833 3997 -781
rect 4049 -833 4061 -781
rect 4113 -833 4223 -781
rect 4275 -833 4287 -781
rect 4339 -833 4351 -781
rect 4403 -833 4419 -781
rect 4471 -833 4483 -781
rect 4535 -833 4547 -781
rect 4599 -833 4649 -781
rect 3683 -959 4649 -833
rect 3683 -993 3737 -959
rect 3789 -993 3801 -959
rect 3683 -1027 3726 -993
rect 3789 -1011 3798 -993
rect 3853 -1011 3865 -959
rect 3917 -1011 3933 -959
rect 3985 -993 3997 -959
rect 4049 -993 4061 -959
rect 4049 -1011 4056 -993
rect 4113 -1011 4223 -959
rect 4275 -993 4287 -959
rect 4339 -993 4351 -959
rect 4276 -1011 4287 -993
rect 4348 -1011 4351 -993
rect 4403 -1011 4419 -959
rect 4471 -1011 4483 -959
rect 4535 -1011 4547 -959
rect 4599 -993 4649 -959
rect 3760 -1027 3798 -1011
rect 3832 -1027 3984 -1011
rect 4018 -1027 4056 -1011
rect 4090 -1027 4242 -1011
rect 4276 -1027 4314 -1011
rect 4348 -1027 4500 -1011
rect 4534 -1027 4572 -1011
rect 4606 -1027 4649 -993
rect 3683 -1033 4649 -1027
rect 4853 -769 5643 -731
rect 4853 -803 5231 -769
rect 5265 -803 5643 -769
rect 4853 -841 5643 -803
rect 4853 -875 5231 -841
rect 5265 -875 5643 -841
rect 4853 -913 5643 -875
rect 4853 -947 5231 -913
rect 5265 -947 5643 -913
rect 4853 -985 5643 -947
rect 4853 -993 5231 -985
rect 4853 -1027 4952 -993
rect 4986 -1027 5024 -993
rect 5058 -1019 5231 -993
rect 5265 -993 5643 -985
rect 5265 -1019 5438 -993
rect 5058 -1027 5438 -1019
rect 5472 -1027 5510 -993
rect 5544 -1027 5643 -993
rect 849 -1091 872 -1057
rect 906 -1091 1285 -1057
rect 4853 -1057 5643 -1027
rect 5846 -781 6812 -763
rect 5846 -833 5896 -781
rect 5948 -833 5960 -781
rect 6012 -833 6024 -781
rect 6076 -833 6092 -781
rect 6144 -833 6156 -781
rect 6208 -833 6220 -781
rect 6272 -833 6382 -781
rect 6434 -833 6446 -781
rect 6498 -833 6510 -781
rect 6562 -833 6578 -781
rect 6630 -833 6642 -781
rect 6694 -833 6706 -781
rect 6758 -833 6812 -781
rect 5846 -959 6812 -833
rect 5846 -993 5896 -959
rect 5846 -1027 5889 -993
rect 5948 -1011 5960 -959
rect 6012 -1011 6024 -959
rect 6076 -1011 6092 -959
rect 6144 -993 6156 -959
rect 6208 -993 6220 -959
rect 6144 -1011 6147 -993
rect 6208 -1011 6219 -993
rect 6272 -1011 6382 -959
rect 6434 -993 6446 -959
rect 6498 -993 6510 -959
rect 6439 -1011 6446 -993
rect 6562 -1011 6578 -959
rect 6630 -1011 6642 -959
rect 6694 -993 6706 -959
rect 6758 -993 6812 -959
rect 6697 -1011 6706 -993
rect 5923 -1027 5961 -1011
rect 5995 -1027 6147 -1011
rect 6181 -1027 6219 -1011
rect 6253 -1027 6405 -1011
rect 6439 -1027 6477 -1011
rect 6511 -1027 6663 -1011
rect 6697 -1027 6735 -1011
rect 6769 -1027 6812 -993
rect 5846 -1033 6812 -1027
rect 6889 -945 6950 -713
rect 7072 -630 7780 -624
rect 7072 -664 7115 -630
rect 7149 -664 7187 -630
rect 7221 -664 7373 -630
rect 7407 -664 7445 -630
rect 7479 -664 7631 -630
rect 7665 -664 7703 -630
rect 7737 -664 7780 -630
rect 7072 -781 7780 -664
rect 7072 -833 7110 -781
rect 7162 -833 7174 -781
rect 7226 -833 7238 -781
rect 7290 -833 7306 -781
rect 7358 -833 7370 -781
rect 7422 -833 7434 -781
rect 7486 -833 7498 -781
rect 7550 -833 7566 -781
rect 7618 -833 7630 -781
rect 7682 -833 7694 -781
rect 7746 -833 7780 -781
rect 7072 -851 7780 -833
rect 7902 -630 9006 -624
rect 7902 -664 8083 -630
rect 8117 -643 8155 -630
rect 8189 -643 8341 -630
rect 8375 -643 8413 -630
rect 8447 -643 8599 -630
rect 8633 -643 8671 -630
rect 8705 -643 8857 -630
rect 8891 -643 8929 -630
rect 8146 -664 8155 -643
rect 7902 -695 8094 -664
rect 8146 -695 8158 -664
rect 8210 -695 8222 -643
rect 8274 -695 8290 -643
rect 8406 -664 8413 -643
rect 8342 -695 8354 -664
rect 8406 -695 8418 -664
rect 8470 -695 8580 -643
rect 8633 -664 8644 -643
rect 8705 -664 8708 -643
rect 8632 -695 8644 -664
rect 8696 -695 8708 -664
rect 8760 -695 8776 -643
rect 8828 -695 8840 -643
rect 8892 -695 8904 -643
rect 8963 -664 9006 -630
rect 8956 -695 9006 -664
rect 7902 -713 9006 -695
rect 9210 -625 9646 -587
rect 9210 -630 9589 -625
rect 9210 -664 9309 -630
rect 9343 -664 9381 -630
rect 9415 -659 9589 -630
rect 9623 -659 9646 -625
rect 9415 -664 9646 -659
rect 9210 -697 9646 -664
rect 7902 -945 7963 -713
rect 9210 -731 9589 -697
rect 9623 -731 9646 -697
rect 6889 -993 7963 -945
rect 6889 -1027 7115 -993
rect 7149 -1027 7187 -993
rect 7221 -1027 7373 -993
rect 7407 -1027 7445 -993
rect 7479 -1027 7631 -993
rect 7665 -1027 7703 -993
rect 7737 -1027 7963 -993
rect 6889 -1033 7963 -1027
rect 8040 -781 9006 -763
rect 8040 -833 8094 -781
rect 8146 -833 8158 -781
rect 8210 -833 8222 -781
rect 8274 -833 8290 -781
rect 8342 -833 8354 -781
rect 8406 -833 8418 -781
rect 8470 -833 8580 -781
rect 8632 -833 8644 -781
rect 8696 -833 8708 -781
rect 8760 -833 8776 -781
rect 8828 -833 8840 -781
rect 8892 -833 8904 -781
rect 8956 -833 9006 -781
rect 8040 -959 9006 -833
rect 8040 -993 8094 -959
rect 8146 -993 8158 -959
rect 8040 -1027 8083 -993
rect 8146 -1011 8155 -993
rect 8210 -1011 8222 -959
rect 8274 -1011 8290 -959
rect 8342 -993 8354 -959
rect 8406 -993 8418 -959
rect 8406 -1011 8413 -993
rect 8470 -1011 8580 -959
rect 8632 -993 8644 -959
rect 8696 -993 8708 -959
rect 8633 -1011 8644 -993
rect 8705 -1011 8708 -993
rect 8760 -1011 8776 -959
rect 8828 -1011 8840 -959
rect 8892 -1011 8904 -959
rect 8956 -993 9006 -959
rect 8117 -1027 8155 -1011
rect 8189 -1027 8341 -1011
rect 8375 -1027 8413 -1011
rect 8447 -1027 8599 -1011
rect 8633 -1027 8671 -1011
rect 8705 -1027 8857 -1011
rect 8891 -1027 8929 -1011
rect 8963 -1027 9006 -993
rect 8040 -1033 9006 -1027
rect 9210 -769 9646 -731
rect 9210 -803 9589 -769
rect 9623 -803 9646 -769
rect 9210 -841 9646 -803
rect 9210 -875 9589 -841
rect 9623 -875 9646 -841
rect 9210 -913 9646 -875
rect 9210 -947 9589 -913
rect 9623 -947 9646 -913
rect 9210 -985 9646 -947
rect 9210 -993 9589 -985
rect 9210 -1027 9309 -993
rect 9343 -1027 9381 -993
rect 9415 -1019 9589 -993
rect 9623 -1019 9646 -985
rect 9415 -1027 9646 -1019
rect 849 -1121 1285 -1091
rect 849 -1129 987 -1121
rect 849 -1163 872 -1129
rect 906 -1155 987 -1129
rect 1021 -1155 1245 -1121
rect 1279 -1155 1285 -1121
rect 906 -1163 1285 -1155
rect 849 -1193 1285 -1163
rect 849 -1201 987 -1193
rect 849 -1235 872 -1201
rect 906 -1227 987 -1201
rect 1021 -1227 1245 -1193
rect 1279 -1227 1285 -1193
rect 906 -1235 1285 -1227
rect 849 -1273 1285 -1235
rect 849 -1307 872 -1273
rect 906 -1307 1285 -1273
rect 849 -1345 1285 -1307
rect 849 -1379 872 -1345
rect 906 -1379 1285 -1345
rect 849 -1417 1285 -1379
rect 1433 -1121 1479 -1074
rect 1433 -1155 1439 -1121
rect 1473 -1155 1479 -1121
rect 1433 -1193 1479 -1155
rect 1433 -1227 1439 -1193
rect 1473 -1227 1479 -1193
rect 1433 -1401 1479 -1227
rect 1691 -1121 1737 -1074
rect 1691 -1155 1697 -1121
rect 1731 -1155 1737 -1121
rect 1691 -1193 1737 -1155
rect 1691 -1227 1697 -1193
rect 1731 -1227 1737 -1193
rect 849 -1451 872 -1417
rect 906 -1451 1285 -1417
rect 849 -1489 1285 -1451
rect 1360 -1409 1556 -1401
rect 1360 -1461 1367 -1409
rect 1419 -1461 1431 -1409
rect 1483 -1461 1495 -1409
rect 1547 -1461 1556 -1409
rect 1360 -1471 1556 -1461
rect 849 -1523 872 -1489
rect 906 -1523 1285 -1489
rect 849 -1561 1285 -1523
rect 849 -1595 872 -1561
rect 906 -1595 1285 -1561
rect 849 -1633 1285 -1595
rect 849 -1667 872 -1633
rect 906 -1667 1285 -1633
rect 849 -1705 1285 -1667
rect 849 -1739 872 -1705
rect 906 -1739 1285 -1705
rect 849 -1777 1285 -1739
rect 849 -1811 872 -1777
rect 906 -1811 1285 -1777
rect 849 -1849 1285 -1811
rect 849 -1883 872 -1849
rect 906 -1883 1285 -1849
rect 849 -1921 1285 -1883
rect 849 -1955 872 -1921
rect 906 -1955 1285 -1921
rect 849 -1993 1285 -1955
rect 849 -2027 872 -1993
rect 906 -2027 1285 -1993
rect 849 -2065 1285 -2027
rect 849 -2099 872 -2065
rect 906 -2077 1285 -2065
rect 906 -2099 987 -2077
rect 849 -2111 987 -2099
rect 1021 -2111 1245 -2077
rect 1279 -2111 1285 -2077
rect 849 -2137 1285 -2111
rect 849 -2171 872 -2137
rect 906 -2149 1285 -2137
rect 906 -2171 987 -2149
rect 849 -2183 987 -2171
rect 1021 -2183 1245 -2149
rect 1279 -2183 1285 -2149
rect 849 -2209 1285 -2183
rect 849 -2243 872 -2209
rect 906 -2243 1285 -2209
rect 1433 -2077 1479 -1471
rect 1691 -1702 1737 -1227
rect 1949 -1121 1995 -1074
rect 1949 -1155 1955 -1121
rect 1989 -1155 1995 -1121
rect 1949 -1193 1995 -1155
rect 1949 -1227 1955 -1193
rect 1989 -1227 1995 -1193
rect 1949 -1401 1995 -1227
rect 2207 -1121 2253 -1074
rect 2207 -1155 2213 -1121
rect 2247 -1155 2253 -1121
rect 2207 -1193 2253 -1155
rect 2207 -1227 2213 -1193
rect 2247 -1227 2253 -1193
rect 1875 -1409 2071 -1401
rect 1875 -1461 1882 -1409
rect 1934 -1461 1946 -1409
rect 1998 -1461 2010 -1409
rect 2062 -1461 2071 -1409
rect 1875 -1471 2071 -1461
rect 1618 -1710 1814 -1702
rect 1618 -1762 1625 -1710
rect 1677 -1762 1689 -1710
rect 1741 -1762 1753 -1710
rect 1805 -1762 1814 -1710
rect 1618 -1772 1814 -1762
rect 1433 -2111 1439 -2077
rect 1473 -2111 1479 -2077
rect 1433 -2149 1479 -2111
rect 1433 -2183 1439 -2149
rect 1473 -2183 1479 -2149
rect 1433 -2230 1479 -2183
rect 1691 -2077 1737 -1772
rect 1691 -2111 1697 -2077
rect 1731 -2111 1737 -2077
rect 1691 -2149 1737 -2111
rect 1691 -2183 1697 -2149
rect 1731 -2183 1737 -2149
rect 1691 -2230 1737 -2183
rect 1949 -2077 1995 -1471
rect 2207 -1702 2253 -1227
rect 2465 -1121 2511 -1074
rect 2465 -1155 2471 -1121
rect 2505 -1155 2511 -1121
rect 2465 -1193 2511 -1155
rect 2465 -1227 2471 -1193
rect 2505 -1227 2511 -1193
rect 2465 -1401 2511 -1227
rect 2659 -1121 2705 -1074
rect 2659 -1155 2665 -1121
rect 2699 -1155 2705 -1121
rect 2659 -1193 2705 -1155
rect 2659 -1227 2665 -1193
rect 2699 -1227 2705 -1193
rect 2392 -1409 2588 -1401
rect 2392 -1461 2399 -1409
rect 2451 -1461 2463 -1409
rect 2515 -1461 2527 -1409
rect 2579 -1461 2588 -1409
rect 2392 -1471 2588 -1461
rect 2135 -1710 2331 -1702
rect 2135 -1762 2142 -1710
rect 2194 -1762 2206 -1710
rect 2258 -1762 2270 -1710
rect 2322 -1762 2331 -1710
rect 2135 -1772 2331 -1762
rect 1949 -2111 1955 -2077
rect 1989 -2111 1995 -2077
rect 1949 -2149 1995 -2111
rect 1949 -2183 1955 -2149
rect 1989 -2183 1995 -2149
rect 1949 -2230 1995 -2183
rect 2207 -2077 2253 -1772
rect 2207 -2111 2213 -2077
rect 2247 -2111 2253 -2077
rect 2207 -2149 2253 -2111
rect 2207 -2183 2213 -2149
rect 2247 -2183 2253 -2149
rect 2207 -2230 2253 -2183
rect 2465 -2077 2511 -1471
rect 2659 -1846 2705 -1227
rect 2917 -1121 2963 -1074
rect 2917 -1155 2923 -1121
rect 2957 -1155 2963 -1121
rect 2917 -1193 2963 -1155
rect 2917 -1227 2923 -1193
rect 2957 -1227 2963 -1193
rect 2917 -1541 2963 -1227
rect 3175 -1121 3221 -1074
rect 3175 -1155 3181 -1121
rect 3215 -1155 3221 -1121
rect 3175 -1193 3221 -1155
rect 3175 -1227 3181 -1193
rect 3215 -1227 3221 -1193
rect 2840 -1549 3036 -1541
rect 2840 -1601 2849 -1549
rect 2901 -1601 2913 -1549
rect 2965 -1601 2977 -1549
rect 3029 -1601 3036 -1549
rect 2840 -1611 3036 -1601
rect 2582 -1854 2778 -1846
rect 2582 -1906 2591 -1854
rect 2643 -1906 2655 -1854
rect 2707 -1906 2719 -1854
rect 2771 -1906 2778 -1854
rect 2582 -1916 2778 -1906
rect 2465 -2111 2471 -2077
rect 2505 -2111 2511 -2077
rect 2465 -2149 2511 -2111
rect 2465 -2183 2471 -2149
rect 2505 -2183 2511 -2149
rect 2465 -2230 2511 -2183
rect 2659 -2077 2705 -1916
rect 2659 -2111 2665 -2077
rect 2699 -2111 2705 -2077
rect 2659 -2149 2705 -2111
rect 2659 -2183 2665 -2149
rect 2699 -2183 2705 -2149
rect 2659 -2230 2705 -2183
rect 2917 -2077 2963 -1611
rect 3175 -1846 3221 -1227
rect 3433 -1121 3479 -1074
rect 3433 -1155 3439 -1121
rect 3473 -1155 3479 -1121
rect 3433 -1193 3479 -1155
rect 3433 -1227 3439 -1193
rect 3473 -1227 3479 -1193
rect 3433 -1541 3479 -1227
rect 3627 -1121 3673 -1074
rect 3627 -1155 3633 -1121
rect 3667 -1155 3673 -1121
rect 3627 -1193 3673 -1155
rect 3627 -1227 3633 -1193
rect 3667 -1227 3673 -1193
rect 3627 -1401 3673 -1227
rect 3885 -1121 3931 -1074
rect 3885 -1155 3891 -1121
rect 3925 -1155 3931 -1121
rect 3885 -1193 3931 -1155
rect 3885 -1227 3891 -1193
rect 3925 -1227 3931 -1193
rect 3552 -1409 3748 -1401
rect 3552 -1461 3559 -1409
rect 3611 -1461 3623 -1409
rect 3675 -1461 3687 -1409
rect 3739 -1461 3748 -1409
rect 3552 -1471 3748 -1461
rect 3357 -1549 3553 -1541
rect 3357 -1601 3366 -1549
rect 3418 -1601 3430 -1549
rect 3482 -1601 3494 -1549
rect 3546 -1601 3553 -1549
rect 3357 -1611 3553 -1601
rect 3099 -1854 3295 -1846
rect 3099 -1906 3108 -1854
rect 3160 -1906 3172 -1854
rect 3224 -1906 3236 -1854
rect 3288 -1906 3295 -1854
rect 3099 -1916 3295 -1906
rect 2917 -2111 2923 -2077
rect 2957 -2111 2963 -2077
rect 2917 -2149 2963 -2111
rect 2917 -2183 2923 -2149
rect 2957 -2183 2963 -2149
rect 2917 -2230 2963 -2183
rect 3175 -2077 3221 -1916
rect 3175 -2111 3181 -2077
rect 3215 -2111 3221 -2077
rect 3175 -2149 3221 -2111
rect 3175 -2183 3181 -2149
rect 3215 -2183 3221 -2149
rect 3175 -2230 3221 -2183
rect 3433 -2077 3479 -1611
rect 3433 -2111 3439 -2077
rect 3473 -2111 3479 -2077
rect 3433 -2149 3479 -2111
rect 3433 -2183 3439 -2149
rect 3473 -2183 3479 -2149
rect 3433 -2230 3479 -2183
rect 3627 -2077 3673 -1471
rect 3885 -1702 3931 -1227
rect 4143 -1121 4189 -1074
rect 4143 -1155 4149 -1121
rect 4183 -1155 4189 -1121
rect 4143 -1193 4189 -1155
rect 4143 -1227 4149 -1193
rect 4183 -1227 4189 -1193
rect 4143 -1401 4189 -1227
rect 4401 -1121 4447 -1074
rect 4401 -1155 4407 -1121
rect 4441 -1155 4447 -1121
rect 4401 -1193 4447 -1155
rect 4401 -1227 4407 -1193
rect 4441 -1227 4447 -1193
rect 4069 -1409 4265 -1401
rect 4069 -1461 4076 -1409
rect 4128 -1461 4140 -1409
rect 4192 -1461 4204 -1409
rect 4256 -1461 4265 -1409
rect 4069 -1471 4265 -1461
rect 3812 -1710 4008 -1702
rect 3812 -1762 3819 -1710
rect 3871 -1762 3883 -1710
rect 3935 -1762 3947 -1710
rect 3999 -1762 4008 -1710
rect 3812 -1772 4008 -1762
rect 3627 -2111 3633 -2077
rect 3667 -2111 3673 -2077
rect 3627 -2149 3673 -2111
rect 3627 -2183 3633 -2149
rect 3667 -2183 3673 -2149
rect 3627 -2230 3673 -2183
rect 3885 -2077 3931 -1772
rect 3885 -2111 3891 -2077
rect 3925 -2111 3931 -2077
rect 3885 -2149 3931 -2111
rect 3885 -2183 3891 -2149
rect 3925 -2183 3931 -2149
rect 3885 -2230 3931 -2183
rect 4143 -2077 4189 -1471
rect 4401 -1702 4447 -1227
rect 4659 -1121 4705 -1074
rect 4659 -1155 4665 -1121
rect 4699 -1155 4705 -1121
rect 4659 -1193 4705 -1155
rect 4659 -1227 4665 -1193
rect 4699 -1227 4705 -1193
rect 4659 -1401 4705 -1227
rect 4853 -1091 5231 -1057
rect 5265 -1091 5643 -1057
rect 9210 -1057 9646 -1027
rect 4853 -1121 5643 -1091
rect 4853 -1155 4859 -1121
rect 4893 -1155 5117 -1121
rect 5151 -1129 5345 -1121
rect 5151 -1155 5231 -1129
rect 4853 -1163 5231 -1155
rect 5265 -1155 5345 -1129
rect 5379 -1155 5603 -1121
rect 5637 -1155 5643 -1121
rect 5265 -1163 5643 -1155
rect 4853 -1193 5643 -1163
rect 4853 -1227 4859 -1193
rect 4893 -1227 5117 -1193
rect 5151 -1201 5345 -1193
rect 5151 -1227 5231 -1201
rect 4853 -1235 5231 -1227
rect 5265 -1227 5345 -1201
rect 5379 -1227 5603 -1193
rect 5637 -1227 5643 -1193
rect 5265 -1235 5643 -1227
rect 4853 -1273 5643 -1235
rect 4853 -1307 5231 -1273
rect 5265 -1307 5643 -1273
rect 4853 -1345 5643 -1307
rect 4853 -1379 5231 -1345
rect 5265 -1379 5643 -1345
rect 4586 -1409 4782 -1401
rect 4586 -1461 4593 -1409
rect 4645 -1461 4657 -1409
rect 4709 -1461 4721 -1409
rect 4773 -1461 4782 -1409
rect 4586 -1471 4782 -1461
rect 4853 -1417 5643 -1379
rect 5790 -1121 5836 -1074
rect 5790 -1155 5796 -1121
rect 5830 -1155 5836 -1121
rect 5790 -1193 5836 -1155
rect 5790 -1227 5796 -1193
rect 5830 -1227 5836 -1193
rect 5790 -1401 5836 -1227
rect 6048 -1121 6094 -1074
rect 6048 -1155 6054 -1121
rect 6088 -1155 6094 -1121
rect 6048 -1193 6094 -1155
rect 6048 -1227 6054 -1193
rect 6088 -1227 6094 -1193
rect 4853 -1451 5231 -1417
rect 5265 -1451 5643 -1417
rect 4329 -1710 4525 -1702
rect 4329 -1762 4336 -1710
rect 4388 -1762 4400 -1710
rect 4452 -1762 4464 -1710
rect 4516 -1762 4525 -1710
rect 4329 -1772 4525 -1762
rect 4143 -2111 4149 -2077
rect 4183 -2111 4189 -2077
rect 4143 -2149 4189 -2111
rect 4143 -2183 4149 -2149
rect 4183 -2183 4189 -2149
rect 4143 -2230 4189 -2183
rect 4401 -2077 4447 -1772
rect 4401 -2111 4407 -2077
rect 4441 -2111 4447 -2077
rect 4401 -2149 4447 -2111
rect 4401 -2183 4407 -2149
rect 4441 -2183 4447 -2149
rect 4401 -2230 4447 -2183
rect 4659 -2077 4705 -1471
rect 4659 -2111 4665 -2077
rect 4699 -2111 4705 -2077
rect 4659 -2149 4705 -2111
rect 4659 -2183 4665 -2149
rect 4699 -2183 4705 -2149
rect 4659 -2230 4705 -2183
rect 4853 -1489 5643 -1451
rect 5713 -1409 5909 -1401
rect 5713 -1461 5722 -1409
rect 5774 -1461 5786 -1409
rect 5838 -1461 5850 -1409
rect 5902 -1461 5909 -1409
rect 5713 -1471 5909 -1461
rect 4853 -1523 5231 -1489
rect 5265 -1523 5643 -1489
rect 4853 -1561 5643 -1523
rect 4853 -1595 5231 -1561
rect 5265 -1595 5643 -1561
rect 4853 -1633 5643 -1595
rect 4853 -1667 5231 -1633
rect 5265 -1667 5643 -1633
rect 4853 -1705 5643 -1667
rect 4853 -1739 5231 -1705
rect 5265 -1739 5643 -1705
rect 4853 -1777 5643 -1739
rect 4853 -1811 5231 -1777
rect 5265 -1811 5643 -1777
rect 4853 -1849 5643 -1811
rect 4853 -1883 5231 -1849
rect 5265 -1883 5643 -1849
rect 4853 -1921 5643 -1883
rect 4853 -1955 5231 -1921
rect 5265 -1955 5643 -1921
rect 4853 -1993 5643 -1955
rect 4853 -2027 5231 -1993
rect 5265 -2027 5643 -1993
rect 4853 -2065 5643 -2027
rect 4853 -2077 5231 -2065
rect 4853 -2111 4859 -2077
rect 4893 -2111 5117 -2077
rect 5151 -2099 5231 -2077
rect 5265 -2077 5643 -2065
rect 5265 -2099 5345 -2077
rect 5151 -2111 5345 -2099
rect 5379 -2111 5603 -2077
rect 5637 -2111 5643 -2077
rect 4853 -2137 5643 -2111
rect 4853 -2149 5231 -2137
rect 4853 -2183 4859 -2149
rect 4893 -2183 5117 -2149
rect 5151 -2171 5231 -2149
rect 5265 -2149 5643 -2137
rect 5265 -2171 5345 -2149
rect 5151 -2183 5345 -2171
rect 5379 -2183 5603 -2149
rect 5637 -2183 5643 -2149
rect 4853 -2209 5643 -2183
rect 849 -2277 1285 -2243
rect 4853 -2243 5231 -2209
rect 5265 -2243 5643 -2209
rect 5790 -2077 5836 -1471
rect 6048 -1702 6094 -1227
rect 6306 -1121 6352 -1074
rect 6306 -1155 6312 -1121
rect 6346 -1155 6352 -1121
rect 6306 -1193 6352 -1155
rect 6306 -1227 6312 -1193
rect 6346 -1227 6352 -1193
rect 6306 -1401 6352 -1227
rect 6564 -1121 6610 -1074
rect 6564 -1155 6570 -1121
rect 6604 -1155 6610 -1121
rect 6564 -1193 6610 -1155
rect 6564 -1227 6570 -1193
rect 6604 -1227 6610 -1193
rect 6230 -1409 6426 -1401
rect 6230 -1461 6239 -1409
rect 6291 -1461 6303 -1409
rect 6355 -1461 6367 -1409
rect 6419 -1461 6426 -1409
rect 6230 -1471 6426 -1461
rect 5970 -1710 6166 -1702
rect 5970 -1762 5979 -1710
rect 6031 -1762 6043 -1710
rect 6095 -1762 6107 -1710
rect 6159 -1762 6166 -1710
rect 5970 -1772 6166 -1762
rect 5790 -2111 5796 -2077
rect 5830 -2111 5836 -2077
rect 5790 -2149 5836 -2111
rect 5790 -2183 5796 -2149
rect 5830 -2183 5836 -2149
rect 5790 -2230 5836 -2183
rect 6048 -2077 6094 -1772
rect 6048 -2111 6054 -2077
rect 6088 -2111 6094 -2077
rect 6048 -2149 6094 -2111
rect 6048 -2183 6054 -2149
rect 6088 -2183 6094 -2149
rect 6048 -2230 6094 -2183
rect 6306 -2077 6352 -1471
rect 6564 -1702 6610 -1227
rect 6822 -1121 6868 -1074
rect 6822 -1155 6828 -1121
rect 6862 -1155 6868 -1121
rect 6822 -1193 6868 -1155
rect 6822 -1227 6828 -1193
rect 6862 -1227 6868 -1193
rect 6822 -1401 6868 -1227
rect 7016 -1121 7062 -1074
rect 7016 -1155 7022 -1121
rect 7056 -1155 7062 -1121
rect 7016 -1193 7062 -1155
rect 7016 -1227 7022 -1193
rect 7056 -1227 7062 -1193
rect 6747 -1409 6943 -1401
rect 6747 -1461 6756 -1409
rect 6808 -1461 6820 -1409
rect 6872 -1461 6884 -1409
rect 6936 -1461 6943 -1409
rect 6747 -1471 6943 -1461
rect 6487 -1710 6683 -1702
rect 6487 -1762 6496 -1710
rect 6548 -1762 6560 -1710
rect 6612 -1762 6624 -1710
rect 6676 -1762 6683 -1710
rect 6487 -1772 6683 -1762
rect 6306 -2111 6312 -2077
rect 6346 -2111 6352 -2077
rect 6306 -2149 6352 -2111
rect 6306 -2183 6312 -2149
rect 6346 -2183 6352 -2149
rect 6306 -2230 6352 -2183
rect 6564 -2077 6610 -1772
rect 6564 -2111 6570 -2077
rect 6604 -2111 6610 -2077
rect 6564 -2149 6610 -2111
rect 6564 -2183 6570 -2149
rect 6604 -2183 6610 -2149
rect 6564 -2230 6610 -2183
rect 6822 -2077 6868 -1471
rect 7016 -1541 7062 -1227
rect 7274 -1121 7320 -1074
rect 7274 -1155 7280 -1121
rect 7314 -1155 7320 -1121
rect 7274 -1193 7320 -1155
rect 7274 -1227 7280 -1193
rect 7314 -1227 7320 -1193
rect 6942 -1549 7138 -1541
rect 6942 -1601 6949 -1549
rect 7001 -1601 7013 -1549
rect 7065 -1601 7077 -1549
rect 7129 -1601 7138 -1549
rect 6942 -1611 7138 -1601
rect 6822 -2111 6828 -2077
rect 6862 -2111 6868 -2077
rect 6822 -2149 6868 -2111
rect 6822 -2183 6828 -2149
rect 6862 -2183 6868 -2149
rect 6822 -2230 6868 -2183
rect 7016 -2077 7062 -1611
rect 7274 -1846 7320 -1227
rect 7532 -1121 7578 -1074
rect 7532 -1155 7538 -1121
rect 7572 -1155 7578 -1121
rect 7532 -1193 7578 -1155
rect 7532 -1227 7538 -1193
rect 7572 -1227 7578 -1193
rect 7532 -1541 7578 -1227
rect 7790 -1121 7836 -1074
rect 7790 -1155 7796 -1121
rect 7830 -1155 7836 -1121
rect 7790 -1193 7836 -1155
rect 7790 -1227 7796 -1193
rect 7830 -1227 7836 -1193
rect 7459 -1549 7655 -1541
rect 7459 -1601 7466 -1549
rect 7518 -1601 7530 -1549
rect 7582 -1601 7594 -1549
rect 7646 -1601 7655 -1549
rect 7459 -1611 7655 -1601
rect 7200 -1854 7396 -1846
rect 7200 -1906 7207 -1854
rect 7259 -1906 7271 -1854
rect 7323 -1906 7335 -1854
rect 7387 -1906 7396 -1854
rect 7200 -1916 7396 -1906
rect 7016 -2111 7022 -2077
rect 7056 -2111 7062 -2077
rect 7016 -2149 7062 -2111
rect 7016 -2183 7022 -2149
rect 7056 -2183 7062 -2149
rect 7016 -2230 7062 -2183
rect 7274 -2077 7320 -1916
rect 7274 -2111 7280 -2077
rect 7314 -2111 7320 -2077
rect 7274 -2149 7320 -2111
rect 7274 -2183 7280 -2149
rect 7314 -2183 7320 -2149
rect 7274 -2230 7320 -2183
rect 7532 -2077 7578 -1611
rect 7790 -1846 7836 -1227
rect 7984 -1121 8030 -1074
rect 7984 -1155 7990 -1121
rect 8024 -1155 8030 -1121
rect 7984 -1193 8030 -1155
rect 7984 -1227 7990 -1193
rect 8024 -1227 8030 -1193
rect 7984 -1401 8030 -1227
rect 8242 -1121 8288 -1074
rect 8242 -1155 8248 -1121
rect 8282 -1155 8288 -1121
rect 8242 -1193 8288 -1155
rect 8242 -1227 8248 -1193
rect 8282 -1227 8288 -1193
rect 7907 -1409 8103 -1401
rect 7907 -1461 7916 -1409
rect 7968 -1461 7980 -1409
rect 8032 -1461 8044 -1409
rect 8096 -1461 8103 -1409
rect 7907 -1471 8103 -1461
rect 7717 -1854 7913 -1846
rect 7717 -1906 7724 -1854
rect 7776 -1906 7788 -1854
rect 7840 -1906 7852 -1854
rect 7904 -1906 7913 -1854
rect 7717 -1916 7913 -1906
rect 7532 -2111 7538 -2077
rect 7572 -2111 7578 -2077
rect 7532 -2149 7578 -2111
rect 7532 -2183 7538 -2149
rect 7572 -2183 7578 -2149
rect 7532 -2230 7578 -2183
rect 7790 -2077 7836 -1916
rect 7790 -2111 7796 -2077
rect 7830 -2111 7836 -2077
rect 7790 -2149 7836 -2111
rect 7790 -2183 7796 -2149
rect 7830 -2183 7836 -2149
rect 7790 -2230 7836 -2183
rect 7984 -2077 8030 -1471
rect 8242 -1702 8288 -1227
rect 8500 -1121 8546 -1074
rect 8500 -1155 8506 -1121
rect 8540 -1155 8546 -1121
rect 8500 -1193 8546 -1155
rect 8500 -1227 8506 -1193
rect 8540 -1227 8546 -1193
rect 8500 -1401 8546 -1227
rect 8758 -1121 8804 -1074
rect 8758 -1155 8764 -1121
rect 8798 -1155 8804 -1121
rect 8758 -1193 8804 -1155
rect 8758 -1227 8764 -1193
rect 8798 -1227 8804 -1193
rect 8425 -1409 8621 -1401
rect 8425 -1461 8434 -1409
rect 8486 -1461 8498 -1409
rect 8550 -1461 8562 -1409
rect 8614 -1461 8621 -1409
rect 8425 -1471 8621 -1461
rect 8164 -1710 8360 -1702
rect 8164 -1762 8173 -1710
rect 8225 -1762 8237 -1710
rect 8289 -1762 8301 -1710
rect 8353 -1762 8360 -1710
rect 8164 -1772 8360 -1762
rect 7984 -2111 7990 -2077
rect 8024 -2111 8030 -2077
rect 7984 -2149 8030 -2111
rect 7984 -2183 7990 -2149
rect 8024 -2183 8030 -2149
rect 7984 -2230 8030 -2183
rect 8242 -2077 8288 -1772
rect 8242 -2111 8248 -2077
rect 8282 -2111 8288 -2077
rect 8242 -2149 8288 -2111
rect 8242 -2183 8248 -2149
rect 8282 -2183 8288 -2149
rect 8242 -2230 8288 -2183
rect 8500 -2077 8546 -1471
rect 8758 -1702 8804 -1227
rect 9016 -1121 9062 -1074
rect 9016 -1155 9022 -1121
rect 9056 -1155 9062 -1121
rect 9016 -1193 9062 -1155
rect 9016 -1227 9022 -1193
rect 9056 -1227 9062 -1193
rect 9016 -1401 9062 -1227
rect 9210 -1091 9589 -1057
rect 9623 -1091 9646 -1057
rect 9210 -1121 9646 -1091
rect 9210 -1155 9216 -1121
rect 9250 -1155 9474 -1121
rect 9508 -1129 9646 -1121
rect 9508 -1155 9589 -1129
rect 9210 -1163 9589 -1155
rect 9623 -1163 9646 -1129
rect 9210 -1193 9646 -1163
rect 9210 -1227 9216 -1193
rect 9250 -1227 9474 -1193
rect 9508 -1201 9646 -1193
rect 9508 -1227 9589 -1201
rect 9210 -1235 9589 -1227
rect 9623 -1235 9646 -1201
rect 9210 -1273 9646 -1235
rect 9210 -1307 9589 -1273
rect 9623 -1307 9646 -1273
rect 9210 -1345 9646 -1307
rect 9210 -1379 9589 -1345
rect 9623 -1379 9646 -1345
rect 8940 -1409 9136 -1401
rect 8940 -1461 8949 -1409
rect 9001 -1461 9013 -1409
rect 9065 -1461 9077 -1409
rect 9129 -1461 9136 -1409
rect 8940 -1471 9136 -1461
rect 9210 -1417 9646 -1379
rect 9210 -1451 9589 -1417
rect 9623 -1451 9646 -1417
rect 8682 -1710 8878 -1702
rect 8682 -1762 8691 -1710
rect 8743 -1762 8755 -1710
rect 8807 -1762 8819 -1710
rect 8871 -1762 8878 -1710
rect 8682 -1772 8878 -1762
rect 8500 -2111 8506 -2077
rect 8540 -2111 8546 -2077
rect 8500 -2149 8546 -2111
rect 8500 -2183 8506 -2149
rect 8540 -2183 8546 -2149
rect 8500 -2230 8546 -2183
rect 8758 -2077 8804 -1772
rect 8758 -2111 8764 -2077
rect 8798 -2111 8804 -2077
rect 8758 -2149 8804 -2111
rect 8758 -2183 8764 -2149
rect 8798 -2183 8804 -2149
rect 8758 -2230 8804 -2183
rect 9016 -2077 9062 -1471
rect 9016 -2111 9022 -2077
rect 9056 -2111 9062 -2077
rect 9016 -2149 9062 -2111
rect 9016 -2183 9022 -2149
rect 9056 -2183 9062 -2149
rect 9016 -2230 9062 -2183
rect 9210 -1489 9646 -1451
rect 9210 -1523 9589 -1489
rect 9623 -1523 9646 -1489
rect 9210 -1561 9646 -1523
rect 9210 -1595 9589 -1561
rect 9623 -1595 9646 -1561
rect 9210 -1633 9646 -1595
rect 9210 -1667 9589 -1633
rect 9623 -1667 9646 -1633
rect 9210 -1705 9646 -1667
rect 9210 -1739 9589 -1705
rect 9623 -1739 9646 -1705
rect 9210 -1777 9646 -1739
rect 9210 -1811 9589 -1777
rect 9623 -1811 9646 -1777
rect 9210 -1849 9646 -1811
rect 9210 -1883 9589 -1849
rect 9623 -1883 9646 -1849
rect 9210 -1921 9646 -1883
rect 9210 -1955 9589 -1921
rect 9623 -1955 9646 -1921
rect 9210 -1993 9646 -1955
rect 9210 -2027 9589 -1993
rect 9623 -2027 9646 -1993
rect 9210 -2065 9646 -2027
rect 9210 -2077 9589 -2065
rect 9210 -2111 9216 -2077
rect 9250 -2111 9474 -2077
rect 9508 -2099 9589 -2077
rect 9623 -2099 9646 -2065
rect 9508 -2111 9646 -2099
rect 9210 -2137 9646 -2111
rect 9210 -2149 9589 -2137
rect 9210 -2183 9216 -2149
rect 9250 -2183 9474 -2149
rect 9508 -2171 9589 -2149
rect 9623 -2171 9646 -2137
rect 9508 -2183 9646 -2171
rect 9210 -2209 9646 -2183
rect 849 -2281 1080 -2277
rect 849 -2315 872 -2281
rect 906 -2311 1080 -2281
rect 1114 -2311 1152 -2277
rect 1186 -2311 1285 -2277
rect 906 -2315 1285 -2311
rect 849 -2353 1285 -2315
rect 849 -2387 872 -2353
rect 906 -2387 1285 -2353
rect 1489 -2277 2593 -2271
rect 1489 -2311 1532 -2277
rect 1566 -2290 1604 -2277
rect 1638 -2290 1790 -2277
rect 1824 -2290 1862 -2277
rect 1896 -2290 2048 -2277
rect 2082 -2290 2120 -2277
rect 2154 -2290 2306 -2277
rect 2340 -2290 2378 -2277
rect 1489 -2342 1539 -2311
rect 1591 -2342 1603 -2290
rect 1655 -2342 1667 -2290
rect 1719 -2342 1735 -2290
rect 1787 -2311 1790 -2290
rect 1851 -2311 1862 -2290
rect 1787 -2342 1799 -2311
rect 1851 -2342 1863 -2311
rect 1915 -2342 2025 -2290
rect 2082 -2311 2089 -2290
rect 2077 -2342 2089 -2311
rect 2141 -2342 2153 -2311
rect 2205 -2342 2221 -2290
rect 2273 -2342 2285 -2290
rect 2340 -2311 2349 -2290
rect 2412 -2311 2593 -2277
rect 2337 -2342 2349 -2311
rect 2401 -2342 2593 -2311
rect 1489 -2360 2593 -2342
rect 849 -2425 1285 -2387
rect 849 -2459 872 -2425
rect 906 -2459 1285 -2425
rect 849 -2497 1285 -2459
rect 849 -2531 872 -2497
rect 906 -2531 1285 -2497
rect 849 -2569 1285 -2531
rect 849 -2603 872 -2569
rect 906 -2603 1285 -2569
rect 849 -2640 1285 -2603
rect 849 -2641 1080 -2640
rect 849 -2675 872 -2641
rect 906 -2674 1080 -2641
rect 1114 -2674 1152 -2640
rect 1186 -2674 1285 -2640
rect 906 -2675 1285 -2674
rect 849 -2713 1285 -2675
rect 1489 -2428 2455 -2410
rect 1489 -2480 1539 -2428
rect 1591 -2480 1603 -2428
rect 1655 -2480 1667 -2428
rect 1719 -2480 1735 -2428
rect 1787 -2480 1799 -2428
rect 1851 -2480 1863 -2428
rect 1915 -2480 2025 -2428
rect 2077 -2480 2089 -2428
rect 2141 -2480 2153 -2428
rect 2205 -2480 2221 -2428
rect 2273 -2480 2285 -2428
rect 2337 -2480 2349 -2428
rect 2401 -2480 2455 -2428
rect 1489 -2606 2455 -2480
rect 1489 -2640 1539 -2606
rect 1489 -2674 1532 -2640
rect 1591 -2658 1603 -2606
rect 1655 -2658 1667 -2606
rect 1719 -2658 1735 -2606
rect 1787 -2640 1799 -2606
rect 1851 -2640 1863 -2606
rect 1787 -2658 1790 -2640
rect 1851 -2658 1862 -2640
rect 1915 -2658 2025 -2606
rect 2077 -2640 2089 -2606
rect 2141 -2640 2153 -2606
rect 2082 -2658 2089 -2640
rect 2205 -2658 2221 -2606
rect 2273 -2658 2285 -2606
rect 2337 -2640 2349 -2606
rect 2401 -2640 2455 -2606
rect 2340 -2658 2349 -2640
rect 1566 -2674 1604 -2658
rect 1638 -2674 1790 -2658
rect 1824 -2674 1862 -2658
rect 1896 -2674 2048 -2658
rect 2082 -2674 2120 -2658
rect 2154 -2674 2306 -2658
rect 2340 -2674 2378 -2658
rect 2412 -2674 2455 -2640
rect 1489 -2680 2455 -2674
rect 2532 -2592 2593 -2360
rect 2715 -2277 3423 -2271
rect 2715 -2311 2758 -2277
rect 2792 -2311 2830 -2277
rect 2864 -2311 3016 -2277
rect 3050 -2311 3088 -2277
rect 3122 -2311 3274 -2277
rect 3308 -2311 3346 -2277
rect 3380 -2311 3423 -2277
rect 2715 -2428 3423 -2311
rect 2715 -2480 2749 -2428
rect 2801 -2480 2813 -2428
rect 2865 -2480 2877 -2428
rect 2929 -2480 2945 -2428
rect 2997 -2480 3009 -2428
rect 3061 -2480 3073 -2428
rect 3125 -2480 3137 -2428
rect 3189 -2480 3205 -2428
rect 3257 -2480 3269 -2428
rect 3321 -2480 3333 -2428
rect 3385 -2480 3423 -2428
rect 2715 -2498 3423 -2480
rect 3545 -2277 4649 -2271
rect 3545 -2311 3726 -2277
rect 3760 -2290 3798 -2277
rect 3832 -2290 3984 -2277
rect 4018 -2290 4056 -2277
rect 4090 -2290 4242 -2277
rect 4276 -2290 4314 -2277
rect 4348 -2290 4500 -2277
rect 4534 -2290 4572 -2277
rect 3789 -2311 3798 -2290
rect 3545 -2342 3737 -2311
rect 3789 -2342 3801 -2311
rect 3853 -2342 3865 -2290
rect 3917 -2342 3933 -2290
rect 4049 -2311 4056 -2290
rect 3985 -2342 3997 -2311
rect 4049 -2342 4061 -2311
rect 4113 -2342 4223 -2290
rect 4276 -2311 4287 -2290
rect 4348 -2311 4351 -2290
rect 4275 -2342 4287 -2311
rect 4339 -2342 4351 -2311
rect 4403 -2342 4419 -2290
rect 4471 -2342 4483 -2290
rect 4535 -2342 4547 -2290
rect 4606 -2311 4649 -2277
rect 4599 -2342 4649 -2311
rect 3545 -2360 4649 -2342
rect 4853 -2277 5643 -2243
rect 9210 -2243 9589 -2209
rect 9623 -2243 9646 -2209
rect 4853 -2311 4952 -2277
rect 4986 -2311 5024 -2277
rect 5058 -2281 5438 -2277
rect 5058 -2311 5231 -2281
rect 4853 -2315 5231 -2311
rect 5265 -2311 5438 -2281
rect 5472 -2311 5510 -2277
rect 5544 -2311 5643 -2277
rect 5265 -2315 5643 -2311
rect 4853 -2353 5643 -2315
rect 3545 -2592 3606 -2360
rect 4853 -2387 5231 -2353
rect 5265 -2387 5643 -2353
rect 5846 -2277 6950 -2271
rect 5846 -2311 5889 -2277
rect 5923 -2290 5961 -2277
rect 5995 -2290 6147 -2277
rect 6181 -2290 6219 -2277
rect 6253 -2290 6405 -2277
rect 6439 -2290 6477 -2277
rect 6511 -2290 6663 -2277
rect 6697 -2290 6735 -2277
rect 5846 -2342 5896 -2311
rect 5948 -2342 5960 -2290
rect 6012 -2342 6024 -2290
rect 6076 -2342 6092 -2290
rect 6144 -2311 6147 -2290
rect 6208 -2311 6219 -2290
rect 6144 -2342 6156 -2311
rect 6208 -2342 6220 -2311
rect 6272 -2342 6382 -2290
rect 6439 -2311 6446 -2290
rect 6434 -2342 6446 -2311
rect 6498 -2342 6510 -2311
rect 6562 -2342 6578 -2290
rect 6630 -2342 6642 -2290
rect 6697 -2311 6706 -2290
rect 6769 -2311 6950 -2277
rect 6694 -2342 6706 -2311
rect 6758 -2342 6950 -2311
rect 5846 -2360 6950 -2342
rect 2532 -2640 3606 -2592
rect 2532 -2674 2758 -2640
rect 2792 -2674 2830 -2640
rect 2864 -2674 3016 -2640
rect 3050 -2674 3088 -2640
rect 3122 -2674 3274 -2640
rect 3308 -2674 3346 -2640
rect 3380 -2674 3606 -2640
rect 2532 -2680 3606 -2674
rect 3683 -2428 4649 -2410
rect 3683 -2480 3737 -2428
rect 3789 -2480 3801 -2428
rect 3853 -2480 3865 -2428
rect 3917 -2480 3933 -2428
rect 3985 -2480 3997 -2428
rect 4049 -2480 4061 -2428
rect 4113 -2480 4223 -2428
rect 4275 -2480 4287 -2428
rect 4339 -2480 4351 -2428
rect 4403 -2480 4419 -2428
rect 4471 -2480 4483 -2428
rect 4535 -2480 4547 -2428
rect 4599 -2480 4649 -2428
rect 3683 -2606 4649 -2480
rect 3683 -2640 3737 -2606
rect 3789 -2640 3801 -2606
rect 3683 -2674 3726 -2640
rect 3789 -2658 3798 -2640
rect 3853 -2658 3865 -2606
rect 3917 -2658 3933 -2606
rect 3985 -2640 3997 -2606
rect 4049 -2640 4061 -2606
rect 4049 -2658 4056 -2640
rect 4113 -2658 4223 -2606
rect 4275 -2640 4287 -2606
rect 4339 -2640 4351 -2606
rect 4276 -2658 4287 -2640
rect 4348 -2658 4351 -2640
rect 4403 -2658 4419 -2606
rect 4471 -2658 4483 -2606
rect 4535 -2658 4547 -2606
rect 4599 -2640 4649 -2606
rect 3760 -2674 3798 -2658
rect 3832 -2674 3984 -2658
rect 4018 -2674 4056 -2658
rect 4090 -2674 4242 -2658
rect 4276 -2674 4314 -2658
rect 4348 -2674 4500 -2658
rect 4534 -2674 4572 -2658
rect 4606 -2674 4649 -2640
rect 3683 -2680 4649 -2674
rect 4853 -2425 5643 -2387
rect 4853 -2459 5231 -2425
rect 5265 -2459 5643 -2425
rect 4853 -2497 5643 -2459
rect 4853 -2531 5231 -2497
rect 5265 -2531 5643 -2497
rect 4853 -2569 5643 -2531
rect 4853 -2603 5231 -2569
rect 5265 -2603 5643 -2569
rect 4853 -2640 5643 -2603
rect 4853 -2674 4952 -2640
rect 4986 -2674 5024 -2640
rect 5058 -2641 5438 -2640
rect 5058 -2674 5231 -2641
rect 4853 -2675 5231 -2674
rect 5265 -2674 5438 -2641
rect 5472 -2674 5510 -2640
rect 5544 -2674 5643 -2640
rect 5265 -2675 5643 -2674
rect 849 -2747 872 -2713
rect 906 -2747 1285 -2713
rect 4853 -2713 5643 -2675
rect 5846 -2428 6812 -2410
rect 5846 -2480 5896 -2428
rect 5948 -2480 5960 -2428
rect 6012 -2480 6024 -2428
rect 6076 -2480 6092 -2428
rect 6144 -2480 6156 -2428
rect 6208 -2480 6220 -2428
rect 6272 -2480 6382 -2428
rect 6434 -2480 6446 -2428
rect 6498 -2480 6510 -2428
rect 6562 -2480 6578 -2428
rect 6630 -2480 6642 -2428
rect 6694 -2480 6706 -2428
rect 6758 -2480 6812 -2428
rect 5846 -2606 6812 -2480
rect 5846 -2640 5896 -2606
rect 5846 -2674 5889 -2640
rect 5948 -2658 5960 -2606
rect 6012 -2658 6024 -2606
rect 6076 -2658 6092 -2606
rect 6144 -2640 6156 -2606
rect 6208 -2640 6220 -2606
rect 6144 -2658 6147 -2640
rect 6208 -2658 6219 -2640
rect 6272 -2658 6382 -2606
rect 6434 -2640 6446 -2606
rect 6498 -2640 6510 -2606
rect 6439 -2658 6446 -2640
rect 6562 -2658 6578 -2606
rect 6630 -2658 6642 -2606
rect 6694 -2640 6706 -2606
rect 6758 -2640 6812 -2606
rect 6697 -2658 6706 -2640
rect 5923 -2674 5961 -2658
rect 5995 -2674 6147 -2658
rect 6181 -2674 6219 -2658
rect 6253 -2674 6405 -2658
rect 6439 -2674 6477 -2658
rect 6511 -2674 6663 -2658
rect 6697 -2674 6735 -2658
rect 6769 -2674 6812 -2640
rect 5846 -2680 6812 -2674
rect 6889 -2592 6950 -2360
rect 7072 -2277 7780 -2271
rect 7072 -2311 7115 -2277
rect 7149 -2311 7187 -2277
rect 7221 -2311 7373 -2277
rect 7407 -2311 7445 -2277
rect 7479 -2311 7631 -2277
rect 7665 -2311 7703 -2277
rect 7737 -2311 7780 -2277
rect 7072 -2428 7780 -2311
rect 7072 -2480 7110 -2428
rect 7162 -2480 7174 -2428
rect 7226 -2480 7238 -2428
rect 7290 -2480 7306 -2428
rect 7358 -2480 7370 -2428
rect 7422 -2480 7434 -2428
rect 7486 -2480 7498 -2428
rect 7550 -2480 7566 -2428
rect 7618 -2480 7630 -2428
rect 7682 -2480 7694 -2428
rect 7746 -2480 7780 -2428
rect 7072 -2498 7780 -2480
rect 7902 -2277 9006 -2271
rect 7902 -2311 8083 -2277
rect 8117 -2290 8155 -2277
rect 8189 -2290 8341 -2277
rect 8375 -2290 8413 -2277
rect 8447 -2290 8599 -2277
rect 8633 -2290 8671 -2277
rect 8705 -2290 8857 -2277
rect 8891 -2290 8929 -2277
rect 8146 -2311 8155 -2290
rect 7902 -2342 8094 -2311
rect 8146 -2342 8158 -2311
rect 8210 -2342 8222 -2290
rect 8274 -2342 8290 -2290
rect 8406 -2311 8413 -2290
rect 8342 -2342 8354 -2311
rect 8406 -2342 8418 -2311
rect 8470 -2342 8580 -2290
rect 8633 -2311 8644 -2290
rect 8705 -2311 8708 -2290
rect 8632 -2342 8644 -2311
rect 8696 -2342 8708 -2311
rect 8760 -2342 8776 -2290
rect 8828 -2342 8840 -2290
rect 8892 -2342 8904 -2290
rect 8963 -2311 9006 -2277
rect 8956 -2342 9006 -2311
rect 7902 -2360 9006 -2342
rect 9210 -2277 9646 -2243
rect 9210 -2311 9309 -2277
rect 9343 -2311 9381 -2277
rect 9415 -2281 9646 -2277
rect 9415 -2311 9589 -2281
rect 9210 -2315 9589 -2311
rect 9623 -2315 9646 -2281
rect 9210 -2353 9646 -2315
rect 7902 -2592 7963 -2360
rect 9210 -2387 9589 -2353
rect 9623 -2387 9646 -2353
rect 6889 -2640 7963 -2592
rect 6889 -2674 7115 -2640
rect 7149 -2674 7187 -2640
rect 7221 -2674 7373 -2640
rect 7407 -2674 7445 -2640
rect 7479 -2674 7631 -2640
rect 7665 -2674 7703 -2640
rect 7737 -2674 7963 -2640
rect 6889 -2680 7963 -2674
rect 8040 -2428 9006 -2410
rect 8040 -2480 8094 -2428
rect 8146 -2480 8158 -2428
rect 8210 -2480 8222 -2428
rect 8274 -2480 8290 -2428
rect 8342 -2480 8354 -2428
rect 8406 -2480 8418 -2428
rect 8470 -2480 8580 -2428
rect 8632 -2480 8644 -2428
rect 8696 -2480 8708 -2428
rect 8760 -2480 8776 -2428
rect 8828 -2480 8840 -2428
rect 8892 -2480 8904 -2428
rect 8956 -2480 9006 -2428
rect 8040 -2606 9006 -2480
rect 8040 -2640 8094 -2606
rect 8146 -2640 8158 -2606
rect 8040 -2674 8083 -2640
rect 8146 -2658 8155 -2640
rect 8210 -2658 8222 -2606
rect 8274 -2658 8290 -2606
rect 8342 -2640 8354 -2606
rect 8406 -2640 8418 -2606
rect 8406 -2658 8413 -2640
rect 8470 -2658 8580 -2606
rect 8632 -2640 8644 -2606
rect 8696 -2640 8708 -2606
rect 8633 -2658 8644 -2640
rect 8705 -2658 8708 -2640
rect 8760 -2658 8776 -2606
rect 8828 -2658 8840 -2606
rect 8892 -2658 8904 -2606
rect 8956 -2640 9006 -2606
rect 8117 -2674 8155 -2658
rect 8189 -2674 8341 -2658
rect 8375 -2674 8413 -2658
rect 8447 -2674 8599 -2658
rect 8633 -2674 8671 -2658
rect 8705 -2674 8857 -2658
rect 8891 -2674 8929 -2658
rect 8963 -2674 9006 -2640
rect 8040 -2680 9006 -2674
rect 9210 -2425 9646 -2387
rect 9210 -2459 9589 -2425
rect 9623 -2459 9646 -2425
rect 9210 -2497 9646 -2459
rect 9210 -2531 9589 -2497
rect 9623 -2531 9646 -2497
rect 9210 -2569 9646 -2531
rect 9210 -2603 9589 -2569
rect 9623 -2603 9646 -2569
rect 9210 -2640 9646 -2603
rect 9210 -2674 9309 -2640
rect 9343 -2674 9381 -2640
rect 9415 -2641 9646 -2640
rect 9415 -2674 9589 -2641
rect 9210 -2675 9589 -2674
rect 9623 -2675 9646 -2641
rect 849 -2768 1285 -2747
rect 849 -2785 987 -2768
rect 849 -2819 872 -2785
rect 906 -2802 987 -2785
rect 1021 -2802 1245 -2768
rect 1279 -2802 1285 -2768
rect 906 -2819 1285 -2802
rect 849 -2840 1285 -2819
rect 849 -2857 987 -2840
rect 849 -2891 872 -2857
rect 906 -2874 987 -2857
rect 1021 -2874 1245 -2840
rect 1279 -2874 1285 -2840
rect 906 -2891 1285 -2874
rect 849 -2929 1285 -2891
rect 849 -2963 872 -2929
rect 906 -2963 1285 -2929
rect 849 -3001 1285 -2963
rect 849 -3035 872 -3001
rect 906 -3035 1285 -3001
rect 849 -3073 1285 -3035
rect 849 -3107 872 -3073
rect 906 -3107 1285 -3073
rect 849 -3145 1285 -3107
rect 849 -3179 872 -3145
rect 906 -3179 1285 -3145
rect 849 -3217 1285 -3179
rect 849 -3251 872 -3217
rect 906 -3251 1285 -3217
rect 849 -3289 1285 -3251
rect 849 -3323 872 -3289
rect 906 -3323 1285 -3289
rect 849 -3361 1285 -3323
rect 1433 -2768 1479 -2721
rect 1433 -2802 1439 -2768
rect 1473 -2802 1479 -2768
rect 1433 -2840 1479 -2802
rect 1433 -2874 1439 -2840
rect 1473 -2874 1479 -2840
rect 1433 -3354 1479 -2874
rect 1691 -2768 1737 -2721
rect 1691 -2802 1697 -2768
rect 1731 -2802 1737 -2768
rect 1691 -2840 1737 -2802
rect 1691 -2874 1697 -2840
rect 1731 -2874 1737 -2840
rect 1691 -3023 1737 -2874
rect 1949 -2768 1995 -2721
rect 1949 -2802 1955 -2768
rect 1989 -2802 1995 -2768
rect 1949 -2840 1995 -2802
rect 1949 -2874 1955 -2840
rect 1989 -2874 1995 -2840
rect 1615 -3033 1811 -3023
rect 1615 -3085 1624 -3033
rect 1676 -3085 1688 -3033
rect 1740 -3085 1752 -3033
rect 1804 -3085 1811 -3033
rect 1615 -3093 1811 -3085
rect 1949 -3354 1995 -2874
rect 2207 -2768 2253 -2721
rect 2207 -2802 2213 -2768
rect 2247 -2802 2253 -2768
rect 2207 -2840 2253 -2802
rect 2207 -2874 2213 -2840
rect 2247 -2874 2253 -2840
rect 2207 -3023 2253 -2874
rect 2465 -2768 2511 -2721
rect 2465 -2802 2471 -2768
rect 2505 -2802 2511 -2768
rect 2465 -2840 2511 -2802
rect 2465 -2874 2471 -2840
rect 2505 -2874 2511 -2840
rect 2132 -3033 2328 -3023
rect 2132 -3085 2141 -3033
rect 2193 -3085 2205 -3033
rect 2257 -3085 2269 -3033
rect 2321 -3085 2328 -3033
rect 2132 -3093 2328 -3085
rect 2465 -3354 2511 -2874
rect 2659 -2768 2705 -2721
rect 2659 -2802 2665 -2768
rect 2699 -2802 2705 -2768
rect 2659 -2840 2705 -2802
rect 2659 -2874 2665 -2840
rect 2699 -2874 2705 -2840
rect 2659 -3192 2705 -2874
rect 2917 -2768 2963 -2721
rect 2917 -2802 2923 -2768
rect 2957 -2802 2963 -2768
rect 2917 -2840 2963 -2802
rect 2917 -2874 2923 -2840
rect 2957 -2874 2963 -2840
rect 2586 -3202 2782 -3192
rect 2586 -3254 2593 -3202
rect 2645 -3254 2657 -3202
rect 2709 -3254 2721 -3202
rect 2773 -3254 2782 -3202
rect 2586 -3262 2782 -3254
rect 849 -3395 872 -3361
rect 906 -3395 1285 -3361
rect 849 -3433 1285 -3395
rect 1355 -3364 1551 -3354
rect 1355 -3416 1364 -3364
rect 1416 -3416 1428 -3364
rect 1480 -3416 1492 -3364
rect 1544 -3416 1551 -3364
rect 1355 -3424 1551 -3416
rect 1873 -3364 2069 -3354
rect 1873 -3416 1882 -3364
rect 1934 -3416 1946 -3364
rect 1998 -3416 2010 -3364
rect 2062 -3416 2069 -3364
rect 1873 -3424 2069 -3416
rect 2389 -3364 2585 -3354
rect 2389 -3416 2398 -3364
rect 2450 -3416 2462 -3364
rect 2514 -3416 2526 -3364
rect 2578 -3416 2585 -3364
rect 2389 -3424 2585 -3416
rect 849 -3467 872 -3433
rect 906 -3467 1285 -3433
rect 849 -3505 1285 -3467
rect 849 -3539 872 -3505
rect 906 -3539 1285 -3505
rect 2917 -3523 2963 -2874
rect 3175 -2768 3221 -2721
rect 3175 -2802 3181 -2768
rect 3215 -2802 3221 -2768
rect 3175 -2840 3221 -2802
rect 3175 -2874 3181 -2840
rect 3215 -2874 3221 -2840
rect 3175 -3192 3221 -2874
rect 3433 -2768 3479 -2721
rect 3433 -2802 3439 -2768
rect 3473 -2802 3479 -2768
rect 3433 -2840 3479 -2802
rect 3433 -2874 3439 -2840
rect 3473 -2874 3479 -2840
rect 3103 -3202 3299 -3192
rect 3103 -3254 3110 -3202
rect 3162 -3254 3174 -3202
rect 3226 -3254 3238 -3202
rect 3290 -3254 3299 -3202
rect 3103 -3262 3299 -3254
rect 3433 -3523 3479 -2874
rect 3627 -2768 3673 -2721
rect 3627 -2802 3633 -2768
rect 3667 -2802 3673 -2768
rect 3627 -2840 3673 -2802
rect 3627 -2874 3633 -2840
rect 3667 -2874 3673 -2840
rect 3627 -3354 3673 -2874
rect 3885 -2768 3931 -2721
rect 3885 -2802 3891 -2768
rect 3925 -2802 3931 -2768
rect 3885 -2840 3931 -2802
rect 3885 -2874 3891 -2840
rect 3925 -2874 3931 -2840
rect 3885 -3023 3931 -2874
rect 4143 -2768 4189 -2721
rect 4143 -2802 4149 -2768
rect 4183 -2802 4189 -2768
rect 4143 -2840 4189 -2802
rect 4143 -2874 4149 -2840
rect 4183 -2874 4189 -2840
rect 3809 -3033 4005 -3023
rect 3809 -3085 3818 -3033
rect 3870 -3085 3882 -3033
rect 3934 -3085 3946 -3033
rect 3998 -3085 4005 -3033
rect 3809 -3093 4005 -3085
rect 4143 -3354 4189 -2874
rect 4401 -2768 4447 -2721
rect 4401 -2802 4407 -2768
rect 4441 -2802 4447 -2768
rect 4401 -2840 4447 -2802
rect 4401 -2874 4407 -2840
rect 4441 -2874 4447 -2840
rect 4401 -3023 4447 -2874
rect 4659 -2768 4705 -2721
rect 4659 -2802 4665 -2768
rect 4699 -2802 4705 -2768
rect 4659 -2840 4705 -2802
rect 4659 -2874 4665 -2840
rect 4699 -2874 4705 -2840
rect 4326 -3033 4522 -3023
rect 4326 -3085 4335 -3033
rect 4387 -3085 4399 -3033
rect 4451 -3085 4463 -3033
rect 4515 -3085 4522 -3033
rect 4326 -3093 4522 -3085
rect 4659 -3354 4705 -2874
rect 4853 -2747 5231 -2713
rect 5265 -2747 5643 -2713
rect 9210 -2713 9646 -2675
rect 4853 -2768 5643 -2747
rect 4853 -2802 4859 -2768
rect 4893 -2802 5117 -2768
rect 5151 -2785 5345 -2768
rect 5151 -2802 5231 -2785
rect 4853 -2819 5231 -2802
rect 5265 -2802 5345 -2785
rect 5379 -2802 5603 -2768
rect 5637 -2802 5643 -2768
rect 5265 -2819 5643 -2802
rect 4853 -2840 5643 -2819
rect 4853 -2874 4859 -2840
rect 4893 -2874 5117 -2840
rect 5151 -2857 5345 -2840
rect 5151 -2874 5231 -2857
rect 4853 -2891 5231 -2874
rect 5265 -2874 5345 -2857
rect 5379 -2874 5603 -2840
rect 5637 -2874 5643 -2840
rect 5265 -2891 5643 -2874
rect 4853 -2929 5643 -2891
rect 4853 -2963 5231 -2929
rect 5265 -2963 5643 -2929
rect 4853 -3001 5643 -2963
rect 4853 -3035 5231 -3001
rect 5265 -3035 5643 -3001
rect 4853 -3073 5643 -3035
rect 4853 -3107 5231 -3073
rect 5265 -3107 5643 -3073
rect 4853 -3145 5643 -3107
rect 4853 -3179 5231 -3145
rect 5265 -3179 5643 -3145
rect 4853 -3217 5643 -3179
rect 4853 -3251 5231 -3217
rect 5265 -3251 5643 -3217
rect 4853 -3289 5643 -3251
rect 4853 -3323 5231 -3289
rect 5265 -3323 5643 -3289
rect 3550 -3364 3746 -3354
rect 3550 -3416 3559 -3364
rect 3611 -3416 3623 -3364
rect 3675 -3416 3687 -3364
rect 3739 -3416 3746 -3364
rect 3550 -3424 3746 -3416
rect 4067 -3364 4263 -3354
rect 4067 -3416 4076 -3364
rect 4128 -3416 4140 -3364
rect 4192 -3416 4204 -3364
rect 4256 -3416 4263 -3364
rect 4067 -3424 4263 -3416
rect 4582 -3364 4778 -3354
rect 4582 -3416 4591 -3364
rect 4643 -3416 4655 -3364
rect 4707 -3416 4719 -3364
rect 4771 -3416 4778 -3364
rect 4582 -3424 4778 -3416
rect 4853 -3361 5643 -3323
rect 5790 -2768 5836 -2721
rect 5790 -2802 5796 -2768
rect 5830 -2802 5836 -2768
rect 5790 -2840 5836 -2802
rect 5790 -2874 5796 -2840
rect 5830 -2874 5836 -2840
rect 5790 -3354 5836 -2874
rect 6048 -2768 6094 -2721
rect 6048 -2802 6054 -2768
rect 6088 -2802 6094 -2768
rect 6048 -2840 6094 -2802
rect 6048 -2874 6054 -2840
rect 6088 -2874 6094 -2840
rect 6048 -3023 6094 -2874
rect 6306 -2768 6352 -2721
rect 6306 -2802 6312 -2768
rect 6346 -2802 6352 -2768
rect 6306 -2840 6352 -2802
rect 6306 -2874 6312 -2840
rect 6346 -2874 6352 -2840
rect 5973 -3033 6169 -3023
rect 5973 -3085 5980 -3033
rect 6032 -3085 6044 -3033
rect 6096 -3085 6108 -3033
rect 6160 -3085 6169 -3033
rect 5973 -3093 6169 -3085
rect 6306 -3354 6352 -2874
rect 6564 -2768 6610 -2721
rect 6564 -2802 6570 -2768
rect 6604 -2802 6610 -2768
rect 6564 -2840 6610 -2802
rect 6564 -2874 6570 -2840
rect 6604 -2874 6610 -2840
rect 6564 -3023 6610 -2874
rect 6822 -2768 6868 -2721
rect 6822 -2802 6828 -2768
rect 6862 -2802 6868 -2768
rect 6822 -2840 6868 -2802
rect 6822 -2874 6828 -2840
rect 6862 -2874 6868 -2840
rect 6490 -3033 6686 -3023
rect 6490 -3085 6497 -3033
rect 6549 -3085 6561 -3033
rect 6613 -3085 6625 -3033
rect 6677 -3085 6686 -3033
rect 6490 -3093 6686 -3085
rect 6822 -3354 6868 -2874
rect 7016 -2768 7062 -2721
rect 7016 -2802 7022 -2768
rect 7056 -2802 7062 -2768
rect 7016 -2840 7062 -2802
rect 7016 -2874 7022 -2840
rect 7056 -2874 7062 -2840
rect 4853 -3395 5231 -3361
rect 5265 -3395 5643 -3361
rect 4853 -3433 5643 -3395
rect 5717 -3364 5913 -3354
rect 5717 -3416 5724 -3364
rect 5776 -3416 5788 -3364
rect 5840 -3416 5852 -3364
rect 5904 -3416 5913 -3364
rect 5717 -3424 5913 -3416
rect 6232 -3364 6428 -3354
rect 6232 -3416 6239 -3364
rect 6291 -3416 6303 -3364
rect 6355 -3416 6367 -3364
rect 6419 -3416 6428 -3364
rect 6232 -3424 6428 -3416
rect 6749 -3364 6945 -3354
rect 6749 -3416 6756 -3364
rect 6808 -3416 6820 -3364
rect 6872 -3416 6884 -3364
rect 6936 -3416 6945 -3364
rect 6749 -3424 6945 -3416
rect 4853 -3467 5231 -3433
rect 5265 -3467 5643 -3433
rect 4853 -3505 5643 -3467
rect 849 -3577 1285 -3539
rect 849 -3611 872 -3577
rect 906 -3611 1285 -3577
rect 2843 -3533 3039 -3523
rect 2843 -3585 2850 -3533
rect 2902 -3585 2914 -3533
rect 2966 -3585 2978 -3533
rect 3030 -3585 3039 -3533
rect 2843 -3593 3039 -3585
rect 3361 -3533 3557 -3523
rect 3361 -3585 3368 -3533
rect 3420 -3585 3432 -3533
rect 3484 -3585 3496 -3533
rect 3548 -3585 3557 -3533
rect 3361 -3593 3557 -3585
rect 4853 -3539 5231 -3505
rect 5265 -3539 5643 -3505
rect 7016 -3523 7062 -2874
rect 7274 -2768 7320 -2721
rect 7274 -2802 7280 -2768
rect 7314 -2802 7320 -2768
rect 7274 -2840 7320 -2802
rect 7274 -2874 7280 -2840
rect 7314 -2874 7320 -2840
rect 7274 -3192 7320 -2874
rect 7532 -2768 7578 -2721
rect 7532 -2802 7538 -2768
rect 7572 -2802 7578 -2768
rect 7532 -2840 7578 -2802
rect 7532 -2874 7538 -2840
rect 7572 -2874 7578 -2840
rect 7196 -3202 7392 -3192
rect 7196 -3254 7205 -3202
rect 7257 -3254 7269 -3202
rect 7321 -3254 7333 -3202
rect 7385 -3254 7392 -3202
rect 7196 -3262 7392 -3254
rect 7532 -3523 7578 -2874
rect 7790 -2768 7836 -2721
rect 7790 -2802 7796 -2768
rect 7830 -2802 7836 -2768
rect 7790 -2840 7836 -2802
rect 7790 -2874 7796 -2840
rect 7830 -2874 7836 -2840
rect 7790 -3192 7836 -2874
rect 7984 -2768 8030 -2721
rect 7984 -2802 7990 -2768
rect 8024 -2802 8030 -2768
rect 7984 -2840 8030 -2802
rect 7984 -2874 7990 -2840
rect 8024 -2874 8030 -2840
rect 7713 -3202 7909 -3192
rect 7713 -3254 7722 -3202
rect 7774 -3254 7786 -3202
rect 7838 -3254 7850 -3202
rect 7902 -3254 7909 -3202
rect 7713 -3262 7909 -3254
rect 7984 -3354 8030 -2874
rect 8242 -2768 8288 -2721
rect 8242 -2802 8248 -2768
rect 8282 -2802 8288 -2768
rect 8242 -2840 8288 -2802
rect 8242 -2874 8248 -2840
rect 8282 -2874 8288 -2840
rect 8242 -3023 8288 -2874
rect 8500 -2768 8546 -2721
rect 8500 -2802 8506 -2768
rect 8540 -2802 8546 -2768
rect 8500 -2840 8546 -2802
rect 8500 -2874 8506 -2840
rect 8540 -2874 8546 -2840
rect 8167 -3033 8363 -3023
rect 8167 -3085 8174 -3033
rect 8226 -3085 8238 -3033
rect 8290 -3085 8302 -3033
rect 8354 -3085 8363 -3033
rect 8167 -3093 8363 -3085
rect 8500 -3354 8546 -2874
rect 8758 -2768 8804 -2721
rect 8758 -2802 8764 -2768
rect 8798 -2802 8804 -2768
rect 8758 -2840 8804 -2802
rect 8758 -2874 8764 -2840
rect 8798 -2874 8804 -2840
rect 8758 -3023 8804 -2874
rect 9016 -2768 9062 -2721
rect 9016 -2802 9022 -2768
rect 9056 -2802 9062 -2768
rect 9016 -2840 9062 -2802
rect 9016 -2874 9022 -2840
rect 9056 -2874 9062 -2840
rect 8685 -3033 8881 -3023
rect 8685 -3085 8692 -3033
rect 8744 -3085 8756 -3033
rect 8808 -3085 8820 -3033
rect 8872 -3085 8881 -3033
rect 8685 -3093 8881 -3085
rect 9016 -3354 9062 -2874
rect 9210 -2747 9589 -2713
rect 9623 -2747 9646 -2713
rect 9210 -2768 9646 -2747
rect 9210 -2802 9216 -2768
rect 9250 -2802 9474 -2768
rect 9508 -2785 9646 -2768
rect 9508 -2802 9589 -2785
rect 9210 -2819 9589 -2802
rect 9623 -2819 9646 -2785
rect 9210 -2840 9646 -2819
rect 9210 -2874 9216 -2840
rect 9250 -2874 9474 -2840
rect 9508 -2857 9646 -2840
rect 9508 -2874 9589 -2857
rect 9210 -2891 9589 -2874
rect 9623 -2891 9646 -2857
rect 9210 -2929 9646 -2891
rect 9210 -2963 9589 -2929
rect 9623 -2963 9646 -2929
rect 9210 -3001 9646 -2963
rect 9210 -3035 9589 -3001
rect 9623 -3035 9646 -3001
rect 9210 -3073 9646 -3035
rect 9210 -3107 9589 -3073
rect 9623 -3107 9646 -3073
rect 9210 -3145 9646 -3107
rect 9210 -3179 9589 -3145
rect 9623 -3179 9646 -3145
rect 9210 -3217 9646 -3179
rect 9210 -3251 9589 -3217
rect 9623 -3251 9646 -3217
rect 9210 -3289 9646 -3251
rect 9210 -3323 9589 -3289
rect 9623 -3323 9646 -3289
rect 7910 -3364 8106 -3354
rect 7910 -3416 7917 -3364
rect 7969 -3416 7981 -3364
rect 8033 -3416 8045 -3364
rect 8097 -3416 8106 -3364
rect 7910 -3424 8106 -3416
rect 8427 -3364 8623 -3354
rect 8427 -3416 8434 -3364
rect 8486 -3416 8498 -3364
rect 8550 -3416 8562 -3364
rect 8614 -3416 8623 -3364
rect 8427 -3424 8623 -3416
rect 8944 -3364 9140 -3354
rect 8944 -3416 8951 -3364
rect 9003 -3416 9015 -3364
rect 9067 -3416 9079 -3364
rect 9131 -3416 9140 -3364
rect 8944 -3424 9140 -3416
rect 9210 -3361 9646 -3323
rect 9210 -3395 9589 -3361
rect 9623 -3395 9646 -3361
rect 9210 -3433 9646 -3395
rect 9210 -3467 9589 -3433
rect 9623 -3467 9646 -3433
rect 9210 -3505 9646 -3467
rect 4853 -3577 5643 -3539
rect 849 -3649 1285 -3611
rect 849 -3683 872 -3649
rect 906 -3683 1285 -3649
rect 849 -3721 1285 -3683
rect 4853 -3611 5231 -3577
rect 5265 -3611 5643 -3577
rect 6939 -3533 7135 -3523
rect 6939 -3585 6948 -3533
rect 7000 -3585 7012 -3533
rect 7064 -3585 7076 -3533
rect 7128 -3585 7135 -3533
rect 6939 -3593 7135 -3585
rect 7456 -3533 7652 -3523
rect 7456 -3585 7465 -3533
rect 7517 -3585 7529 -3533
rect 7581 -3585 7593 -3533
rect 7645 -3585 7652 -3533
rect 7456 -3593 7652 -3585
rect 9210 -3539 9589 -3505
rect 9623 -3539 9646 -3505
rect 9210 -3577 9646 -3539
rect 4853 -3649 5643 -3611
rect 4853 -3683 5231 -3649
rect 5265 -3683 5643 -3649
rect 849 -3755 872 -3721
rect 906 -3755 1285 -3721
rect 849 -3758 1285 -3755
rect 849 -3792 987 -3758
rect 1021 -3792 1245 -3758
rect 1279 -3792 1285 -3758
rect 849 -3793 1285 -3792
rect 849 -3827 872 -3793
rect 906 -3827 1285 -3793
rect 849 -3830 1285 -3827
rect 849 -3864 987 -3830
rect 1021 -3864 1245 -3830
rect 1279 -3864 1285 -3830
rect 849 -3865 1285 -3864
rect 849 -3899 872 -3865
rect 906 -3899 1285 -3865
rect 849 -3937 1285 -3899
rect 849 -3952 872 -3937
rect 847 -3971 872 -3952
rect 906 -3952 1285 -3937
rect 1433 -3758 1479 -3711
rect 1433 -3792 1439 -3758
rect 1473 -3792 1479 -3758
rect 1433 -3830 1479 -3792
rect 1433 -3864 1439 -3830
rect 1473 -3864 1479 -3830
rect 1433 -3952 1479 -3864
rect 1691 -3758 1737 -3711
rect 1691 -3792 1697 -3758
rect 1731 -3792 1737 -3758
rect 1691 -3830 1737 -3792
rect 1691 -3864 1697 -3830
rect 1731 -3864 1737 -3830
rect 1691 -3952 1737 -3864
rect 1949 -3758 1995 -3711
rect 1949 -3792 1955 -3758
rect 1989 -3792 1995 -3758
rect 1949 -3830 1995 -3792
rect 1949 -3864 1955 -3830
rect 1989 -3864 1995 -3830
rect 1949 -3952 1995 -3864
rect 2207 -3758 2253 -3711
rect 2207 -3792 2213 -3758
rect 2247 -3792 2253 -3758
rect 2207 -3830 2253 -3792
rect 2207 -3864 2213 -3830
rect 2247 -3864 2253 -3830
rect 2207 -3952 2253 -3864
rect 2465 -3758 2511 -3711
rect 2465 -3792 2471 -3758
rect 2505 -3792 2511 -3758
rect 2465 -3830 2511 -3792
rect 2465 -3864 2471 -3830
rect 2505 -3864 2511 -3830
rect 2465 -3952 2511 -3864
rect 2659 -3758 2705 -3711
rect 2659 -3792 2665 -3758
rect 2699 -3792 2705 -3758
rect 2659 -3830 2705 -3792
rect 2659 -3864 2665 -3830
rect 2699 -3864 2705 -3830
rect 2659 -3952 2705 -3864
rect 2917 -3758 2963 -3711
rect 2917 -3792 2923 -3758
rect 2957 -3792 2963 -3758
rect 2917 -3830 2963 -3792
rect 2917 -3864 2923 -3830
rect 2957 -3864 2963 -3830
rect 2917 -3952 2963 -3864
rect 3175 -3758 3221 -3711
rect 3175 -3792 3181 -3758
rect 3215 -3792 3221 -3758
rect 3175 -3830 3221 -3792
rect 3175 -3864 3181 -3830
rect 3215 -3864 3221 -3830
rect 3175 -3952 3221 -3864
rect 3433 -3758 3479 -3711
rect 3433 -3792 3439 -3758
rect 3473 -3792 3479 -3758
rect 3433 -3830 3479 -3792
rect 3433 -3864 3439 -3830
rect 3473 -3864 3479 -3830
rect 3433 -3952 3479 -3864
rect 3627 -3758 3673 -3711
rect 3627 -3792 3633 -3758
rect 3667 -3792 3673 -3758
rect 3627 -3830 3673 -3792
rect 3627 -3864 3633 -3830
rect 3667 -3864 3673 -3830
rect 3627 -3952 3673 -3864
rect 3885 -3758 3931 -3711
rect 3885 -3792 3891 -3758
rect 3925 -3792 3931 -3758
rect 3885 -3830 3931 -3792
rect 3885 -3864 3891 -3830
rect 3925 -3864 3931 -3830
rect 3885 -3952 3931 -3864
rect 4143 -3758 4189 -3711
rect 4143 -3792 4149 -3758
rect 4183 -3792 4189 -3758
rect 4143 -3830 4189 -3792
rect 4143 -3864 4149 -3830
rect 4183 -3864 4189 -3830
rect 4143 -3952 4189 -3864
rect 4401 -3758 4447 -3711
rect 4401 -3792 4407 -3758
rect 4441 -3792 4447 -3758
rect 4401 -3830 4447 -3792
rect 4401 -3864 4407 -3830
rect 4441 -3864 4447 -3830
rect 4401 -3952 4447 -3864
rect 4659 -3758 4705 -3711
rect 4659 -3792 4665 -3758
rect 4699 -3792 4705 -3758
rect 4659 -3830 4705 -3792
rect 4659 -3864 4665 -3830
rect 4699 -3864 4705 -3830
rect 4659 -3952 4705 -3864
rect 4853 -3721 5643 -3683
rect 9210 -3611 9589 -3577
rect 9623 -3611 9646 -3577
rect 9210 -3649 9646 -3611
rect 9210 -3683 9589 -3649
rect 9623 -3683 9646 -3649
rect 4853 -3755 5231 -3721
rect 5265 -3755 5643 -3721
rect 4853 -3758 5643 -3755
rect 4853 -3792 4859 -3758
rect 4893 -3792 5117 -3758
rect 5151 -3792 5345 -3758
rect 5379 -3792 5603 -3758
rect 5637 -3792 5643 -3758
rect 4853 -3793 5643 -3792
rect 4853 -3827 5231 -3793
rect 5265 -3827 5643 -3793
rect 4853 -3830 5643 -3827
rect 4853 -3864 4859 -3830
rect 4893 -3864 5117 -3830
rect 5151 -3864 5345 -3830
rect 5379 -3864 5603 -3830
rect 5637 -3864 5643 -3830
rect 4853 -3865 5643 -3864
rect 4853 -3899 5231 -3865
rect 5265 -3899 5643 -3865
rect 4853 -3937 5643 -3899
rect 4853 -3952 5231 -3937
rect 906 -3958 5231 -3952
rect 906 -3971 1080 -3958
rect 847 -3992 1080 -3971
rect 1114 -3992 1152 -3958
rect 1186 -3992 1532 -3958
rect 1566 -3992 1604 -3958
rect 1638 -3992 1790 -3958
rect 1824 -3992 1862 -3958
rect 1896 -3992 2048 -3958
rect 2082 -3992 2120 -3958
rect 2154 -3992 2306 -3958
rect 2340 -3992 2378 -3958
rect 2412 -3992 2758 -3958
rect 2792 -3992 2830 -3958
rect 2864 -3992 3016 -3958
rect 3050 -3992 3088 -3958
rect 3122 -3992 3274 -3958
rect 3308 -3992 3346 -3958
rect 3380 -3992 3726 -3958
rect 3760 -3992 3798 -3958
rect 3832 -3992 3984 -3958
rect 4018 -3992 4056 -3958
rect 4090 -3992 4242 -3958
rect 4276 -3992 4314 -3958
rect 4348 -3992 4500 -3958
rect 4534 -3992 4572 -3958
rect 4606 -3992 4952 -3958
rect 4986 -3992 5024 -3958
rect 5058 -3971 5231 -3958
rect 5265 -3952 5643 -3937
rect 5790 -3758 5836 -3711
rect 5790 -3792 5796 -3758
rect 5830 -3792 5836 -3758
rect 5790 -3830 5836 -3792
rect 5790 -3864 5796 -3830
rect 5830 -3864 5836 -3830
rect 5790 -3952 5836 -3864
rect 6048 -3758 6094 -3711
rect 6048 -3792 6054 -3758
rect 6088 -3792 6094 -3758
rect 6048 -3830 6094 -3792
rect 6048 -3864 6054 -3830
rect 6088 -3864 6094 -3830
rect 6048 -3952 6094 -3864
rect 6306 -3758 6352 -3711
rect 6306 -3792 6312 -3758
rect 6346 -3792 6352 -3758
rect 6306 -3830 6352 -3792
rect 6306 -3864 6312 -3830
rect 6346 -3864 6352 -3830
rect 6306 -3952 6352 -3864
rect 6564 -3758 6610 -3711
rect 6564 -3792 6570 -3758
rect 6604 -3792 6610 -3758
rect 6564 -3830 6610 -3792
rect 6564 -3864 6570 -3830
rect 6604 -3864 6610 -3830
rect 6564 -3952 6610 -3864
rect 6822 -3758 6868 -3711
rect 6822 -3792 6828 -3758
rect 6862 -3792 6868 -3758
rect 6822 -3830 6868 -3792
rect 6822 -3864 6828 -3830
rect 6862 -3864 6868 -3830
rect 6822 -3952 6868 -3864
rect 7016 -3758 7062 -3711
rect 7016 -3792 7022 -3758
rect 7056 -3792 7062 -3758
rect 7016 -3830 7062 -3792
rect 7016 -3864 7022 -3830
rect 7056 -3864 7062 -3830
rect 7016 -3952 7062 -3864
rect 7274 -3758 7320 -3711
rect 7274 -3792 7280 -3758
rect 7314 -3792 7320 -3758
rect 7274 -3830 7320 -3792
rect 7274 -3864 7280 -3830
rect 7314 -3864 7320 -3830
rect 7274 -3952 7320 -3864
rect 7532 -3758 7578 -3711
rect 7532 -3792 7538 -3758
rect 7572 -3792 7578 -3758
rect 7532 -3830 7578 -3792
rect 7532 -3864 7538 -3830
rect 7572 -3864 7578 -3830
rect 7532 -3952 7578 -3864
rect 7790 -3758 7836 -3711
rect 7790 -3792 7796 -3758
rect 7830 -3792 7836 -3758
rect 7790 -3830 7836 -3792
rect 7790 -3864 7796 -3830
rect 7830 -3864 7836 -3830
rect 7790 -3952 7836 -3864
rect 7984 -3758 8030 -3711
rect 7984 -3792 7990 -3758
rect 8024 -3792 8030 -3758
rect 7984 -3830 8030 -3792
rect 7984 -3864 7990 -3830
rect 8024 -3864 8030 -3830
rect 7984 -3952 8030 -3864
rect 8242 -3758 8288 -3711
rect 8242 -3792 8248 -3758
rect 8282 -3792 8288 -3758
rect 8242 -3830 8288 -3792
rect 8242 -3864 8248 -3830
rect 8282 -3864 8288 -3830
rect 8242 -3952 8288 -3864
rect 8500 -3758 8546 -3711
rect 8500 -3792 8506 -3758
rect 8540 -3792 8546 -3758
rect 8500 -3830 8546 -3792
rect 8500 -3864 8506 -3830
rect 8540 -3864 8546 -3830
rect 8500 -3952 8546 -3864
rect 8758 -3758 8804 -3711
rect 8758 -3792 8764 -3758
rect 8798 -3792 8804 -3758
rect 8758 -3830 8804 -3792
rect 8758 -3864 8764 -3830
rect 8798 -3864 8804 -3830
rect 8758 -3952 8804 -3864
rect 9016 -3758 9062 -3711
rect 9016 -3792 9022 -3758
rect 9056 -3792 9062 -3758
rect 9016 -3830 9062 -3792
rect 9016 -3864 9022 -3830
rect 9056 -3864 9062 -3830
rect 9016 -3952 9062 -3864
rect 9210 -3721 9646 -3683
rect 9210 -3755 9589 -3721
rect 9623 -3755 9646 -3721
rect 9210 -3758 9646 -3755
rect 9210 -3792 9216 -3758
rect 9250 -3792 9474 -3758
rect 9508 -3792 9646 -3758
rect 9210 -3793 9646 -3792
rect 9210 -3827 9589 -3793
rect 9623 -3827 9646 -3793
rect 9210 -3830 9646 -3827
rect 9210 -3864 9216 -3830
rect 9250 -3864 9474 -3830
rect 9508 -3864 9646 -3830
rect 9210 -3865 9646 -3864
rect 9210 -3899 9589 -3865
rect 9623 -3899 9646 -3865
rect 9210 -3937 9646 -3899
rect 9210 -3952 9589 -3937
rect 5265 -3958 9589 -3952
rect 5265 -3971 5438 -3958
rect 5058 -3992 5438 -3971
rect 5472 -3992 5510 -3958
rect 5544 -3992 5889 -3958
rect 5923 -3992 5961 -3958
rect 5995 -3992 6147 -3958
rect 6181 -3992 6219 -3958
rect 6253 -3992 6405 -3958
rect 6439 -3992 6477 -3958
rect 6511 -3992 6663 -3958
rect 6697 -3992 6735 -3958
rect 6769 -3992 7115 -3958
rect 7149 -3992 7187 -3958
rect 7221 -3992 7373 -3958
rect 7407 -3992 7445 -3958
rect 7479 -3992 7631 -3958
rect 7665 -3992 7703 -3958
rect 7737 -3992 8083 -3958
rect 8117 -3992 8155 -3958
rect 8189 -3992 8341 -3958
rect 8375 -3992 8413 -3958
rect 8447 -3992 8599 -3958
rect 8633 -3992 8671 -3958
rect 8705 -3992 8857 -3958
rect 8891 -3992 8929 -3958
rect 8963 -3992 9309 -3958
rect 9343 -3992 9381 -3958
rect 9415 -3971 9589 -3958
rect 9623 -3952 9646 -3937
rect 9623 -3971 9648 -3952
rect 9415 -3992 9648 -3971
rect 847 -4009 9648 -3992
rect 847 -4043 872 -4009
rect 906 -4043 5231 -4009
rect 5265 -4043 9589 -4009
rect 9623 -4043 9648 -4009
rect 847 -4072 9648 -4043
rect 847 -4106 946 -4072
rect 980 -4106 1018 -4072
rect 1052 -4106 1090 -4072
rect 1124 -4106 1162 -4072
rect 1196 -4106 1234 -4072
rect 1268 -4106 1306 -4072
rect 1340 -4106 1378 -4072
rect 1412 -4106 1450 -4072
rect 1484 -4106 1522 -4072
rect 1556 -4106 1594 -4072
rect 1628 -4106 1666 -4072
rect 1700 -4106 1738 -4072
rect 1772 -4106 1810 -4072
rect 1844 -4106 1882 -4072
rect 1916 -4106 1954 -4072
rect 1988 -4106 2026 -4072
rect 2060 -4106 2098 -4072
rect 2132 -4106 2170 -4072
rect 2204 -4106 2242 -4072
rect 2276 -4106 2314 -4072
rect 2348 -4106 2386 -4072
rect 2420 -4106 2458 -4072
rect 2492 -4106 2530 -4072
rect 2564 -4106 2602 -4072
rect 2636 -4106 2674 -4072
rect 2708 -4106 2746 -4072
rect 2780 -4106 2818 -4072
rect 2852 -4106 2890 -4072
rect 2924 -4106 2962 -4072
rect 2996 -4106 3034 -4072
rect 3068 -4106 3106 -4072
rect 3140 -4106 3178 -4072
rect 3212 -4106 3250 -4072
rect 3284 -4106 3322 -4072
rect 3356 -4106 3394 -4072
rect 3428 -4106 3466 -4072
rect 3500 -4106 3538 -4072
rect 3572 -4106 3610 -4072
rect 3644 -4106 3682 -4072
rect 3716 -4106 3754 -4072
rect 3788 -4106 3826 -4072
rect 3860 -4106 3898 -4072
rect 3932 -4106 3970 -4072
rect 4004 -4106 4042 -4072
rect 4076 -4106 4114 -4072
rect 4148 -4106 4186 -4072
rect 4220 -4106 4258 -4072
rect 4292 -4106 4330 -4072
rect 4364 -4106 4402 -4072
rect 4436 -4106 4474 -4072
rect 4508 -4106 4546 -4072
rect 4580 -4106 4618 -4072
rect 4652 -4106 4690 -4072
rect 4724 -4106 4762 -4072
rect 4796 -4106 4834 -4072
rect 4868 -4106 4906 -4072
rect 4940 -4106 4978 -4072
rect 5012 -4106 5050 -4072
rect 5084 -4106 5122 -4072
rect 5156 -4106 5339 -4072
rect 5373 -4106 5411 -4072
rect 5445 -4106 5483 -4072
rect 5517 -4106 5555 -4072
rect 5589 -4106 5627 -4072
rect 5661 -4106 5699 -4072
rect 5733 -4106 5771 -4072
rect 5805 -4106 5843 -4072
rect 5877 -4106 5915 -4072
rect 5949 -4106 5987 -4072
rect 6021 -4106 6059 -4072
rect 6093 -4106 6131 -4072
rect 6165 -4106 6203 -4072
rect 6237 -4106 6275 -4072
rect 6309 -4106 6347 -4072
rect 6381 -4106 6419 -4072
rect 6453 -4106 6491 -4072
rect 6525 -4106 6563 -4072
rect 6597 -4106 6635 -4072
rect 6669 -4106 6707 -4072
rect 6741 -4106 6779 -4072
rect 6813 -4106 6851 -4072
rect 6885 -4106 6923 -4072
rect 6957 -4106 6995 -4072
rect 7029 -4106 7067 -4072
rect 7101 -4106 7139 -4072
rect 7173 -4106 7211 -4072
rect 7245 -4106 7283 -4072
rect 7317 -4106 7355 -4072
rect 7389 -4106 7427 -4072
rect 7461 -4106 7499 -4072
rect 7533 -4106 7571 -4072
rect 7605 -4106 7643 -4072
rect 7677 -4106 7715 -4072
rect 7749 -4106 7787 -4072
rect 7821 -4106 7859 -4072
rect 7893 -4106 7931 -4072
rect 7965 -4106 8003 -4072
rect 8037 -4106 8075 -4072
rect 8109 -4106 8147 -4072
rect 8181 -4106 8219 -4072
rect 8253 -4106 8291 -4072
rect 8325 -4106 8363 -4072
rect 8397 -4106 8435 -4072
rect 8469 -4106 8507 -4072
rect 8541 -4106 8579 -4072
rect 8613 -4106 8651 -4072
rect 8685 -4106 8723 -4072
rect 8757 -4106 8795 -4072
rect 8829 -4106 8867 -4072
rect 8901 -4106 8939 -4072
rect 8973 -4106 9011 -4072
rect 9045 -4106 9083 -4072
rect 9117 -4106 9155 -4072
rect 9189 -4106 9227 -4072
rect 9261 -4106 9299 -4072
rect 9333 -4106 9371 -4072
rect 9405 -4106 9443 -4072
rect 9477 -4106 9515 -4072
rect 9549 -4106 9648 -4072
rect 847 -4135 9648 -4106
rect 847 -4169 872 -4135
rect 906 -4169 5231 -4135
rect 5265 -4169 9589 -4135
rect 9623 -4169 9648 -4135
rect 847 -4186 9648 -4169
rect 847 -4207 1080 -4186
rect 847 -4226 872 -4207
rect 849 -4241 872 -4226
rect 906 -4220 1080 -4207
rect 1114 -4220 1152 -4186
rect 1186 -4220 1532 -4186
rect 1566 -4220 1604 -4186
rect 1638 -4220 1790 -4186
rect 1824 -4220 1862 -4186
rect 1896 -4220 2048 -4186
rect 2082 -4220 2120 -4186
rect 2154 -4220 2306 -4186
rect 2340 -4220 2378 -4186
rect 2412 -4220 2758 -4186
rect 2792 -4220 2830 -4186
rect 2864 -4220 3016 -4186
rect 3050 -4220 3088 -4186
rect 3122 -4220 3274 -4186
rect 3308 -4220 3346 -4186
rect 3380 -4220 3726 -4186
rect 3760 -4220 3798 -4186
rect 3832 -4220 3984 -4186
rect 4018 -4220 4056 -4186
rect 4090 -4220 4242 -4186
rect 4276 -4220 4314 -4186
rect 4348 -4220 4500 -4186
rect 4534 -4220 4572 -4186
rect 4606 -4220 4952 -4186
rect 4986 -4220 5024 -4186
rect 5058 -4207 5438 -4186
rect 5058 -4220 5231 -4207
rect 906 -4226 5231 -4220
rect 906 -4241 1285 -4226
rect 849 -4279 1285 -4241
rect 849 -4313 872 -4279
rect 906 -4313 1285 -4279
rect 849 -4314 1285 -4313
rect 849 -4348 987 -4314
rect 1021 -4348 1245 -4314
rect 1279 -4348 1285 -4314
rect 849 -4351 1285 -4348
rect 849 -4385 872 -4351
rect 906 -4385 1285 -4351
rect 849 -4386 1285 -4385
rect 849 -4420 987 -4386
rect 1021 -4420 1245 -4386
rect 1279 -4420 1285 -4386
rect 849 -4423 1285 -4420
rect 849 -4457 872 -4423
rect 906 -4457 1285 -4423
rect 849 -4495 1285 -4457
rect 1433 -4314 1479 -4226
rect 1433 -4348 1439 -4314
rect 1473 -4348 1479 -4314
rect 1433 -4386 1479 -4348
rect 1433 -4420 1439 -4386
rect 1473 -4420 1479 -4386
rect 1433 -4467 1479 -4420
rect 1691 -4314 1737 -4226
rect 1691 -4348 1697 -4314
rect 1731 -4348 1737 -4314
rect 1691 -4386 1737 -4348
rect 1691 -4420 1697 -4386
rect 1731 -4420 1737 -4386
rect 1691 -4467 1737 -4420
rect 1949 -4314 1995 -4226
rect 1949 -4348 1955 -4314
rect 1989 -4348 1995 -4314
rect 1949 -4386 1995 -4348
rect 1949 -4420 1955 -4386
rect 1989 -4420 1995 -4386
rect 1949 -4467 1995 -4420
rect 2207 -4314 2253 -4226
rect 2207 -4348 2213 -4314
rect 2247 -4348 2253 -4314
rect 2207 -4386 2253 -4348
rect 2207 -4420 2213 -4386
rect 2247 -4420 2253 -4386
rect 2207 -4467 2253 -4420
rect 2465 -4314 2511 -4226
rect 2465 -4348 2471 -4314
rect 2505 -4348 2511 -4314
rect 2465 -4386 2511 -4348
rect 2465 -4420 2471 -4386
rect 2505 -4420 2511 -4386
rect 2465 -4467 2511 -4420
rect 2659 -4314 2705 -4226
rect 2659 -4348 2665 -4314
rect 2699 -4348 2705 -4314
rect 2659 -4386 2705 -4348
rect 2659 -4420 2665 -4386
rect 2699 -4420 2705 -4386
rect 2659 -4467 2705 -4420
rect 2917 -4314 2963 -4226
rect 2917 -4348 2923 -4314
rect 2957 -4348 2963 -4314
rect 2917 -4386 2963 -4348
rect 2917 -4420 2923 -4386
rect 2957 -4420 2963 -4386
rect 2917 -4467 2963 -4420
rect 3175 -4314 3221 -4226
rect 3175 -4348 3181 -4314
rect 3215 -4348 3221 -4314
rect 3175 -4386 3221 -4348
rect 3175 -4420 3181 -4386
rect 3215 -4420 3221 -4386
rect 3175 -4467 3221 -4420
rect 3433 -4314 3479 -4226
rect 3433 -4348 3439 -4314
rect 3473 -4348 3479 -4314
rect 3433 -4386 3479 -4348
rect 3433 -4420 3439 -4386
rect 3473 -4420 3479 -4386
rect 3433 -4467 3479 -4420
rect 3627 -4314 3673 -4226
rect 3627 -4348 3633 -4314
rect 3667 -4348 3673 -4314
rect 3627 -4386 3673 -4348
rect 3627 -4420 3633 -4386
rect 3667 -4420 3673 -4386
rect 3627 -4467 3673 -4420
rect 3885 -4314 3931 -4226
rect 3885 -4348 3891 -4314
rect 3925 -4348 3931 -4314
rect 3885 -4386 3931 -4348
rect 3885 -4420 3891 -4386
rect 3925 -4420 3931 -4386
rect 3885 -4467 3931 -4420
rect 4143 -4314 4189 -4226
rect 4143 -4348 4149 -4314
rect 4183 -4348 4189 -4314
rect 4143 -4386 4189 -4348
rect 4143 -4420 4149 -4386
rect 4183 -4420 4189 -4386
rect 4143 -4467 4189 -4420
rect 4401 -4314 4447 -4226
rect 4401 -4348 4407 -4314
rect 4441 -4348 4447 -4314
rect 4401 -4386 4447 -4348
rect 4401 -4420 4407 -4386
rect 4441 -4420 4447 -4386
rect 4401 -4467 4447 -4420
rect 4659 -4314 4705 -4226
rect 4659 -4348 4665 -4314
rect 4699 -4348 4705 -4314
rect 4659 -4386 4705 -4348
rect 4659 -4420 4665 -4386
rect 4699 -4420 4705 -4386
rect 4659 -4467 4705 -4420
rect 4853 -4241 5231 -4226
rect 5265 -4220 5438 -4207
rect 5472 -4220 5510 -4186
rect 5544 -4220 5889 -4186
rect 5923 -4220 5961 -4186
rect 5995 -4220 6147 -4186
rect 6181 -4220 6219 -4186
rect 6253 -4220 6405 -4186
rect 6439 -4220 6477 -4186
rect 6511 -4220 6663 -4186
rect 6697 -4220 6735 -4186
rect 6769 -4220 7115 -4186
rect 7149 -4220 7187 -4186
rect 7221 -4220 7373 -4186
rect 7407 -4220 7445 -4186
rect 7479 -4220 7631 -4186
rect 7665 -4220 7703 -4186
rect 7737 -4220 8083 -4186
rect 8117 -4220 8155 -4186
rect 8189 -4220 8341 -4186
rect 8375 -4220 8413 -4186
rect 8447 -4220 8599 -4186
rect 8633 -4220 8671 -4186
rect 8705 -4220 8857 -4186
rect 8891 -4220 8929 -4186
rect 8963 -4220 9309 -4186
rect 9343 -4220 9381 -4186
rect 9415 -4207 9648 -4186
rect 9415 -4220 9589 -4207
rect 5265 -4226 9589 -4220
rect 5265 -4241 5643 -4226
rect 4853 -4279 5643 -4241
rect 4853 -4313 5231 -4279
rect 5265 -4313 5643 -4279
rect 4853 -4314 5643 -4313
rect 4853 -4348 4859 -4314
rect 4893 -4348 5117 -4314
rect 5151 -4348 5345 -4314
rect 5379 -4348 5603 -4314
rect 5637 -4348 5643 -4314
rect 4853 -4351 5643 -4348
rect 4853 -4385 5231 -4351
rect 5265 -4385 5643 -4351
rect 4853 -4386 5643 -4385
rect 4853 -4420 4859 -4386
rect 4893 -4420 5117 -4386
rect 5151 -4420 5345 -4386
rect 5379 -4420 5603 -4386
rect 5637 -4420 5643 -4386
rect 4853 -4423 5643 -4420
rect 4853 -4457 5231 -4423
rect 5265 -4457 5643 -4423
rect 849 -4529 872 -4495
rect 906 -4529 1285 -4495
rect 849 -4567 1285 -4529
rect 849 -4601 872 -4567
rect 906 -4601 1285 -4567
rect 4853 -4495 5643 -4457
rect 5790 -4314 5836 -4226
rect 5790 -4348 5796 -4314
rect 5830 -4348 5836 -4314
rect 5790 -4386 5836 -4348
rect 5790 -4420 5796 -4386
rect 5830 -4420 5836 -4386
rect 5790 -4467 5836 -4420
rect 6048 -4314 6094 -4226
rect 6048 -4348 6054 -4314
rect 6088 -4348 6094 -4314
rect 6048 -4386 6094 -4348
rect 6048 -4420 6054 -4386
rect 6088 -4420 6094 -4386
rect 6048 -4467 6094 -4420
rect 6306 -4314 6352 -4226
rect 6306 -4348 6312 -4314
rect 6346 -4348 6352 -4314
rect 6306 -4386 6352 -4348
rect 6306 -4420 6312 -4386
rect 6346 -4420 6352 -4386
rect 6306 -4467 6352 -4420
rect 6564 -4314 6610 -4226
rect 6564 -4348 6570 -4314
rect 6604 -4348 6610 -4314
rect 6564 -4386 6610 -4348
rect 6564 -4420 6570 -4386
rect 6604 -4420 6610 -4386
rect 6564 -4467 6610 -4420
rect 6822 -4314 6868 -4226
rect 6822 -4348 6828 -4314
rect 6862 -4348 6868 -4314
rect 6822 -4386 6868 -4348
rect 6822 -4420 6828 -4386
rect 6862 -4420 6868 -4386
rect 6822 -4467 6868 -4420
rect 7016 -4314 7062 -4226
rect 7016 -4348 7022 -4314
rect 7056 -4348 7062 -4314
rect 7016 -4386 7062 -4348
rect 7016 -4420 7022 -4386
rect 7056 -4420 7062 -4386
rect 7016 -4467 7062 -4420
rect 7274 -4314 7320 -4226
rect 7274 -4348 7280 -4314
rect 7314 -4348 7320 -4314
rect 7274 -4386 7320 -4348
rect 7274 -4420 7280 -4386
rect 7314 -4420 7320 -4386
rect 7274 -4467 7320 -4420
rect 7532 -4314 7578 -4226
rect 7532 -4348 7538 -4314
rect 7572 -4348 7578 -4314
rect 7532 -4386 7578 -4348
rect 7532 -4420 7538 -4386
rect 7572 -4420 7578 -4386
rect 7532 -4467 7578 -4420
rect 7790 -4314 7836 -4226
rect 7790 -4348 7796 -4314
rect 7830 -4348 7836 -4314
rect 7790 -4386 7836 -4348
rect 7790 -4420 7796 -4386
rect 7830 -4420 7836 -4386
rect 7790 -4467 7836 -4420
rect 7984 -4314 8030 -4226
rect 7984 -4348 7990 -4314
rect 8024 -4348 8030 -4314
rect 7984 -4386 8030 -4348
rect 7984 -4420 7990 -4386
rect 8024 -4420 8030 -4386
rect 7984 -4467 8030 -4420
rect 8242 -4314 8288 -4226
rect 8242 -4348 8248 -4314
rect 8282 -4348 8288 -4314
rect 8242 -4386 8288 -4348
rect 8242 -4420 8248 -4386
rect 8282 -4420 8288 -4386
rect 8242 -4467 8288 -4420
rect 8500 -4314 8546 -4226
rect 8500 -4348 8506 -4314
rect 8540 -4348 8546 -4314
rect 8500 -4386 8546 -4348
rect 8500 -4420 8506 -4386
rect 8540 -4420 8546 -4386
rect 8500 -4467 8546 -4420
rect 8758 -4314 8804 -4226
rect 8758 -4348 8764 -4314
rect 8798 -4348 8804 -4314
rect 8758 -4386 8804 -4348
rect 8758 -4420 8764 -4386
rect 8798 -4420 8804 -4386
rect 8758 -4467 8804 -4420
rect 9016 -4314 9062 -4226
rect 9016 -4348 9022 -4314
rect 9056 -4348 9062 -4314
rect 9016 -4386 9062 -4348
rect 9016 -4420 9022 -4386
rect 9056 -4420 9062 -4386
rect 9016 -4467 9062 -4420
rect 9210 -4241 9589 -4226
rect 9623 -4226 9648 -4207
rect 9623 -4241 9646 -4226
rect 9210 -4279 9646 -4241
rect 9210 -4313 9589 -4279
rect 9623 -4313 9646 -4279
rect 9210 -4314 9646 -4313
rect 9210 -4348 9216 -4314
rect 9250 -4348 9474 -4314
rect 9508 -4348 9646 -4314
rect 9210 -4351 9646 -4348
rect 9210 -4385 9589 -4351
rect 9623 -4385 9646 -4351
rect 9210 -4386 9646 -4385
rect 9210 -4420 9216 -4386
rect 9250 -4420 9474 -4386
rect 9508 -4420 9646 -4386
rect 9210 -4423 9646 -4420
rect 9210 -4457 9589 -4423
rect 9623 -4457 9646 -4423
rect 4853 -4529 5231 -4495
rect 5265 -4529 5643 -4495
rect 4853 -4567 5643 -4529
rect 849 -4639 1285 -4601
rect 849 -4673 872 -4639
rect 906 -4673 1285 -4639
rect 2843 -4592 3039 -4584
rect 2843 -4644 2850 -4592
rect 2902 -4644 2914 -4592
rect 2966 -4644 2978 -4592
rect 3030 -4644 3039 -4592
rect 2843 -4654 3039 -4644
rect 3361 -4592 3557 -4584
rect 3361 -4644 3368 -4592
rect 3420 -4644 3432 -4592
rect 3484 -4644 3496 -4592
rect 3548 -4644 3557 -4592
rect 3361 -4654 3557 -4644
rect 4853 -4601 5231 -4567
rect 5265 -4601 5643 -4567
rect 9210 -4495 9646 -4457
rect 9210 -4529 9589 -4495
rect 9623 -4529 9646 -4495
rect 9210 -4567 9646 -4529
rect 4853 -4639 5643 -4601
rect 849 -4711 1285 -4673
rect 849 -4745 872 -4711
rect 906 -4745 1285 -4711
rect 849 -4783 1285 -4745
rect 849 -4817 872 -4783
rect 906 -4817 1285 -4783
rect 849 -4855 1285 -4817
rect 1355 -4761 1551 -4753
rect 1355 -4813 1364 -4761
rect 1416 -4813 1428 -4761
rect 1480 -4813 1492 -4761
rect 1544 -4813 1551 -4761
rect 1355 -4823 1551 -4813
rect 1873 -4761 2069 -4753
rect 1873 -4813 1882 -4761
rect 1934 -4813 1946 -4761
rect 1998 -4813 2010 -4761
rect 2062 -4813 2069 -4761
rect 1873 -4823 2069 -4813
rect 2389 -4761 2585 -4753
rect 2389 -4813 2398 -4761
rect 2450 -4813 2462 -4761
rect 2514 -4813 2526 -4761
rect 2578 -4813 2585 -4761
rect 2389 -4823 2585 -4813
rect 849 -4889 872 -4855
rect 906 -4889 1285 -4855
rect 849 -4927 1285 -4889
rect 849 -4961 872 -4927
rect 906 -4961 1285 -4927
rect 849 -4999 1285 -4961
rect 849 -5033 872 -4999
rect 906 -5033 1285 -4999
rect 849 -5071 1285 -5033
rect 849 -5105 872 -5071
rect 906 -5105 1285 -5071
rect 849 -5143 1285 -5105
rect 849 -5177 872 -5143
rect 906 -5177 1285 -5143
rect 849 -5215 1285 -5177
rect 849 -5249 872 -5215
rect 906 -5249 1285 -5215
rect 849 -5287 1285 -5249
rect 849 -5321 872 -5287
rect 906 -5304 1285 -5287
rect 906 -5321 987 -5304
rect 849 -5338 987 -5321
rect 1021 -5338 1245 -5304
rect 1279 -5338 1285 -5304
rect 849 -5359 1285 -5338
rect 849 -5393 872 -5359
rect 906 -5376 1285 -5359
rect 906 -5393 987 -5376
rect 849 -5410 987 -5393
rect 1021 -5410 1245 -5376
rect 1279 -5410 1285 -5376
rect 849 -5431 1285 -5410
rect 849 -5465 872 -5431
rect 906 -5465 1285 -5431
rect 1433 -5304 1479 -4823
rect 1615 -5093 1811 -5085
rect 1615 -5145 1624 -5093
rect 1676 -5145 1688 -5093
rect 1740 -5145 1752 -5093
rect 1804 -5145 1811 -5093
rect 1615 -5155 1811 -5145
rect 1433 -5338 1439 -5304
rect 1473 -5338 1479 -5304
rect 1433 -5376 1479 -5338
rect 1433 -5410 1439 -5376
rect 1473 -5410 1479 -5376
rect 1433 -5457 1479 -5410
rect 1691 -5304 1737 -5155
rect 1691 -5338 1697 -5304
rect 1731 -5338 1737 -5304
rect 1691 -5376 1737 -5338
rect 1691 -5410 1697 -5376
rect 1731 -5410 1737 -5376
rect 1691 -5457 1737 -5410
rect 1949 -5304 1995 -4823
rect 2132 -5093 2328 -5085
rect 2132 -5145 2141 -5093
rect 2193 -5145 2205 -5093
rect 2257 -5145 2269 -5093
rect 2321 -5145 2328 -5093
rect 2132 -5155 2328 -5145
rect 1949 -5338 1955 -5304
rect 1989 -5338 1995 -5304
rect 1949 -5376 1995 -5338
rect 1949 -5410 1955 -5376
rect 1989 -5410 1995 -5376
rect 1949 -5457 1995 -5410
rect 2207 -5304 2253 -5155
rect 2207 -5338 2213 -5304
rect 2247 -5338 2253 -5304
rect 2207 -5376 2253 -5338
rect 2207 -5410 2213 -5376
rect 2247 -5410 2253 -5376
rect 2207 -5457 2253 -5410
rect 2465 -5304 2511 -4823
rect 2586 -4924 2782 -4916
rect 2586 -4976 2593 -4924
rect 2645 -4976 2657 -4924
rect 2709 -4976 2721 -4924
rect 2773 -4976 2782 -4924
rect 2586 -4986 2782 -4976
rect 2465 -5338 2471 -5304
rect 2505 -5338 2511 -5304
rect 2465 -5376 2511 -5338
rect 2465 -5410 2471 -5376
rect 2505 -5410 2511 -5376
rect 2465 -5457 2511 -5410
rect 2659 -5304 2705 -4986
rect 2659 -5338 2665 -5304
rect 2699 -5338 2705 -5304
rect 2659 -5376 2705 -5338
rect 2659 -5410 2665 -5376
rect 2699 -5410 2705 -5376
rect 2659 -5457 2705 -5410
rect 2917 -5304 2963 -4654
rect 3103 -4924 3299 -4916
rect 3103 -4976 3110 -4924
rect 3162 -4976 3174 -4924
rect 3226 -4976 3238 -4924
rect 3290 -4976 3299 -4924
rect 3103 -4986 3299 -4976
rect 2917 -5338 2923 -5304
rect 2957 -5338 2963 -5304
rect 2917 -5376 2963 -5338
rect 2917 -5410 2923 -5376
rect 2957 -5410 2963 -5376
rect 2917 -5457 2963 -5410
rect 3175 -5304 3221 -4986
rect 3175 -5338 3181 -5304
rect 3215 -5338 3221 -5304
rect 3175 -5376 3221 -5338
rect 3175 -5410 3181 -5376
rect 3215 -5410 3221 -5376
rect 3175 -5457 3221 -5410
rect 3433 -5304 3479 -4654
rect 4853 -4673 5231 -4639
rect 5265 -4673 5643 -4639
rect 6939 -4592 7135 -4584
rect 6939 -4644 6948 -4592
rect 7000 -4644 7012 -4592
rect 7064 -4644 7076 -4592
rect 7128 -4644 7135 -4592
rect 6939 -4654 7135 -4644
rect 7456 -4592 7652 -4584
rect 7456 -4644 7465 -4592
rect 7517 -4644 7529 -4592
rect 7581 -4644 7593 -4592
rect 7645 -4644 7652 -4592
rect 7456 -4654 7652 -4644
rect 9210 -4601 9589 -4567
rect 9623 -4601 9646 -4567
rect 9210 -4639 9646 -4601
rect 4853 -4711 5643 -4673
rect 4853 -4745 5231 -4711
rect 5265 -4745 5643 -4711
rect 3550 -4761 3746 -4753
rect 3550 -4813 3559 -4761
rect 3611 -4813 3623 -4761
rect 3675 -4813 3687 -4761
rect 3739 -4813 3746 -4761
rect 3550 -4823 3746 -4813
rect 4067 -4761 4263 -4753
rect 4067 -4813 4076 -4761
rect 4128 -4813 4140 -4761
rect 4192 -4813 4204 -4761
rect 4256 -4813 4263 -4761
rect 4067 -4823 4263 -4813
rect 4582 -4761 4778 -4753
rect 4582 -4813 4591 -4761
rect 4643 -4813 4655 -4761
rect 4707 -4813 4719 -4761
rect 4771 -4813 4778 -4761
rect 4582 -4823 4778 -4813
rect 4853 -4783 5643 -4745
rect 4853 -4817 5231 -4783
rect 5265 -4817 5643 -4783
rect 3433 -5338 3439 -5304
rect 3473 -5338 3479 -5304
rect 3433 -5376 3479 -5338
rect 3433 -5410 3439 -5376
rect 3473 -5410 3479 -5376
rect 3433 -5457 3479 -5410
rect 3627 -5304 3673 -4823
rect 3809 -5093 4005 -5085
rect 3809 -5145 3818 -5093
rect 3870 -5145 3882 -5093
rect 3934 -5145 3946 -5093
rect 3998 -5145 4005 -5093
rect 3809 -5155 4005 -5145
rect 3627 -5338 3633 -5304
rect 3667 -5338 3673 -5304
rect 3627 -5376 3673 -5338
rect 3627 -5410 3633 -5376
rect 3667 -5410 3673 -5376
rect 3627 -5457 3673 -5410
rect 3885 -5304 3931 -5155
rect 3885 -5338 3891 -5304
rect 3925 -5338 3931 -5304
rect 3885 -5376 3931 -5338
rect 3885 -5410 3891 -5376
rect 3925 -5410 3931 -5376
rect 3885 -5457 3931 -5410
rect 4143 -5304 4189 -4823
rect 4326 -5093 4522 -5085
rect 4326 -5145 4335 -5093
rect 4387 -5145 4399 -5093
rect 4451 -5145 4463 -5093
rect 4515 -5145 4522 -5093
rect 4326 -5155 4522 -5145
rect 4143 -5338 4149 -5304
rect 4183 -5338 4189 -5304
rect 4143 -5376 4189 -5338
rect 4143 -5410 4149 -5376
rect 4183 -5410 4189 -5376
rect 4143 -5457 4189 -5410
rect 4401 -5304 4447 -5155
rect 4401 -5338 4407 -5304
rect 4441 -5338 4447 -5304
rect 4401 -5376 4447 -5338
rect 4401 -5410 4407 -5376
rect 4441 -5410 4447 -5376
rect 4401 -5457 4447 -5410
rect 4659 -5304 4705 -4823
rect 4659 -5338 4665 -5304
rect 4699 -5338 4705 -5304
rect 4659 -5376 4705 -5338
rect 4659 -5410 4665 -5376
rect 4699 -5410 4705 -5376
rect 4659 -5457 4705 -5410
rect 4853 -4855 5643 -4817
rect 5717 -4761 5913 -4753
rect 5717 -4813 5724 -4761
rect 5776 -4813 5788 -4761
rect 5840 -4813 5852 -4761
rect 5904 -4813 5913 -4761
rect 5717 -4823 5913 -4813
rect 6232 -4761 6428 -4753
rect 6232 -4813 6239 -4761
rect 6291 -4813 6303 -4761
rect 6355 -4813 6367 -4761
rect 6419 -4813 6428 -4761
rect 6232 -4823 6428 -4813
rect 6749 -4761 6945 -4753
rect 6749 -4813 6756 -4761
rect 6808 -4813 6820 -4761
rect 6872 -4813 6884 -4761
rect 6936 -4813 6945 -4761
rect 6749 -4823 6945 -4813
rect 4853 -4889 5231 -4855
rect 5265 -4889 5643 -4855
rect 4853 -4927 5643 -4889
rect 4853 -4961 5231 -4927
rect 5265 -4961 5643 -4927
rect 4853 -4999 5643 -4961
rect 4853 -5033 5231 -4999
rect 5265 -5033 5643 -4999
rect 4853 -5071 5643 -5033
rect 4853 -5105 5231 -5071
rect 5265 -5105 5643 -5071
rect 4853 -5143 5643 -5105
rect 4853 -5177 5231 -5143
rect 5265 -5177 5643 -5143
rect 4853 -5215 5643 -5177
rect 4853 -5249 5231 -5215
rect 5265 -5249 5643 -5215
rect 4853 -5287 5643 -5249
rect 4853 -5304 5231 -5287
rect 4853 -5338 4859 -5304
rect 4893 -5338 5117 -5304
rect 5151 -5321 5231 -5304
rect 5265 -5304 5643 -5287
rect 5265 -5321 5345 -5304
rect 5151 -5338 5345 -5321
rect 5379 -5338 5603 -5304
rect 5637 -5338 5643 -5304
rect 4853 -5359 5643 -5338
rect 4853 -5376 5231 -5359
rect 4853 -5410 4859 -5376
rect 4893 -5410 5117 -5376
rect 5151 -5393 5231 -5376
rect 5265 -5376 5643 -5359
rect 5265 -5393 5345 -5376
rect 5151 -5410 5345 -5393
rect 5379 -5410 5603 -5376
rect 5637 -5410 5643 -5376
rect 4853 -5431 5643 -5410
rect 849 -5503 1285 -5465
rect 4853 -5465 5231 -5431
rect 5265 -5465 5643 -5431
rect 5790 -5304 5836 -4823
rect 5973 -5093 6169 -5085
rect 5973 -5145 5980 -5093
rect 6032 -5145 6044 -5093
rect 6096 -5145 6108 -5093
rect 6160 -5145 6169 -5093
rect 5973 -5155 6169 -5145
rect 5790 -5338 5796 -5304
rect 5830 -5338 5836 -5304
rect 5790 -5376 5836 -5338
rect 5790 -5410 5796 -5376
rect 5830 -5410 5836 -5376
rect 5790 -5457 5836 -5410
rect 6048 -5304 6094 -5155
rect 6048 -5338 6054 -5304
rect 6088 -5338 6094 -5304
rect 6048 -5376 6094 -5338
rect 6048 -5410 6054 -5376
rect 6088 -5410 6094 -5376
rect 6048 -5457 6094 -5410
rect 6306 -5304 6352 -4823
rect 6490 -5093 6686 -5085
rect 6490 -5145 6497 -5093
rect 6549 -5145 6561 -5093
rect 6613 -5145 6625 -5093
rect 6677 -5145 6686 -5093
rect 6490 -5155 6686 -5145
rect 6306 -5338 6312 -5304
rect 6346 -5338 6352 -5304
rect 6306 -5376 6352 -5338
rect 6306 -5410 6312 -5376
rect 6346 -5410 6352 -5376
rect 6306 -5457 6352 -5410
rect 6564 -5304 6610 -5155
rect 6564 -5338 6570 -5304
rect 6604 -5338 6610 -5304
rect 6564 -5376 6610 -5338
rect 6564 -5410 6570 -5376
rect 6604 -5410 6610 -5376
rect 6564 -5457 6610 -5410
rect 6822 -5304 6868 -4823
rect 6822 -5338 6828 -5304
rect 6862 -5338 6868 -5304
rect 6822 -5376 6868 -5338
rect 6822 -5410 6828 -5376
rect 6862 -5410 6868 -5376
rect 6822 -5457 6868 -5410
rect 7016 -5304 7062 -4654
rect 7196 -4924 7392 -4916
rect 7196 -4976 7205 -4924
rect 7257 -4976 7269 -4924
rect 7321 -4976 7333 -4924
rect 7385 -4976 7392 -4924
rect 7196 -4986 7392 -4976
rect 7016 -5338 7022 -5304
rect 7056 -5338 7062 -5304
rect 7016 -5376 7062 -5338
rect 7016 -5410 7022 -5376
rect 7056 -5410 7062 -5376
rect 7016 -5457 7062 -5410
rect 7274 -5304 7320 -4986
rect 7274 -5338 7280 -5304
rect 7314 -5338 7320 -5304
rect 7274 -5376 7320 -5338
rect 7274 -5410 7280 -5376
rect 7314 -5410 7320 -5376
rect 7274 -5457 7320 -5410
rect 7532 -5304 7578 -4654
rect 9210 -4673 9589 -4639
rect 9623 -4673 9646 -4639
rect 9210 -4711 9646 -4673
rect 9210 -4745 9589 -4711
rect 9623 -4745 9646 -4711
rect 7910 -4761 8106 -4753
rect 7910 -4813 7917 -4761
rect 7969 -4813 7981 -4761
rect 8033 -4813 8045 -4761
rect 8097 -4813 8106 -4761
rect 7910 -4823 8106 -4813
rect 8427 -4761 8623 -4753
rect 8427 -4813 8434 -4761
rect 8486 -4813 8498 -4761
rect 8550 -4813 8562 -4761
rect 8614 -4813 8623 -4761
rect 8427 -4823 8623 -4813
rect 8944 -4761 9140 -4753
rect 8944 -4813 8951 -4761
rect 9003 -4813 9015 -4761
rect 9067 -4813 9079 -4761
rect 9131 -4813 9140 -4761
rect 8944 -4823 9140 -4813
rect 9210 -4783 9646 -4745
rect 9210 -4817 9589 -4783
rect 9623 -4817 9646 -4783
rect 7713 -4924 7909 -4916
rect 7713 -4976 7722 -4924
rect 7774 -4976 7786 -4924
rect 7838 -4976 7850 -4924
rect 7902 -4976 7909 -4924
rect 7713 -4986 7909 -4976
rect 7532 -5338 7538 -5304
rect 7572 -5338 7578 -5304
rect 7532 -5376 7578 -5338
rect 7532 -5410 7538 -5376
rect 7572 -5410 7578 -5376
rect 7532 -5457 7578 -5410
rect 7790 -5304 7836 -4986
rect 7790 -5338 7796 -5304
rect 7830 -5338 7836 -5304
rect 7790 -5376 7836 -5338
rect 7790 -5410 7796 -5376
rect 7830 -5410 7836 -5376
rect 7790 -5457 7836 -5410
rect 7984 -5304 8030 -4823
rect 8167 -5093 8363 -5085
rect 8167 -5145 8174 -5093
rect 8226 -5145 8238 -5093
rect 8290 -5145 8302 -5093
rect 8354 -5145 8363 -5093
rect 8167 -5155 8363 -5145
rect 7984 -5338 7990 -5304
rect 8024 -5338 8030 -5304
rect 7984 -5376 8030 -5338
rect 7984 -5410 7990 -5376
rect 8024 -5410 8030 -5376
rect 7984 -5457 8030 -5410
rect 8242 -5304 8288 -5155
rect 8242 -5338 8248 -5304
rect 8282 -5338 8288 -5304
rect 8242 -5376 8288 -5338
rect 8242 -5410 8248 -5376
rect 8282 -5410 8288 -5376
rect 8242 -5457 8288 -5410
rect 8500 -5304 8546 -4823
rect 8685 -5093 8881 -5085
rect 8685 -5145 8692 -5093
rect 8744 -5145 8756 -5093
rect 8808 -5145 8820 -5093
rect 8872 -5145 8881 -5093
rect 8685 -5155 8881 -5145
rect 8500 -5338 8506 -5304
rect 8540 -5338 8546 -5304
rect 8500 -5376 8546 -5338
rect 8500 -5410 8506 -5376
rect 8540 -5410 8546 -5376
rect 8500 -5457 8546 -5410
rect 8758 -5304 8804 -5155
rect 8758 -5338 8764 -5304
rect 8798 -5338 8804 -5304
rect 8758 -5376 8804 -5338
rect 8758 -5410 8764 -5376
rect 8798 -5410 8804 -5376
rect 8758 -5457 8804 -5410
rect 9016 -5304 9062 -4823
rect 9016 -5338 9022 -5304
rect 9056 -5338 9062 -5304
rect 9016 -5376 9062 -5338
rect 9016 -5410 9022 -5376
rect 9056 -5410 9062 -5376
rect 9016 -5457 9062 -5410
rect 9210 -4855 9646 -4817
rect 9210 -4889 9589 -4855
rect 9623 -4889 9646 -4855
rect 9210 -4927 9646 -4889
rect 9210 -4961 9589 -4927
rect 9623 -4961 9646 -4927
rect 9210 -4999 9646 -4961
rect 9210 -5033 9589 -4999
rect 9623 -5033 9646 -4999
rect 9210 -5071 9646 -5033
rect 9210 -5105 9589 -5071
rect 9623 -5105 9646 -5071
rect 9210 -5143 9646 -5105
rect 9210 -5177 9589 -5143
rect 9623 -5177 9646 -5143
rect 9210 -5215 9646 -5177
rect 9210 -5249 9589 -5215
rect 9623 -5249 9646 -5215
rect 9210 -5287 9646 -5249
rect 9210 -5304 9589 -5287
rect 9210 -5338 9216 -5304
rect 9250 -5338 9474 -5304
rect 9508 -5321 9589 -5304
rect 9623 -5321 9646 -5287
rect 9508 -5338 9646 -5321
rect 9210 -5359 9646 -5338
rect 9210 -5376 9589 -5359
rect 9210 -5410 9216 -5376
rect 9250 -5410 9474 -5376
rect 9508 -5393 9589 -5376
rect 9623 -5393 9646 -5359
rect 9508 -5410 9646 -5393
rect 9210 -5431 9646 -5410
rect 849 -5537 872 -5503
rect 906 -5504 1285 -5503
rect 906 -5537 1080 -5504
rect 849 -5538 1080 -5537
rect 1114 -5538 1152 -5504
rect 1186 -5538 1285 -5504
rect 849 -5575 1285 -5538
rect 849 -5609 872 -5575
rect 906 -5609 1285 -5575
rect 849 -5647 1285 -5609
rect 849 -5681 872 -5647
rect 906 -5681 1285 -5647
rect 849 -5719 1285 -5681
rect 849 -5753 872 -5719
rect 906 -5753 1285 -5719
rect 849 -5791 1285 -5753
rect 1489 -5504 2455 -5498
rect 1489 -5538 1532 -5504
rect 1566 -5519 1604 -5504
rect 1638 -5519 1790 -5504
rect 1824 -5519 1862 -5504
rect 1896 -5519 2048 -5504
rect 2082 -5519 2120 -5504
rect 2154 -5519 2306 -5504
rect 2340 -5519 2378 -5504
rect 1489 -5571 1539 -5538
rect 1591 -5571 1603 -5519
rect 1655 -5571 1667 -5519
rect 1719 -5571 1735 -5519
rect 1787 -5538 1790 -5519
rect 1851 -5538 1862 -5519
rect 1787 -5571 1799 -5538
rect 1851 -5571 1863 -5538
rect 1915 -5571 2025 -5519
rect 2082 -5538 2089 -5519
rect 2077 -5571 2089 -5538
rect 2141 -5571 2153 -5538
rect 2205 -5571 2221 -5519
rect 2273 -5571 2285 -5519
rect 2340 -5538 2349 -5519
rect 2412 -5538 2455 -5504
rect 2337 -5571 2349 -5538
rect 2401 -5571 2455 -5538
rect 1489 -5697 2455 -5571
rect 1489 -5749 1539 -5697
rect 1591 -5749 1603 -5697
rect 1655 -5749 1667 -5697
rect 1719 -5749 1735 -5697
rect 1787 -5749 1799 -5697
rect 1851 -5749 1863 -5697
rect 1915 -5749 2025 -5697
rect 2077 -5749 2089 -5697
rect 2141 -5749 2153 -5697
rect 2205 -5749 2221 -5697
rect 2273 -5749 2285 -5697
rect 2337 -5749 2349 -5697
rect 2401 -5749 2455 -5697
rect 1489 -5768 2455 -5749
rect 2532 -5504 3606 -5498
rect 2532 -5538 2758 -5504
rect 2792 -5538 2830 -5504
rect 2864 -5538 3016 -5504
rect 3050 -5538 3088 -5504
rect 3122 -5538 3274 -5504
rect 3308 -5538 3346 -5504
rect 3380 -5538 3606 -5504
rect 2532 -5586 3606 -5538
rect 849 -5825 872 -5791
rect 906 -5825 1285 -5791
rect 2532 -5818 2593 -5586
rect 849 -5863 1285 -5825
rect 849 -5897 872 -5863
rect 906 -5866 1285 -5863
rect 906 -5897 1080 -5866
rect 849 -5900 1080 -5897
rect 1114 -5900 1152 -5866
rect 1186 -5900 1285 -5866
rect 849 -5935 1285 -5900
rect 1489 -5836 2593 -5818
rect 1489 -5866 1539 -5836
rect 1489 -5900 1532 -5866
rect 1591 -5888 1603 -5836
rect 1655 -5888 1667 -5836
rect 1719 -5888 1735 -5836
rect 1787 -5866 1799 -5836
rect 1851 -5866 1863 -5836
rect 1787 -5888 1790 -5866
rect 1851 -5888 1862 -5866
rect 1915 -5888 2025 -5836
rect 2077 -5866 2089 -5836
rect 2141 -5866 2153 -5836
rect 2082 -5888 2089 -5866
rect 2205 -5888 2221 -5836
rect 2273 -5888 2285 -5836
rect 2337 -5866 2349 -5836
rect 2401 -5866 2593 -5836
rect 2340 -5888 2349 -5866
rect 1566 -5900 1604 -5888
rect 1638 -5900 1790 -5888
rect 1824 -5900 1862 -5888
rect 1896 -5900 2048 -5888
rect 2082 -5900 2120 -5888
rect 2154 -5900 2306 -5888
rect 2340 -5900 2378 -5888
rect 2412 -5900 2593 -5866
rect 1489 -5906 2593 -5900
rect 2715 -5697 3423 -5680
rect 2715 -5749 2749 -5697
rect 2801 -5749 2813 -5697
rect 2865 -5749 2877 -5697
rect 2929 -5749 2945 -5697
rect 2997 -5749 3009 -5697
rect 3061 -5749 3073 -5697
rect 3125 -5749 3137 -5697
rect 3189 -5749 3205 -5697
rect 3257 -5749 3269 -5697
rect 3321 -5749 3333 -5697
rect 3385 -5749 3423 -5697
rect 2715 -5866 3423 -5749
rect 2715 -5900 2758 -5866
rect 2792 -5900 2830 -5866
rect 2864 -5900 3016 -5866
rect 3050 -5900 3088 -5866
rect 3122 -5900 3274 -5866
rect 3308 -5900 3346 -5866
rect 3380 -5900 3423 -5866
rect 2715 -5906 3423 -5900
rect 3545 -5818 3606 -5586
rect 3683 -5504 4649 -5498
rect 3683 -5538 3726 -5504
rect 3760 -5519 3798 -5504
rect 3832 -5519 3984 -5504
rect 4018 -5519 4056 -5504
rect 4090 -5519 4242 -5504
rect 4276 -5519 4314 -5504
rect 4348 -5519 4500 -5504
rect 4534 -5519 4572 -5504
rect 3789 -5538 3798 -5519
rect 3683 -5571 3737 -5538
rect 3789 -5571 3801 -5538
rect 3853 -5571 3865 -5519
rect 3917 -5571 3933 -5519
rect 4049 -5538 4056 -5519
rect 3985 -5571 3997 -5538
rect 4049 -5571 4061 -5538
rect 4113 -5571 4223 -5519
rect 4276 -5538 4287 -5519
rect 4348 -5538 4351 -5519
rect 4275 -5571 4287 -5538
rect 4339 -5571 4351 -5538
rect 4403 -5571 4419 -5519
rect 4471 -5571 4483 -5519
rect 4535 -5571 4547 -5519
rect 4606 -5538 4649 -5504
rect 4599 -5571 4649 -5538
rect 3683 -5697 4649 -5571
rect 3683 -5749 3737 -5697
rect 3789 -5749 3801 -5697
rect 3853 -5749 3865 -5697
rect 3917 -5749 3933 -5697
rect 3985 -5749 3997 -5697
rect 4049 -5749 4061 -5697
rect 4113 -5749 4223 -5697
rect 4275 -5749 4287 -5697
rect 4339 -5749 4351 -5697
rect 4403 -5749 4419 -5697
rect 4471 -5749 4483 -5697
rect 4535 -5749 4547 -5697
rect 4599 -5749 4649 -5697
rect 3683 -5768 4649 -5749
rect 4853 -5503 5643 -5465
rect 9210 -5465 9589 -5431
rect 9623 -5465 9646 -5431
rect 4853 -5504 5231 -5503
rect 4853 -5538 4952 -5504
rect 4986 -5538 5024 -5504
rect 5058 -5537 5231 -5504
rect 5265 -5504 5643 -5503
rect 5265 -5537 5438 -5504
rect 5058 -5538 5438 -5537
rect 5472 -5538 5510 -5504
rect 5544 -5538 5643 -5504
rect 4853 -5575 5643 -5538
rect 4853 -5609 5231 -5575
rect 5265 -5609 5643 -5575
rect 4853 -5647 5643 -5609
rect 4853 -5681 5231 -5647
rect 5265 -5681 5643 -5647
rect 4853 -5719 5643 -5681
rect 4853 -5753 5231 -5719
rect 5265 -5753 5643 -5719
rect 4853 -5791 5643 -5753
rect 5846 -5504 6812 -5498
rect 5846 -5538 5889 -5504
rect 5923 -5519 5961 -5504
rect 5995 -5519 6147 -5504
rect 6181 -5519 6219 -5504
rect 6253 -5519 6405 -5504
rect 6439 -5519 6477 -5504
rect 6511 -5519 6663 -5504
rect 6697 -5519 6735 -5504
rect 5846 -5571 5896 -5538
rect 5948 -5571 5960 -5519
rect 6012 -5571 6024 -5519
rect 6076 -5571 6092 -5519
rect 6144 -5538 6147 -5519
rect 6208 -5538 6219 -5519
rect 6144 -5571 6156 -5538
rect 6208 -5571 6220 -5538
rect 6272 -5571 6382 -5519
rect 6439 -5538 6446 -5519
rect 6434 -5571 6446 -5538
rect 6498 -5571 6510 -5538
rect 6562 -5571 6578 -5519
rect 6630 -5571 6642 -5519
rect 6697 -5538 6706 -5519
rect 6769 -5538 6812 -5504
rect 6694 -5571 6706 -5538
rect 6758 -5571 6812 -5538
rect 5846 -5697 6812 -5571
rect 5846 -5749 5896 -5697
rect 5948 -5749 5960 -5697
rect 6012 -5749 6024 -5697
rect 6076 -5749 6092 -5697
rect 6144 -5749 6156 -5697
rect 6208 -5749 6220 -5697
rect 6272 -5749 6382 -5697
rect 6434 -5749 6446 -5697
rect 6498 -5749 6510 -5697
rect 6562 -5749 6578 -5697
rect 6630 -5749 6642 -5697
rect 6694 -5749 6706 -5697
rect 6758 -5749 6812 -5697
rect 5846 -5768 6812 -5749
rect 6889 -5504 7963 -5498
rect 6889 -5538 7115 -5504
rect 7149 -5538 7187 -5504
rect 7221 -5538 7373 -5504
rect 7407 -5538 7445 -5504
rect 7479 -5538 7631 -5504
rect 7665 -5538 7703 -5504
rect 7737 -5538 7963 -5504
rect 6889 -5586 7963 -5538
rect 3545 -5836 4649 -5818
rect 3545 -5866 3737 -5836
rect 3789 -5866 3801 -5836
rect 3545 -5900 3726 -5866
rect 3789 -5888 3798 -5866
rect 3853 -5888 3865 -5836
rect 3917 -5888 3933 -5836
rect 3985 -5866 3997 -5836
rect 4049 -5866 4061 -5836
rect 4049 -5888 4056 -5866
rect 4113 -5888 4223 -5836
rect 4275 -5866 4287 -5836
rect 4339 -5866 4351 -5836
rect 4276 -5888 4287 -5866
rect 4348 -5888 4351 -5866
rect 4403 -5888 4419 -5836
rect 4471 -5888 4483 -5836
rect 4535 -5888 4547 -5836
rect 4599 -5866 4649 -5836
rect 3760 -5900 3798 -5888
rect 3832 -5900 3984 -5888
rect 4018 -5900 4056 -5888
rect 4090 -5900 4242 -5888
rect 4276 -5900 4314 -5888
rect 4348 -5900 4500 -5888
rect 4534 -5900 4572 -5888
rect 4606 -5900 4649 -5866
rect 3545 -5906 4649 -5900
rect 4853 -5825 5231 -5791
rect 5265 -5825 5643 -5791
rect 6889 -5818 6950 -5586
rect 4853 -5863 5643 -5825
rect 4853 -5866 5231 -5863
rect 4853 -5900 4952 -5866
rect 4986 -5900 5024 -5866
rect 5058 -5897 5231 -5866
rect 5265 -5866 5643 -5863
rect 5265 -5897 5438 -5866
rect 5058 -5900 5438 -5897
rect 5472 -5900 5510 -5866
rect 5544 -5900 5643 -5866
rect 849 -5969 872 -5935
rect 906 -5969 1285 -5935
rect 4853 -5935 5643 -5900
rect 5846 -5836 6950 -5818
rect 5846 -5866 5896 -5836
rect 5846 -5900 5889 -5866
rect 5948 -5888 5960 -5836
rect 6012 -5888 6024 -5836
rect 6076 -5888 6092 -5836
rect 6144 -5866 6156 -5836
rect 6208 -5866 6220 -5836
rect 6144 -5888 6147 -5866
rect 6208 -5888 6219 -5866
rect 6272 -5888 6382 -5836
rect 6434 -5866 6446 -5836
rect 6498 -5866 6510 -5836
rect 6439 -5888 6446 -5866
rect 6562 -5888 6578 -5836
rect 6630 -5888 6642 -5836
rect 6694 -5866 6706 -5836
rect 6758 -5866 6950 -5836
rect 6697 -5888 6706 -5866
rect 5923 -5900 5961 -5888
rect 5995 -5900 6147 -5888
rect 6181 -5900 6219 -5888
rect 6253 -5900 6405 -5888
rect 6439 -5900 6477 -5888
rect 6511 -5900 6663 -5888
rect 6697 -5900 6735 -5888
rect 6769 -5900 6950 -5866
rect 5846 -5906 6950 -5900
rect 7072 -5697 7780 -5680
rect 7072 -5749 7110 -5697
rect 7162 -5749 7174 -5697
rect 7226 -5749 7238 -5697
rect 7290 -5749 7306 -5697
rect 7358 -5749 7370 -5697
rect 7422 -5749 7434 -5697
rect 7486 -5749 7498 -5697
rect 7550 -5749 7566 -5697
rect 7618 -5749 7630 -5697
rect 7682 -5749 7694 -5697
rect 7746 -5749 7780 -5697
rect 7072 -5866 7780 -5749
rect 7072 -5900 7115 -5866
rect 7149 -5900 7187 -5866
rect 7221 -5900 7373 -5866
rect 7407 -5900 7445 -5866
rect 7479 -5900 7631 -5866
rect 7665 -5900 7703 -5866
rect 7737 -5900 7780 -5866
rect 7072 -5906 7780 -5900
rect 7902 -5818 7963 -5586
rect 8040 -5504 9006 -5498
rect 8040 -5538 8083 -5504
rect 8117 -5519 8155 -5504
rect 8189 -5519 8341 -5504
rect 8375 -5519 8413 -5504
rect 8447 -5519 8599 -5504
rect 8633 -5519 8671 -5504
rect 8705 -5519 8857 -5504
rect 8891 -5519 8929 -5504
rect 8146 -5538 8155 -5519
rect 8040 -5571 8094 -5538
rect 8146 -5571 8158 -5538
rect 8210 -5571 8222 -5519
rect 8274 -5571 8290 -5519
rect 8406 -5538 8413 -5519
rect 8342 -5571 8354 -5538
rect 8406 -5571 8418 -5538
rect 8470 -5571 8580 -5519
rect 8633 -5538 8644 -5519
rect 8705 -5538 8708 -5519
rect 8632 -5571 8644 -5538
rect 8696 -5571 8708 -5538
rect 8760 -5571 8776 -5519
rect 8828 -5571 8840 -5519
rect 8892 -5571 8904 -5519
rect 8963 -5538 9006 -5504
rect 8956 -5571 9006 -5538
rect 8040 -5697 9006 -5571
rect 8040 -5749 8094 -5697
rect 8146 -5749 8158 -5697
rect 8210 -5749 8222 -5697
rect 8274 -5749 8290 -5697
rect 8342 -5749 8354 -5697
rect 8406 -5749 8418 -5697
rect 8470 -5749 8580 -5697
rect 8632 -5749 8644 -5697
rect 8696 -5749 8708 -5697
rect 8760 -5749 8776 -5697
rect 8828 -5749 8840 -5697
rect 8892 -5749 8904 -5697
rect 8956 -5749 9006 -5697
rect 8040 -5768 9006 -5749
rect 9210 -5503 9646 -5465
rect 9210 -5504 9589 -5503
rect 9210 -5538 9309 -5504
rect 9343 -5538 9381 -5504
rect 9415 -5537 9589 -5504
rect 9623 -5537 9646 -5503
rect 9415 -5538 9646 -5537
rect 9210 -5575 9646 -5538
rect 9210 -5609 9589 -5575
rect 9623 -5609 9646 -5575
rect 9210 -5647 9646 -5609
rect 9210 -5681 9589 -5647
rect 9623 -5681 9646 -5647
rect 9210 -5719 9646 -5681
rect 9210 -5753 9589 -5719
rect 9623 -5753 9646 -5719
rect 9210 -5791 9646 -5753
rect 7902 -5836 9006 -5818
rect 7902 -5866 8094 -5836
rect 8146 -5866 8158 -5836
rect 7902 -5900 8083 -5866
rect 8146 -5888 8155 -5866
rect 8210 -5888 8222 -5836
rect 8274 -5888 8290 -5836
rect 8342 -5866 8354 -5836
rect 8406 -5866 8418 -5836
rect 8406 -5888 8413 -5866
rect 8470 -5888 8580 -5836
rect 8632 -5866 8644 -5836
rect 8696 -5866 8708 -5836
rect 8633 -5888 8644 -5866
rect 8705 -5888 8708 -5866
rect 8760 -5888 8776 -5836
rect 8828 -5888 8840 -5836
rect 8892 -5888 8904 -5836
rect 8956 -5866 9006 -5836
rect 8117 -5900 8155 -5888
rect 8189 -5900 8341 -5888
rect 8375 -5900 8413 -5888
rect 8447 -5900 8599 -5888
rect 8633 -5900 8671 -5888
rect 8705 -5900 8857 -5888
rect 8891 -5900 8929 -5888
rect 8963 -5900 9006 -5866
rect 7902 -5906 9006 -5900
rect 9210 -5825 9589 -5791
rect 9623 -5825 9646 -5791
rect 9210 -5863 9646 -5825
rect 9210 -5866 9589 -5863
rect 9210 -5900 9309 -5866
rect 9343 -5900 9381 -5866
rect 9415 -5897 9589 -5866
rect 9623 -5897 9646 -5863
rect 9415 -5900 9646 -5897
rect 849 -5994 1285 -5969
rect 849 -6007 987 -5994
rect 849 -6041 872 -6007
rect 906 -6028 987 -6007
rect 1021 -6028 1245 -5994
rect 1279 -6028 1285 -5994
rect 906 -6041 1285 -6028
rect 849 -6066 1285 -6041
rect 849 -6079 987 -6066
rect 849 -6113 872 -6079
rect 906 -6100 987 -6079
rect 1021 -6100 1245 -6066
rect 1279 -6100 1285 -6066
rect 906 -6113 1285 -6100
rect 849 -6151 1285 -6113
rect 849 -6185 872 -6151
rect 906 -6185 1285 -6151
rect 849 -6223 1285 -6185
rect 849 -6257 872 -6223
rect 906 -6257 1285 -6223
rect 849 -6295 1285 -6257
rect 849 -6329 872 -6295
rect 906 -6329 1285 -6295
rect 849 -6367 1285 -6329
rect 849 -6401 872 -6367
rect 906 -6401 1285 -6367
rect 849 -6439 1285 -6401
rect 849 -6473 872 -6439
rect 906 -6473 1285 -6439
rect 849 -6511 1285 -6473
rect 849 -6545 872 -6511
rect 906 -6545 1285 -6511
rect 849 -6583 1285 -6545
rect 849 -6617 872 -6583
rect 906 -6617 1285 -6583
rect 849 -6655 1285 -6617
rect 849 -6689 872 -6655
rect 906 -6689 1285 -6655
rect 849 -6727 1285 -6689
rect 1433 -5994 1479 -5947
rect 1433 -6028 1439 -5994
rect 1473 -6028 1479 -5994
rect 1433 -6066 1479 -6028
rect 1433 -6100 1439 -6066
rect 1473 -6100 1479 -6066
rect 1433 -6707 1479 -6100
rect 1691 -5994 1737 -5947
rect 1691 -6028 1697 -5994
rect 1731 -6028 1737 -5994
rect 1691 -6066 1737 -6028
rect 1691 -6100 1697 -6066
rect 1731 -6100 1737 -6066
rect 1691 -6406 1737 -6100
rect 1949 -5994 1995 -5947
rect 1949 -6028 1955 -5994
rect 1989 -6028 1995 -5994
rect 1949 -6066 1995 -6028
rect 1949 -6100 1955 -6066
rect 1989 -6100 1995 -6066
rect 1618 -6416 1814 -6406
rect 1618 -6468 1625 -6416
rect 1677 -6468 1689 -6416
rect 1741 -6468 1753 -6416
rect 1805 -6468 1814 -6416
rect 1618 -6476 1814 -6468
rect 849 -6761 872 -6727
rect 906 -6761 1285 -6727
rect 849 -6799 1285 -6761
rect 1360 -6717 1556 -6707
rect 1360 -6769 1367 -6717
rect 1419 -6769 1431 -6717
rect 1483 -6769 1495 -6717
rect 1547 -6769 1556 -6717
rect 1360 -6777 1556 -6769
rect 849 -6833 872 -6799
rect 906 -6833 1285 -6799
rect 849 -6871 1285 -6833
rect 849 -6905 872 -6871
rect 906 -6905 1285 -6871
rect 849 -6943 1285 -6905
rect 849 -6977 872 -6943
rect 906 -6951 1285 -6943
rect 906 -6977 987 -6951
rect 849 -6985 987 -6977
rect 1021 -6985 1245 -6951
rect 1279 -6985 1285 -6951
rect 849 -7015 1285 -6985
rect 849 -7049 872 -7015
rect 906 -7023 1285 -7015
rect 906 -7049 987 -7023
rect 849 -7057 987 -7049
rect 1021 -7057 1245 -7023
rect 1279 -7057 1285 -7023
rect 849 -7087 1285 -7057
rect 849 -7121 872 -7087
rect 906 -7121 1285 -7087
rect 1433 -6951 1479 -6777
rect 1433 -6985 1439 -6951
rect 1473 -6985 1479 -6951
rect 1433 -7023 1479 -6985
rect 1433 -7057 1439 -7023
rect 1473 -7057 1479 -7023
rect 1433 -7104 1479 -7057
rect 1691 -6951 1737 -6476
rect 1949 -6707 1995 -6100
rect 2207 -5994 2253 -5947
rect 2207 -6028 2213 -5994
rect 2247 -6028 2253 -5994
rect 2207 -6066 2253 -6028
rect 2207 -6100 2213 -6066
rect 2247 -6100 2253 -6066
rect 2207 -6406 2253 -6100
rect 2465 -5994 2511 -5947
rect 2465 -6028 2471 -5994
rect 2505 -6028 2511 -5994
rect 2465 -6066 2511 -6028
rect 2465 -6100 2471 -6066
rect 2505 -6100 2511 -6066
rect 2135 -6416 2331 -6406
rect 2135 -6468 2142 -6416
rect 2194 -6468 2206 -6416
rect 2258 -6468 2270 -6416
rect 2322 -6468 2331 -6416
rect 2135 -6476 2331 -6468
rect 1875 -6717 2071 -6707
rect 1875 -6769 1882 -6717
rect 1934 -6769 1946 -6717
rect 1998 -6769 2010 -6717
rect 2062 -6769 2071 -6717
rect 1875 -6777 2071 -6769
rect 1691 -6985 1697 -6951
rect 1731 -6985 1737 -6951
rect 1691 -7023 1737 -6985
rect 1691 -7057 1697 -7023
rect 1731 -7057 1737 -7023
rect 1691 -7104 1737 -7057
rect 1949 -6951 1995 -6777
rect 1949 -6985 1955 -6951
rect 1989 -6985 1995 -6951
rect 1949 -7023 1995 -6985
rect 1949 -7057 1955 -7023
rect 1989 -7057 1995 -7023
rect 1949 -7104 1995 -7057
rect 2207 -6951 2253 -6476
rect 2465 -6707 2511 -6100
rect 2659 -5994 2705 -5947
rect 2659 -6028 2665 -5994
rect 2699 -6028 2705 -5994
rect 2659 -6066 2705 -6028
rect 2659 -6100 2665 -6066
rect 2699 -6100 2705 -6066
rect 2659 -6261 2705 -6100
rect 2917 -5994 2963 -5947
rect 2917 -6028 2923 -5994
rect 2957 -6028 2963 -5994
rect 2917 -6066 2963 -6028
rect 2917 -6100 2923 -6066
rect 2957 -6100 2963 -6066
rect 2582 -6271 2778 -6261
rect 2582 -6323 2591 -6271
rect 2643 -6323 2655 -6271
rect 2707 -6323 2719 -6271
rect 2771 -6323 2778 -6271
rect 2582 -6331 2778 -6323
rect 2392 -6717 2588 -6707
rect 2392 -6769 2399 -6717
rect 2451 -6769 2463 -6717
rect 2515 -6769 2527 -6717
rect 2579 -6769 2588 -6717
rect 2392 -6777 2588 -6769
rect 2207 -6985 2213 -6951
rect 2247 -6985 2253 -6951
rect 2207 -7023 2253 -6985
rect 2207 -7057 2213 -7023
rect 2247 -7057 2253 -7023
rect 2207 -7104 2253 -7057
rect 2465 -6951 2511 -6777
rect 2465 -6985 2471 -6951
rect 2505 -6985 2511 -6951
rect 2465 -7023 2511 -6985
rect 2465 -7057 2471 -7023
rect 2505 -7057 2511 -7023
rect 2465 -7104 2511 -7057
rect 2659 -6951 2705 -6331
rect 2917 -6567 2963 -6100
rect 3175 -5994 3221 -5947
rect 3175 -6028 3181 -5994
rect 3215 -6028 3221 -5994
rect 3175 -6066 3221 -6028
rect 3175 -6100 3181 -6066
rect 3215 -6100 3221 -6066
rect 3175 -6261 3221 -6100
rect 3433 -5994 3479 -5947
rect 3433 -6028 3439 -5994
rect 3473 -6028 3479 -5994
rect 3433 -6066 3479 -6028
rect 3433 -6100 3439 -6066
rect 3473 -6100 3479 -6066
rect 3099 -6271 3295 -6261
rect 3099 -6323 3108 -6271
rect 3160 -6323 3172 -6271
rect 3224 -6323 3236 -6271
rect 3288 -6323 3295 -6271
rect 3099 -6331 3295 -6323
rect 2840 -6577 3036 -6567
rect 2840 -6629 2849 -6577
rect 2901 -6629 2913 -6577
rect 2965 -6629 2977 -6577
rect 3029 -6629 3036 -6577
rect 2840 -6637 3036 -6629
rect 2659 -6985 2665 -6951
rect 2699 -6985 2705 -6951
rect 2659 -7023 2705 -6985
rect 2659 -7057 2665 -7023
rect 2699 -7057 2705 -7023
rect 2659 -7104 2705 -7057
rect 2917 -6951 2963 -6637
rect 2917 -6985 2923 -6951
rect 2957 -6985 2963 -6951
rect 2917 -7023 2963 -6985
rect 2917 -7057 2923 -7023
rect 2957 -7057 2963 -7023
rect 2917 -7104 2963 -7057
rect 3175 -6951 3221 -6331
rect 3433 -6567 3479 -6100
rect 3627 -5994 3673 -5947
rect 3627 -6028 3633 -5994
rect 3667 -6028 3673 -5994
rect 3627 -6066 3673 -6028
rect 3627 -6100 3633 -6066
rect 3667 -6100 3673 -6066
rect 3357 -6577 3553 -6567
rect 3357 -6629 3366 -6577
rect 3418 -6629 3430 -6577
rect 3482 -6629 3494 -6577
rect 3546 -6629 3553 -6577
rect 3357 -6637 3553 -6629
rect 3175 -6985 3181 -6951
rect 3215 -6985 3221 -6951
rect 3175 -7023 3221 -6985
rect 3175 -7057 3181 -7023
rect 3215 -7057 3221 -7023
rect 3175 -7104 3221 -7057
rect 3433 -6951 3479 -6637
rect 3627 -6707 3673 -6100
rect 3885 -5994 3931 -5947
rect 3885 -6028 3891 -5994
rect 3925 -6028 3931 -5994
rect 3885 -6066 3931 -6028
rect 3885 -6100 3891 -6066
rect 3925 -6100 3931 -6066
rect 3885 -6406 3931 -6100
rect 4143 -5994 4189 -5947
rect 4143 -6028 4149 -5994
rect 4183 -6028 4189 -5994
rect 4143 -6066 4189 -6028
rect 4143 -6100 4149 -6066
rect 4183 -6100 4189 -6066
rect 3812 -6416 4008 -6406
rect 3812 -6468 3819 -6416
rect 3871 -6468 3883 -6416
rect 3935 -6468 3947 -6416
rect 3999 -6468 4008 -6416
rect 3812 -6476 4008 -6468
rect 3552 -6717 3748 -6707
rect 3552 -6769 3559 -6717
rect 3611 -6769 3623 -6717
rect 3675 -6769 3687 -6717
rect 3739 -6769 3748 -6717
rect 3552 -6777 3748 -6769
rect 3433 -6985 3439 -6951
rect 3473 -6985 3479 -6951
rect 3433 -7023 3479 -6985
rect 3433 -7057 3439 -7023
rect 3473 -7057 3479 -7023
rect 3433 -7104 3479 -7057
rect 3627 -6951 3673 -6777
rect 3627 -6985 3633 -6951
rect 3667 -6985 3673 -6951
rect 3627 -7023 3673 -6985
rect 3627 -7057 3633 -7023
rect 3667 -7057 3673 -7023
rect 3627 -7104 3673 -7057
rect 3885 -6951 3931 -6476
rect 4143 -6707 4189 -6100
rect 4401 -5994 4447 -5947
rect 4401 -6028 4407 -5994
rect 4441 -6028 4447 -5994
rect 4401 -6066 4447 -6028
rect 4401 -6100 4407 -6066
rect 4441 -6100 4447 -6066
rect 4401 -6406 4447 -6100
rect 4659 -5994 4705 -5947
rect 4659 -6028 4665 -5994
rect 4699 -6028 4705 -5994
rect 4659 -6066 4705 -6028
rect 4659 -6100 4665 -6066
rect 4699 -6100 4705 -6066
rect 4329 -6416 4525 -6406
rect 4329 -6468 4336 -6416
rect 4388 -6468 4400 -6416
rect 4452 -6468 4464 -6416
rect 4516 -6468 4525 -6416
rect 4329 -6476 4525 -6468
rect 4069 -6717 4265 -6707
rect 4069 -6769 4076 -6717
rect 4128 -6769 4140 -6717
rect 4192 -6769 4204 -6717
rect 4256 -6769 4265 -6717
rect 4069 -6777 4265 -6769
rect 3885 -6985 3891 -6951
rect 3925 -6985 3931 -6951
rect 3885 -7023 3931 -6985
rect 3885 -7057 3891 -7023
rect 3925 -7057 3931 -7023
rect 3885 -7104 3931 -7057
rect 4143 -6951 4189 -6777
rect 4143 -6985 4149 -6951
rect 4183 -6985 4189 -6951
rect 4143 -7023 4189 -6985
rect 4143 -7057 4149 -7023
rect 4183 -7057 4189 -7023
rect 4143 -7104 4189 -7057
rect 4401 -6951 4447 -6476
rect 4659 -6707 4705 -6100
rect 4853 -5969 5231 -5935
rect 5265 -5969 5643 -5935
rect 9210 -5935 9646 -5900
rect 4853 -5994 5643 -5969
rect 4853 -6028 4859 -5994
rect 4893 -6028 5117 -5994
rect 5151 -6007 5345 -5994
rect 5151 -6028 5231 -6007
rect 4853 -6041 5231 -6028
rect 5265 -6028 5345 -6007
rect 5379 -6028 5603 -5994
rect 5637 -6028 5643 -5994
rect 5265 -6041 5643 -6028
rect 4853 -6066 5643 -6041
rect 4853 -6100 4859 -6066
rect 4893 -6100 5117 -6066
rect 5151 -6079 5345 -6066
rect 5151 -6100 5231 -6079
rect 4853 -6113 5231 -6100
rect 5265 -6100 5345 -6079
rect 5379 -6100 5603 -6066
rect 5637 -6100 5643 -6066
rect 5265 -6113 5643 -6100
rect 4853 -6151 5643 -6113
rect 4853 -6185 5231 -6151
rect 5265 -6185 5643 -6151
rect 4853 -6223 5643 -6185
rect 4853 -6257 5231 -6223
rect 5265 -6257 5643 -6223
rect 4853 -6295 5643 -6257
rect 4853 -6329 5231 -6295
rect 5265 -6329 5643 -6295
rect 4853 -6367 5643 -6329
rect 4853 -6401 5231 -6367
rect 5265 -6401 5643 -6367
rect 4853 -6439 5643 -6401
rect 4853 -6473 5231 -6439
rect 5265 -6473 5643 -6439
rect 4853 -6511 5643 -6473
rect 4853 -6545 5231 -6511
rect 5265 -6545 5643 -6511
rect 4853 -6583 5643 -6545
rect 4853 -6617 5231 -6583
rect 5265 -6617 5643 -6583
rect 4853 -6655 5643 -6617
rect 4853 -6689 5231 -6655
rect 5265 -6689 5643 -6655
rect 4586 -6717 4782 -6707
rect 4586 -6769 4593 -6717
rect 4645 -6769 4657 -6717
rect 4709 -6769 4721 -6717
rect 4773 -6769 4782 -6717
rect 4586 -6777 4782 -6769
rect 4853 -6727 5643 -6689
rect 5790 -5994 5836 -5947
rect 5790 -6028 5796 -5994
rect 5830 -6028 5836 -5994
rect 5790 -6066 5836 -6028
rect 5790 -6100 5796 -6066
rect 5830 -6100 5836 -6066
rect 5790 -6707 5836 -6100
rect 6048 -5994 6094 -5947
rect 6048 -6028 6054 -5994
rect 6088 -6028 6094 -5994
rect 6048 -6066 6094 -6028
rect 6048 -6100 6054 -6066
rect 6088 -6100 6094 -6066
rect 6048 -6406 6094 -6100
rect 6306 -5994 6352 -5947
rect 6306 -6028 6312 -5994
rect 6346 -6028 6352 -5994
rect 6306 -6066 6352 -6028
rect 6306 -6100 6312 -6066
rect 6346 -6100 6352 -6066
rect 5970 -6416 6166 -6406
rect 5970 -6468 5979 -6416
rect 6031 -6468 6043 -6416
rect 6095 -6468 6107 -6416
rect 6159 -6468 6166 -6416
rect 5970 -6476 6166 -6468
rect 4853 -6761 5231 -6727
rect 5265 -6761 5643 -6727
rect 4401 -6985 4407 -6951
rect 4441 -6985 4447 -6951
rect 4401 -7023 4447 -6985
rect 4401 -7057 4407 -7023
rect 4441 -7057 4447 -7023
rect 4401 -7104 4447 -7057
rect 4659 -6951 4705 -6777
rect 4659 -6985 4665 -6951
rect 4699 -6985 4705 -6951
rect 4659 -7023 4705 -6985
rect 4659 -7057 4665 -7023
rect 4699 -7057 4705 -7023
rect 4659 -7104 4705 -7057
rect 4853 -6799 5643 -6761
rect 5713 -6717 5909 -6707
rect 5713 -6769 5722 -6717
rect 5774 -6769 5786 -6717
rect 5838 -6769 5850 -6717
rect 5902 -6769 5909 -6717
rect 5713 -6777 5909 -6769
rect 4853 -6833 5231 -6799
rect 5265 -6833 5643 -6799
rect 4853 -6871 5643 -6833
rect 4853 -6905 5231 -6871
rect 5265 -6905 5643 -6871
rect 4853 -6943 5643 -6905
rect 4853 -6951 5231 -6943
rect 4853 -6985 4859 -6951
rect 4893 -6985 5117 -6951
rect 5151 -6977 5231 -6951
rect 5265 -6951 5643 -6943
rect 5265 -6977 5345 -6951
rect 5151 -6985 5345 -6977
rect 5379 -6985 5603 -6951
rect 5637 -6985 5643 -6951
rect 4853 -7015 5643 -6985
rect 4853 -7023 5231 -7015
rect 4853 -7057 4859 -7023
rect 4893 -7057 5117 -7023
rect 5151 -7049 5231 -7023
rect 5265 -7023 5643 -7015
rect 5265 -7049 5345 -7023
rect 5151 -7057 5345 -7049
rect 5379 -7057 5603 -7023
rect 5637 -7057 5643 -7023
rect 4853 -7087 5643 -7057
rect 849 -7151 1285 -7121
rect 4853 -7121 5231 -7087
rect 5265 -7121 5643 -7087
rect 5790 -6951 5836 -6777
rect 5790 -6985 5796 -6951
rect 5830 -6985 5836 -6951
rect 5790 -7023 5836 -6985
rect 5790 -7057 5796 -7023
rect 5830 -7057 5836 -7023
rect 5790 -7104 5836 -7057
rect 6048 -6951 6094 -6476
rect 6306 -6707 6352 -6100
rect 6564 -5994 6610 -5947
rect 6564 -6028 6570 -5994
rect 6604 -6028 6610 -5994
rect 6564 -6066 6610 -6028
rect 6564 -6100 6570 -6066
rect 6604 -6100 6610 -6066
rect 6564 -6406 6610 -6100
rect 6822 -5994 6868 -5947
rect 6822 -6028 6828 -5994
rect 6862 -6028 6868 -5994
rect 6822 -6066 6868 -6028
rect 6822 -6100 6828 -6066
rect 6862 -6100 6868 -6066
rect 6487 -6416 6683 -6406
rect 6487 -6468 6496 -6416
rect 6548 -6468 6560 -6416
rect 6612 -6468 6624 -6416
rect 6676 -6468 6683 -6416
rect 6487 -6476 6683 -6468
rect 6230 -6717 6426 -6707
rect 6230 -6769 6239 -6717
rect 6291 -6769 6303 -6717
rect 6355 -6769 6367 -6717
rect 6419 -6769 6426 -6717
rect 6230 -6777 6426 -6769
rect 6048 -6985 6054 -6951
rect 6088 -6985 6094 -6951
rect 6048 -7023 6094 -6985
rect 6048 -7057 6054 -7023
rect 6088 -7057 6094 -7023
rect 6048 -7104 6094 -7057
rect 6306 -6951 6352 -6777
rect 6306 -6985 6312 -6951
rect 6346 -6985 6352 -6951
rect 6306 -7023 6352 -6985
rect 6306 -7057 6312 -7023
rect 6346 -7057 6352 -7023
rect 6306 -7104 6352 -7057
rect 6564 -6951 6610 -6476
rect 6822 -6707 6868 -6100
rect 7016 -5994 7062 -5947
rect 7016 -6028 7022 -5994
rect 7056 -6028 7062 -5994
rect 7016 -6066 7062 -6028
rect 7016 -6100 7022 -6066
rect 7056 -6100 7062 -6066
rect 7016 -6567 7062 -6100
rect 7274 -5994 7320 -5947
rect 7274 -6028 7280 -5994
rect 7314 -6028 7320 -5994
rect 7274 -6066 7320 -6028
rect 7274 -6100 7280 -6066
rect 7314 -6100 7320 -6066
rect 7274 -6261 7320 -6100
rect 7532 -5994 7578 -5947
rect 7532 -6028 7538 -5994
rect 7572 -6028 7578 -5994
rect 7532 -6066 7578 -6028
rect 7532 -6100 7538 -6066
rect 7572 -6100 7578 -6066
rect 7200 -6271 7396 -6261
rect 7200 -6323 7207 -6271
rect 7259 -6323 7271 -6271
rect 7323 -6323 7335 -6271
rect 7387 -6323 7396 -6271
rect 7200 -6331 7396 -6323
rect 6942 -6577 7138 -6567
rect 6942 -6629 6949 -6577
rect 7001 -6629 7013 -6577
rect 7065 -6629 7077 -6577
rect 7129 -6629 7138 -6577
rect 6942 -6637 7138 -6629
rect 6747 -6717 6943 -6707
rect 6747 -6769 6756 -6717
rect 6808 -6769 6820 -6717
rect 6872 -6769 6884 -6717
rect 6936 -6769 6943 -6717
rect 6747 -6777 6943 -6769
rect 6564 -6985 6570 -6951
rect 6604 -6985 6610 -6951
rect 6564 -7023 6610 -6985
rect 6564 -7057 6570 -7023
rect 6604 -7057 6610 -7023
rect 6564 -7104 6610 -7057
rect 6822 -6951 6868 -6777
rect 6822 -6985 6828 -6951
rect 6862 -6985 6868 -6951
rect 6822 -7023 6868 -6985
rect 6822 -7057 6828 -7023
rect 6862 -7057 6868 -7023
rect 6822 -7104 6868 -7057
rect 7016 -6951 7062 -6637
rect 7016 -6985 7022 -6951
rect 7056 -6985 7062 -6951
rect 7016 -7023 7062 -6985
rect 7016 -7057 7022 -7023
rect 7056 -7057 7062 -7023
rect 7016 -7104 7062 -7057
rect 7274 -6951 7320 -6331
rect 7532 -6567 7578 -6100
rect 7790 -5994 7836 -5947
rect 7790 -6028 7796 -5994
rect 7830 -6028 7836 -5994
rect 7790 -6066 7836 -6028
rect 7790 -6100 7796 -6066
rect 7830 -6100 7836 -6066
rect 7790 -6261 7836 -6100
rect 7984 -5994 8030 -5947
rect 7984 -6028 7990 -5994
rect 8024 -6028 8030 -5994
rect 7984 -6066 8030 -6028
rect 7984 -6100 7990 -6066
rect 8024 -6100 8030 -6066
rect 7717 -6271 7913 -6261
rect 7717 -6323 7724 -6271
rect 7776 -6323 7788 -6271
rect 7840 -6323 7852 -6271
rect 7904 -6323 7913 -6271
rect 7717 -6331 7913 -6323
rect 7459 -6577 7655 -6567
rect 7459 -6629 7466 -6577
rect 7518 -6629 7530 -6577
rect 7582 -6629 7594 -6577
rect 7646 -6629 7655 -6577
rect 7459 -6637 7655 -6629
rect 7274 -6985 7280 -6951
rect 7314 -6985 7320 -6951
rect 7274 -7023 7320 -6985
rect 7274 -7057 7280 -7023
rect 7314 -7057 7320 -7023
rect 7274 -7104 7320 -7057
rect 7532 -6951 7578 -6637
rect 7532 -6985 7538 -6951
rect 7572 -6985 7578 -6951
rect 7532 -7023 7578 -6985
rect 7532 -7057 7538 -7023
rect 7572 -7057 7578 -7023
rect 7532 -7104 7578 -7057
rect 7790 -6951 7836 -6331
rect 7984 -6707 8030 -6100
rect 8242 -5994 8288 -5947
rect 8242 -6028 8248 -5994
rect 8282 -6028 8288 -5994
rect 8242 -6066 8288 -6028
rect 8242 -6100 8248 -6066
rect 8282 -6100 8288 -6066
rect 8242 -6406 8288 -6100
rect 8500 -5994 8546 -5947
rect 8500 -6028 8506 -5994
rect 8540 -6028 8546 -5994
rect 8500 -6066 8546 -6028
rect 8500 -6100 8506 -6066
rect 8540 -6100 8546 -6066
rect 8164 -6416 8360 -6406
rect 8164 -6468 8173 -6416
rect 8225 -6468 8237 -6416
rect 8289 -6468 8301 -6416
rect 8353 -6468 8360 -6416
rect 8164 -6476 8360 -6468
rect 7907 -6717 8103 -6707
rect 7907 -6769 7916 -6717
rect 7968 -6769 7980 -6717
rect 8032 -6769 8044 -6717
rect 8096 -6769 8103 -6717
rect 7907 -6777 8103 -6769
rect 7790 -6985 7796 -6951
rect 7830 -6985 7836 -6951
rect 7790 -7023 7836 -6985
rect 7790 -7057 7796 -7023
rect 7830 -7057 7836 -7023
rect 7790 -7104 7836 -7057
rect 7984 -6951 8030 -6777
rect 7984 -6985 7990 -6951
rect 8024 -6985 8030 -6951
rect 7984 -7023 8030 -6985
rect 7984 -7057 7990 -7023
rect 8024 -7057 8030 -7023
rect 7984 -7104 8030 -7057
rect 8242 -6951 8288 -6476
rect 8500 -6707 8546 -6100
rect 8758 -5994 8804 -5947
rect 8758 -6028 8764 -5994
rect 8798 -6028 8804 -5994
rect 8758 -6066 8804 -6028
rect 8758 -6100 8764 -6066
rect 8798 -6100 8804 -6066
rect 8758 -6406 8804 -6100
rect 9016 -5994 9062 -5947
rect 9016 -6028 9022 -5994
rect 9056 -6028 9062 -5994
rect 9016 -6066 9062 -6028
rect 9016 -6100 9022 -6066
rect 9056 -6100 9062 -6066
rect 8682 -6416 8878 -6406
rect 8682 -6468 8691 -6416
rect 8743 -6468 8755 -6416
rect 8807 -6468 8819 -6416
rect 8871 -6468 8878 -6416
rect 8682 -6476 8878 -6468
rect 8425 -6717 8621 -6707
rect 8425 -6769 8434 -6717
rect 8486 -6769 8498 -6717
rect 8550 -6769 8562 -6717
rect 8614 -6769 8621 -6717
rect 8425 -6777 8621 -6769
rect 8242 -6985 8248 -6951
rect 8282 -6985 8288 -6951
rect 8242 -7023 8288 -6985
rect 8242 -7057 8248 -7023
rect 8282 -7057 8288 -7023
rect 8242 -7104 8288 -7057
rect 8500 -6951 8546 -6777
rect 8500 -6985 8506 -6951
rect 8540 -6985 8546 -6951
rect 8500 -7023 8546 -6985
rect 8500 -7057 8506 -7023
rect 8540 -7057 8546 -7023
rect 8500 -7104 8546 -7057
rect 8758 -6951 8804 -6476
rect 9016 -6707 9062 -6100
rect 9210 -5969 9589 -5935
rect 9623 -5969 9646 -5935
rect 9210 -5994 9646 -5969
rect 9210 -6028 9216 -5994
rect 9250 -6028 9474 -5994
rect 9508 -6007 9646 -5994
rect 9508 -6028 9589 -6007
rect 9210 -6041 9589 -6028
rect 9623 -6041 9646 -6007
rect 9210 -6066 9646 -6041
rect 9210 -6100 9216 -6066
rect 9250 -6100 9474 -6066
rect 9508 -6079 9646 -6066
rect 9508 -6100 9589 -6079
rect 9210 -6113 9589 -6100
rect 9623 -6113 9646 -6079
rect 9210 -6151 9646 -6113
rect 9210 -6185 9589 -6151
rect 9623 -6185 9646 -6151
rect 9210 -6223 9646 -6185
rect 9210 -6257 9589 -6223
rect 9623 -6257 9646 -6223
rect 9210 -6295 9646 -6257
rect 9210 -6329 9589 -6295
rect 9623 -6329 9646 -6295
rect 9210 -6367 9646 -6329
rect 9210 -6401 9589 -6367
rect 9623 -6401 9646 -6367
rect 9210 -6439 9646 -6401
rect 9210 -6473 9589 -6439
rect 9623 -6473 9646 -6439
rect 9210 -6511 9646 -6473
rect 9210 -6545 9589 -6511
rect 9623 -6545 9646 -6511
rect 9210 -6583 9646 -6545
rect 9210 -6617 9589 -6583
rect 9623 -6617 9646 -6583
rect 9210 -6655 9646 -6617
rect 9210 -6689 9589 -6655
rect 9623 -6689 9646 -6655
rect 8940 -6717 9136 -6707
rect 8940 -6769 8949 -6717
rect 9001 -6769 9013 -6717
rect 9065 -6769 9077 -6717
rect 9129 -6769 9136 -6717
rect 8940 -6777 9136 -6769
rect 9210 -6727 9646 -6689
rect 9210 -6761 9589 -6727
rect 9623 -6761 9646 -6727
rect 8758 -6985 8764 -6951
rect 8798 -6985 8804 -6951
rect 8758 -7023 8804 -6985
rect 8758 -7057 8764 -7023
rect 8798 -7057 8804 -7023
rect 8758 -7104 8804 -7057
rect 9016 -6951 9062 -6777
rect 9016 -6985 9022 -6951
rect 9056 -6985 9062 -6951
rect 9016 -7023 9062 -6985
rect 9016 -7057 9022 -7023
rect 9056 -7057 9062 -7023
rect 9016 -7104 9062 -7057
rect 9210 -6799 9646 -6761
rect 9210 -6833 9589 -6799
rect 9623 -6833 9646 -6799
rect 9210 -6871 9646 -6833
rect 9210 -6905 9589 -6871
rect 9623 -6905 9646 -6871
rect 9210 -6943 9646 -6905
rect 9210 -6951 9589 -6943
rect 9210 -6985 9216 -6951
rect 9250 -6985 9474 -6951
rect 9508 -6977 9589 -6951
rect 9623 -6977 9646 -6943
rect 9508 -6985 9646 -6977
rect 9210 -7015 9646 -6985
rect 9210 -7023 9589 -7015
rect 9210 -7057 9216 -7023
rect 9250 -7057 9474 -7023
rect 9508 -7049 9589 -7023
rect 9623 -7049 9646 -7015
rect 9508 -7057 9646 -7049
rect 9210 -7087 9646 -7057
rect 849 -7159 1080 -7151
rect 849 -7193 872 -7159
rect 906 -7185 1080 -7159
rect 1114 -7185 1152 -7151
rect 1186 -7185 1285 -7151
rect 906 -7193 1285 -7185
rect 849 -7231 1285 -7193
rect 849 -7265 872 -7231
rect 906 -7265 1285 -7231
rect 849 -7303 1285 -7265
rect 849 -7337 872 -7303
rect 906 -7337 1285 -7303
rect 849 -7375 1285 -7337
rect 849 -7409 872 -7375
rect 906 -7409 1285 -7375
rect 849 -7447 1285 -7409
rect 1489 -7151 2455 -7145
rect 1489 -7185 1532 -7151
rect 1566 -7166 1604 -7151
rect 1638 -7166 1790 -7151
rect 1824 -7166 1862 -7151
rect 1896 -7166 2048 -7151
rect 2082 -7166 2120 -7151
rect 2154 -7166 2306 -7151
rect 2340 -7166 2378 -7151
rect 1489 -7218 1539 -7185
rect 1591 -7218 1603 -7166
rect 1655 -7218 1667 -7166
rect 1719 -7218 1735 -7166
rect 1787 -7185 1790 -7166
rect 1851 -7185 1862 -7166
rect 1787 -7218 1799 -7185
rect 1851 -7218 1863 -7185
rect 1915 -7218 2025 -7166
rect 2082 -7185 2089 -7166
rect 2077 -7218 2089 -7185
rect 2141 -7218 2153 -7185
rect 2205 -7218 2221 -7166
rect 2273 -7218 2285 -7166
rect 2340 -7185 2349 -7166
rect 2412 -7185 2455 -7151
rect 2337 -7218 2349 -7185
rect 2401 -7218 2455 -7185
rect 1489 -7344 2455 -7218
rect 1489 -7396 1539 -7344
rect 1591 -7396 1603 -7344
rect 1655 -7396 1667 -7344
rect 1719 -7396 1735 -7344
rect 1787 -7396 1799 -7344
rect 1851 -7396 1863 -7344
rect 1915 -7396 2025 -7344
rect 2077 -7396 2089 -7344
rect 2141 -7396 2153 -7344
rect 2205 -7396 2221 -7344
rect 2273 -7396 2285 -7344
rect 2337 -7396 2349 -7344
rect 2401 -7396 2455 -7344
rect 1489 -7415 2455 -7396
rect 2532 -7151 3606 -7145
rect 2532 -7185 2758 -7151
rect 2792 -7185 2830 -7151
rect 2864 -7185 3016 -7151
rect 3050 -7185 3088 -7151
rect 3122 -7185 3274 -7151
rect 3308 -7185 3346 -7151
rect 3380 -7185 3606 -7151
rect 2532 -7233 3606 -7185
rect 849 -7481 872 -7447
rect 906 -7481 1285 -7447
rect 2532 -7465 2593 -7233
rect 849 -7513 1285 -7481
rect 849 -7519 1080 -7513
rect 849 -7553 872 -7519
rect 906 -7547 1080 -7519
rect 1114 -7547 1152 -7513
rect 1186 -7547 1285 -7513
rect 906 -7553 1285 -7547
rect 1489 -7483 2593 -7465
rect 1489 -7513 1539 -7483
rect 1489 -7547 1532 -7513
rect 1591 -7535 1603 -7483
rect 1655 -7535 1667 -7483
rect 1719 -7535 1735 -7483
rect 1787 -7513 1799 -7483
rect 1851 -7513 1863 -7483
rect 1787 -7535 1790 -7513
rect 1851 -7535 1862 -7513
rect 1915 -7535 2025 -7483
rect 2077 -7513 2089 -7483
rect 2141 -7513 2153 -7483
rect 2082 -7535 2089 -7513
rect 2205 -7535 2221 -7483
rect 2273 -7535 2285 -7483
rect 2337 -7513 2349 -7483
rect 2401 -7513 2593 -7483
rect 2340 -7535 2349 -7513
rect 1566 -7547 1604 -7535
rect 1638 -7547 1790 -7535
rect 1824 -7547 1862 -7535
rect 1896 -7547 2048 -7535
rect 2082 -7547 2120 -7535
rect 2154 -7547 2306 -7535
rect 2340 -7547 2378 -7535
rect 2412 -7547 2593 -7513
rect 1489 -7553 2593 -7547
rect 2715 -7344 3423 -7327
rect 2715 -7396 2749 -7344
rect 2801 -7396 2813 -7344
rect 2865 -7396 2877 -7344
rect 2929 -7396 2945 -7344
rect 2997 -7396 3009 -7344
rect 3061 -7396 3073 -7344
rect 3125 -7396 3137 -7344
rect 3189 -7396 3205 -7344
rect 3257 -7396 3269 -7344
rect 3321 -7396 3333 -7344
rect 3385 -7396 3423 -7344
rect 2715 -7513 3423 -7396
rect 2715 -7547 2758 -7513
rect 2792 -7547 2830 -7513
rect 2864 -7547 3016 -7513
rect 3050 -7547 3088 -7513
rect 3122 -7547 3274 -7513
rect 3308 -7547 3346 -7513
rect 3380 -7547 3423 -7513
rect 2715 -7553 3423 -7547
rect 3545 -7465 3606 -7233
rect 3683 -7151 4649 -7145
rect 3683 -7185 3726 -7151
rect 3760 -7166 3798 -7151
rect 3832 -7166 3984 -7151
rect 4018 -7166 4056 -7151
rect 4090 -7166 4242 -7151
rect 4276 -7166 4314 -7151
rect 4348 -7166 4500 -7151
rect 4534 -7166 4572 -7151
rect 3789 -7185 3798 -7166
rect 3683 -7218 3737 -7185
rect 3789 -7218 3801 -7185
rect 3853 -7218 3865 -7166
rect 3917 -7218 3933 -7166
rect 4049 -7185 4056 -7166
rect 3985 -7218 3997 -7185
rect 4049 -7218 4061 -7185
rect 4113 -7218 4223 -7166
rect 4276 -7185 4287 -7166
rect 4348 -7185 4351 -7166
rect 4275 -7218 4287 -7185
rect 4339 -7218 4351 -7185
rect 4403 -7218 4419 -7166
rect 4471 -7218 4483 -7166
rect 4535 -7218 4547 -7166
rect 4606 -7185 4649 -7151
rect 4599 -7218 4649 -7185
rect 3683 -7344 4649 -7218
rect 3683 -7396 3737 -7344
rect 3789 -7396 3801 -7344
rect 3853 -7396 3865 -7344
rect 3917 -7396 3933 -7344
rect 3985 -7396 3997 -7344
rect 4049 -7396 4061 -7344
rect 4113 -7396 4223 -7344
rect 4275 -7396 4287 -7344
rect 4339 -7396 4351 -7344
rect 4403 -7396 4419 -7344
rect 4471 -7396 4483 -7344
rect 4535 -7396 4547 -7344
rect 4599 -7396 4649 -7344
rect 3683 -7415 4649 -7396
rect 4853 -7151 5643 -7121
rect 9210 -7121 9589 -7087
rect 9623 -7121 9646 -7087
rect 4853 -7185 4952 -7151
rect 4986 -7185 5024 -7151
rect 5058 -7159 5438 -7151
rect 5058 -7185 5231 -7159
rect 4853 -7193 5231 -7185
rect 5265 -7185 5438 -7159
rect 5472 -7185 5510 -7151
rect 5544 -7185 5643 -7151
rect 5265 -7193 5643 -7185
rect 4853 -7231 5643 -7193
rect 4853 -7265 5231 -7231
rect 5265 -7265 5643 -7231
rect 4853 -7303 5643 -7265
rect 4853 -7337 5231 -7303
rect 5265 -7337 5643 -7303
rect 4853 -7375 5643 -7337
rect 4853 -7409 5231 -7375
rect 5265 -7409 5643 -7375
rect 4853 -7447 5643 -7409
rect 5846 -7151 6812 -7145
rect 5846 -7185 5889 -7151
rect 5923 -7166 5961 -7151
rect 5995 -7166 6147 -7151
rect 6181 -7166 6219 -7151
rect 6253 -7166 6405 -7151
rect 6439 -7166 6477 -7151
rect 6511 -7166 6663 -7151
rect 6697 -7166 6735 -7151
rect 5846 -7218 5896 -7185
rect 5948 -7218 5960 -7166
rect 6012 -7218 6024 -7166
rect 6076 -7218 6092 -7166
rect 6144 -7185 6147 -7166
rect 6208 -7185 6219 -7166
rect 6144 -7218 6156 -7185
rect 6208 -7218 6220 -7185
rect 6272 -7218 6382 -7166
rect 6439 -7185 6446 -7166
rect 6434 -7218 6446 -7185
rect 6498 -7218 6510 -7185
rect 6562 -7218 6578 -7166
rect 6630 -7218 6642 -7166
rect 6697 -7185 6706 -7166
rect 6769 -7185 6812 -7151
rect 6694 -7218 6706 -7185
rect 6758 -7218 6812 -7185
rect 5846 -7344 6812 -7218
rect 5846 -7396 5896 -7344
rect 5948 -7396 5960 -7344
rect 6012 -7396 6024 -7344
rect 6076 -7396 6092 -7344
rect 6144 -7396 6156 -7344
rect 6208 -7396 6220 -7344
rect 6272 -7396 6382 -7344
rect 6434 -7396 6446 -7344
rect 6498 -7396 6510 -7344
rect 6562 -7396 6578 -7344
rect 6630 -7396 6642 -7344
rect 6694 -7396 6706 -7344
rect 6758 -7396 6812 -7344
rect 5846 -7415 6812 -7396
rect 6889 -7151 7963 -7145
rect 6889 -7185 7115 -7151
rect 7149 -7185 7187 -7151
rect 7221 -7185 7373 -7151
rect 7407 -7185 7445 -7151
rect 7479 -7185 7631 -7151
rect 7665 -7185 7703 -7151
rect 7737 -7185 7963 -7151
rect 6889 -7233 7963 -7185
rect 3545 -7483 4649 -7465
rect 3545 -7513 3737 -7483
rect 3789 -7513 3801 -7483
rect 3545 -7547 3726 -7513
rect 3789 -7535 3798 -7513
rect 3853 -7535 3865 -7483
rect 3917 -7535 3933 -7483
rect 3985 -7513 3997 -7483
rect 4049 -7513 4061 -7483
rect 4049 -7535 4056 -7513
rect 4113 -7535 4223 -7483
rect 4275 -7513 4287 -7483
rect 4339 -7513 4351 -7483
rect 4276 -7535 4287 -7513
rect 4348 -7535 4351 -7513
rect 4403 -7535 4419 -7483
rect 4471 -7535 4483 -7483
rect 4535 -7535 4547 -7483
rect 4599 -7513 4649 -7483
rect 3760 -7547 3798 -7535
rect 3832 -7547 3984 -7535
rect 4018 -7547 4056 -7535
rect 4090 -7547 4242 -7535
rect 4276 -7547 4314 -7535
rect 4348 -7547 4500 -7535
rect 4534 -7547 4572 -7535
rect 4606 -7547 4649 -7513
rect 3545 -7553 4649 -7547
rect 4853 -7481 5231 -7447
rect 5265 -7481 5643 -7447
rect 6889 -7465 6950 -7233
rect 4853 -7513 5643 -7481
rect 4853 -7547 4952 -7513
rect 4986 -7547 5024 -7513
rect 5058 -7519 5438 -7513
rect 5058 -7547 5231 -7519
rect 4853 -7553 5231 -7547
rect 5265 -7547 5438 -7519
rect 5472 -7547 5510 -7513
rect 5544 -7547 5643 -7513
rect 5265 -7553 5643 -7547
rect 5846 -7483 6950 -7465
rect 5846 -7513 5896 -7483
rect 5846 -7547 5889 -7513
rect 5948 -7535 5960 -7483
rect 6012 -7535 6024 -7483
rect 6076 -7535 6092 -7483
rect 6144 -7513 6156 -7483
rect 6208 -7513 6220 -7483
rect 6144 -7535 6147 -7513
rect 6208 -7535 6219 -7513
rect 6272 -7535 6382 -7483
rect 6434 -7513 6446 -7483
rect 6498 -7513 6510 -7483
rect 6439 -7535 6446 -7513
rect 6562 -7535 6578 -7483
rect 6630 -7535 6642 -7483
rect 6694 -7513 6706 -7483
rect 6758 -7513 6950 -7483
rect 6697 -7535 6706 -7513
rect 5923 -7547 5961 -7535
rect 5995 -7547 6147 -7535
rect 6181 -7547 6219 -7535
rect 6253 -7547 6405 -7535
rect 6439 -7547 6477 -7535
rect 6511 -7547 6663 -7535
rect 6697 -7547 6735 -7535
rect 6769 -7547 6950 -7513
rect 5846 -7553 6950 -7547
rect 7072 -7344 7780 -7327
rect 7072 -7396 7110 -7344
rect 7162 -7396 7174 -7344
rect 7226 -7396 7238 -7344
rect 7290 -7396 7306 -7344
rect 7358 -7396 7370 -7344
rect 7422 -7396 7434 -7344
rect 7486 -7396 7498 -7344
rect 7550 -7396 7566 -7344
rect 7618 -7396 7630 -7344
rect 7682 -7396 7694 -7344
rect 7746 -7396 7780 -7344
rect 7072 -7513 7780 -7396
rect 7072 -7547 7115 -7513
rect 7149 -7547 7187 -7513
rect 7221 -7547 7373 -7513
rect 7407 -7547 7445 -7513
rect 7479 -7547 7631 -7513
rect 7665 -7547 7703 -7513
rect 7737 -7547 7780 -7513
rect 7072 -7553 7780 -7547
rect 7902 -7465 7963 -7233
rect 8040 -7151 9006 -7145
rect 8040 -7185 8083 -7151
rect 8117 -7166 8155 -7151
rect 8189 -7166 8341 -7151
rect 8375 -7166 8413 -7151
rect 8447 -7166 8599 -7151
rect 8633 -7166 8671 -7151
rect 8705 -7166 8857 -7151
rect 8891 -7166 8929 -7151
rect 8146 -7185 8155 -7166
rect 8040 -7218 8094 -7185
rect 8146 -7218 8158 -7185
rect 8210 -7218 8222 -7166
rect 8274 -7218 8290 -7166
rect 8406 -7185 8413 -7166
rect 8342 -7218 8354 -7185
rect 8406 -7218 8418 -7185
rect 8470 -7218 8580 -7166
rect 8633 -7185 8644 -7166
rect 8705 -7185 8708 -7166
rect 8632 -7218 8644 -7185
rect 8696 -7218 8708 -7185
rect 8760 -7218 8776 -7166
rect 8828 -7218 8840 -7166
rect 8892 -7218 8904 -7166
rect 8963 -7185 9006 -7151
rect 8956 -7218 9006 -7185
rect 8040 -7344 9006 -7218
rect 8040 -7396 8094 -7344
rect 8146 -7396 8158 -7344
rect 8210 -7396 8222 -7344
rect 8274 -7396 8290 -7344
rect 8342 -7396 8354 -7344
rect 8406 -7396 8418 -7344
rect 8470 -7396 8580 -7344
rect 8632 -7396 8644 -7344
rect 8696 -7396 8708 -7344
rect 8760 -7396 8776 -7344
rect 8828 -7396 8840 -7344
rect 8892 -7396 8904 -7344
rect 8956 -7396 9006 -7344
rect 8040 -7415 9006 -7396
rect 9210 -7151 9646 -7121
rect 9210 -7185 9309 -7151
rect 9343 -7185 9381 -7151
rect 9415 -7159 9646 -7151
rect 9415 -7185 9589 -7159
rect 9210 -7193 9589 -7185
rect 9623 -7193 9646 -7159
rect 9210 -7231 9646 -7193
rect 9210 -7265 9589 -7231
rect 9623 -7265 9646 -7231
rect 9210 -7303 9646 -7265
rect 9210 -7337 9589 -7303
rect 9623 -7337 9646 -7303
rect 9210 -7375 9646 -7337
rect 9210 -7409 9589 -7375
rect 9623 -7409 9646 -7375
rect 9210 -7447 9646 -7409
rect 7902 -7483 9006 -7465
rect 7902 -7513 8094 -7483
rect 8146 -7513 8158 -7483
rect 7902 -7547 8083 -7513
rect 8146 -7535 8155 -7513
rect 8210 -7535 8222 -7483
rect 8274 -7535 8290 -7483
rect 8342 -7513 8354 -7483
rect 8406 -7513 8418 -7483
rect 8406 -7535 8413 -7513
rect 8470 -7535 8580 -7483
rect 8632 -7513 8644 -7483
rect 8696 -7513 8708 -7483
rect 8633 -7535 8644 -7513
rect 8705 -7535 8708 -7513
rect 8760 -7535 8776 -7483
rect 8828 -7535 8840 -7483
rect 8892 -7535 8904 -7483
rect 8956 -7513 9006 -7483
rect 8117 -7547 8155 -7535
rect 8189 -7547 8341 -7535
rect 8375 -7547 8413 -7535
rect 8447 -7547 8599 -7535
rect 8633 -7547 8671 -7535
rect 8705 -7547 8857 -7535
rect 8891 -7547 8929 -7535
rect 8963 -7547 9006 -7513
rect 7902 -7553 9006 -7547
rect 9210 -7481 9589 -7447
rect 9623 -7481 9646 -7447
rect 9210 -7513 9646 -7481
rect 9210 -7547 9309 -7513
rect 9343 -7547 9381 -7513
rect 9415 -7519 9646 -7513
rect 9415 -7547 9589 -7519
rect 9210 -7553 9589 -7547
rect 9623 -7553 9646 -7519
rect 849 -7591 1285 -7553
rect 849 -7625 872 -7591
rect 906 -7625 1285 -7591
rect 4853 -7591 5643 -7553
rect 849 -7641 1285 -7625
rect 849 -7663 987 -7641
rect 849 -7697 872 -7663
rect 906 -7675 987 -7663
rect 1021 -7675 1245 -7641
rect 1279 -7675 1285 -7641
rect 906 -7697 1285 -7675
rect 849 -7713 1285 -7697
rect 849 -7735 987 -7713
rect 849 -7769 872 -7735
rect 906 -7747 987 -7735
rect 1021 -7747 1245 -7713
rect 1279 -7747 1285 -7713
rect 906 -7769 1285 -7747
rect 849 -7807 1285 -7769
rect 849 -7841 872 -7807
rect 906 -7841 1285 -7807
rect 849 -7879 1285 -7841
rect 849 -7913 872 -7879
rect 906 -7913 1285 -7879
rect 849 -7951 1285 -7913
rect 849 -7985 872 -7951
rect 906 -7985 1285 -7951
rect 849 -8023 1285 -7985
rect 849 -8057 872 -8023
rect 906 -8057 1285 -8023
rect 849 -8095 1285 -8057
rect 849 -8129 872 -8095
rect 906 -8129 1285 -8095
rect 849 -8167 1285 -8129
rect 849 -8201 872 -8167
rect 906 -8201 1285 -8167
rect 849 -8239 1285 -8201
rect 1433 -7641 1479 -7594
rect 1433 -7675 1439 -7641
rect 1473 -7675 1479 -7641
rect 1433 -7713 1479 -7675
rect 1433 -7747 1439 -7713
rect 1473 -7747 1479 -7713
rect 1433 -8228 1479 -7747
rect 1691 -7641 1737 -7594
rect 1691 -7675 1697 -7641
rect 1731 -7675 1737 -7641
rect 1691 -7713 1737 -7675
rect 1691 -7747 1697 -7713
rect 1731 -7747 1737 -7713
rect 1691 -7896 1737 -7747
rect 1949 -7641 1995 -7594
rect 1949 -7675 1955 -7641
rect 1989 -7675 1995 -7641
rect 1949 -7713 1995 -7675
rect 1949 -7747 1955 -7713
rect 1989 -7747 1995 -7713
rect 1615 -7906 1811 -7896
rect 1615 -7958 1624 -7906
rect 1676 -7958 1688 -7906
rect 1740 -7958 1752 -7906
rect 1804 -7958 1811 -7906
rect 1615 -7966 1811 -7958
rect 1949 -8228 1995 -7747
rect 2207 -7641 2253 -7594
rect 2207 -7675 2213 -7641
rect 2247 -7675 2253 -7641
rect 2207 -7713 2253 -7675
rect 2207 -7747 2213 -7713
rect 2247 -7747 2253 -7713
rect 2207 -7896 2253 -7747
rect 2465 -7641 2511 -7594
rect 2465 -7675 2471 -7641
rect 2505 -7675 2511 -7641
rect 2465 -7713 2511 -7675
rect 2465 -7747 2471 -7713
rect 2505 -7747 2511 -7713
rect 2132 -7906 2328 -7896
rect 2132 -7958 2141 -7906
rect 2193 -7958 2205 -7906
rect 2257 -7958 2269 -7906
rect 2321 -7958 2328 -7906
rect 2132 -7966 2328 -7958
rect 2465 -8228 2511 -7747
rect 2659 -7641 2705 -7594
rect 2659 -7675 2665 -7641
rect 2699 -7675 2705 -7641
rect 2659 -7713 2705 -7675
rect 2659 -7747 2665 -7713
rect 2699 -7747 2705 -7713
rect 2659 -8065 2705 -7747
rect 2917 -7641 2963 -7594
rect 2917 -7675 2923 -7641
rect 2957 -7675 2963 -7641
rect 2917 -7713 2963 -7675
rect 2917 -7747 2923 -7713
rect 2957 -7747 2963 -7713
rect 2586 -8075 2782 -8065
rect 2586 -8127 2593 -8075
rect 2645 -8127 2657 -8075
rect 2709 -8127 2721 -8075
rect 2773 -8127 2782 -8075
rect 2586 -8135 2782 -8127
rect 849 -8273 872 -8239
rect 906 -8273 1285 -8239
rect 849 -8311 1285 -8273
rect 1355 -8238 1551 -8228
rect 1355 -8290 1364 -8238
rect 1416 -8290 1428 -8238
rect 1480 -8290 1492 -8238
rect 1544 -8290 1551 -8238
rect 1355 -8298 1551 -8290
rect 1873 -8238 2069 -8228
rect 1873 -8290 1882 -8238
rect 1934 -8290 1946 -8238
rect 1998 -8290 2010 -8238
rect 2062 -8290 2069 -8238
rect 1873 -8298 2069 -8290
rect 2389 -8238 2585 -8228
rect 2389 -8290 2398 -8238
rect 2450 -8290 2462 -8238
rect 2514 -8290 2526 -8238
rect 2578 -8290 2585 -8238
rect 2389 -8298 2585 -8290
rect 849 -8345 872 -8311
rect 906 -8345 1285 -8311
rect 849 -8383 1285 -8345
rect 849 -8417 872 -8383
rect 906 -8417 1285 -8383
rect 2917 -8396 2963 -7747
rect 3175 -7641 3221 -7594
rect 3175 -7675 3181 -7641
rect 3215 -7675 3221 -7641
rect 3175 -7713 3221 -7675
rect 3175 -7747 3181 -7713
rect 3215 -7747 3221 -7713
rect 3175 -8065 3221 -7747
rect 3433 -7641 3479 -7594
rect 3433 -7675 3439 -7641
rect 3473 -7675 3479 -7641
rect 3433 -7713 3479 -7675
rect 3433 -7747 3439 -7713
rect 3473 -7747 3479 -7713
rect 3103 -8075 3299 -8065
rect 3103 -8127 3110 -8075
rect 3162 -8127 3174 -8075
rect 3226 -8127 3238 -8075
rect 3290 -8127 3299 -8075
rect 3103 -8135 3299 -8127
rect 3433 -8396 3479 -7747
rect 3627 -7641 3673 -7594
rect 3627 -7675 3633 -7641
rect 3667 -7675 3673 -7641
rect 3627 -7713 3673 -7675
rect 3627 -7747 3633 -7713
rect 3667 -7747 3673 -7713
rect 3627 -8228 3673 -7747
rect 3885 -7641 3931 -7594
rect 3885 -7675 3891 -7641
rect 3925 -7675 3931 -7641
rect 3885 -7713 3931 -7675
rect 3885 -7747 3891 -7713
rect 3925 -7747 3931 -7713
rect 3885 -7896 3931 -7747
rect 4143 -7641 4189 -7594
rect 4143 -7675 4149 -7641
rect 4183 -7675 4189 -7641
rect 4143 -7713 4189 -7675
rect 4143 -7747 4149 -7713
rect 4183 -7747 4189 -7713
rect 3809 -7906 4005 -7896
rect 3809 -7958 3818 -7906
rect 3870 -7958 3882 -7906
rect 3934 -7958 3946 -7906
rect 3998 -7958 4005 -7906
rect 3809 -7966 4005 -7958
rect 4143 -8228 4189 -7747
rect 4401 -7641 4447 -7594
rect 4401 -7675 4407 -7641
rect 4441 -7675 4447 -7641
rect 4401 -7713 4447 -7675
rect 4401 -7747 4407 -7713
rect 4441 -7747 4447 -7713
rect 4401 -7896 4447 -7747
rect 4659 -7641 4705 -7594
rect 4659 -7675 4665 -7641
rect 4699 -7675 4705 -7641
rect 4659 -7713 4705 -7675
rect 4659 -7747 4665 -7713
rect 4699 -7747 4705 -7713
rect 4326 -7906 4522 -7896
rect 4326 -7958 4335 -7906
rect 4387 -7958 4399 -7906
rect 4451 -7958 4463 -7906
rect 4515 -7958 4522 -7906
rect 4326 -7966 4522 -7958
rect 4659 -8228 4705 -7747
rect 4853 -7625 5231 -7591
rect 5265 -7625 5643 -7591
rect 9210 -7591 9646 -7553
rect 4853 -7641 5643 -7625
rect 4853 -7675 4859 -7641
rect 4893 -7675 5117 -7641
rect 5151 -7663 5345 -7641
rect 5151 -7675 5231 -7663
rect 4853 -7697 5231 -7675
rect 5265 -7675 5345 -7663
rect 5379 -7675 5603 -7641
rect 5637 -7675 5643 -7641
rect 5265 -7697 5643 -7675
rect 4853 -7713 5643 -7697
rect 4853 -7747 4859 -7713
rect 4893 -7747 5117 -7713
rect 5151 -7735 5345 -7713
rect 5151 -7747 5231 -7735
rect 4853 -7769 5231 -7747
rect 5265 -7747 5345 -7735
rect 5379 -7747 5603 -7713
rect 5637 -7747 5643 -7713
rect 5265 -7769 5643 -7747
rect 4853 -7807 5643 -7769
rect 4853 -7841 5231 -7807
rect 5265 -7841 5643 -7807
rect 4853 -7879 5643 -7841
rect 4853 -7913 5231 -7879
rect 5265 -7913 5643 -7879
rect 4853 -7951 5643 -7913
rect 4853 -7985 5231 -7951
rect 5265 -7985 5643 -7951
rect 4853 -8023 5643 -7985
rect 4853 -8057 5231 -8023
rect 5265 -8057 5643 -8023
rect 4853 -8095 5643 -8057
rect 4853 -8129 5231 -8095
rect 5265 -8129 5643 -8095
rect 4853 -8167 5643 -8129
rect 4853 -8201 5231 -8167
rect 5265 -8201 5643 -8167
rect 3550 -8238 3746 -8228
rect 3550 -8290 3559 -8238
rect 3611 -8290 3623 -8238
rect 3675 -8290 3687 -8238
rect 3739 -8290 3746 -8238
rect 3550 -8298 3746 -8290
rect 4067 -8238 4263 -8228
rect 4067 -8290 4076 -8238
rect 4128 -8290 4140 -8238
rect 4192 -8290 4204 -8238
rect 4256 -8290 4263 -8238
rect 4067 -8298 4263 -8290
rect 4582 -8238 4778 -8228
rect 4582 -8290 4591 -8238
rect 4643 -8290 4655 -8238
rect 4707 -8290 4719 -8238
rect 4771 -8290 4778 -8238
rect 4582 -8298 4778 -8290
rect 4853 -8239 5643 -8201
rect 5790 -7641 5836 -7594
rect 5790 -7675 5796 -7641
rect 5830 -7675 5836 -7641
rect 5790 -7713 5836 -7675
rect 5790 -7747 5796 -7713
rect 5830 -7747 5836 -7713
rect 5790 -8228 5836 -7747
rect 6048 -7641 6094 -7594
rect 6048 -7675 6054 -7641
rect 6088 -7675 6094 -7641
rect 6048 -7713 6094 -7675
rect 6048 -7747 6054 -7713
rect 6088 -7747 6094 -7713
rect 6048 -7896 6094 -7747
rect 6306 -7641 6352 -7594
rect 6306 -7675 6312 -7641
rect 6346 -7675 6352 -7641
rect 6306 -7713 6352 -7675
rect 6306 -7747 6312 -7713
rect 6346 -7747 6352 -7713
rect 5973 -7906 6169 -7896
rect 5973 -7958 5980 -7906
rect 6032 -7958 6044 -7906
rect 6096 -7958 6108 -7906
rect 6160 -7958 6169 -7906
rect 5973 -7966 6169 -7958
rect 6306 -8228 6352 -7747
rect 6564 -7641 6610 -7594
rect 6564 -7675 6570 -7641
rect 6604 -7675 6610 -7641
rect 6564 -7713 6610 -7675
rect 6564 -7747 6570 -7713
rect 6604 -7747 6610 -7713
rect 6564 -7896 6610 -7747
rect 6822 -7641 6868 -7594
rect 6822 -7675 6828 -7641
rect 6862 -7675 6868 -7641
rect 6822 -7713 6868 -7675
rect 6822 -7747 6828 -7713
rect 6862 -7747 6868 -7713
rect 6490 -7906 6686 -7896
rect 6490 -7958 6497 -7906
rect 6549 -7958 6561 -7906
rect 6613 -7958 6625 -7906
rect 6677 -7958 6686 -7906
rect 6490 -7966 6686 -7958
rect 6822 -8228 6868 -7747
rect 7016 -7641 7062 -7594
rect 7016 -7675 7022 -7641
rect 7056 -7675 7062 -7641
rect 7016 -7713 7062 -7675
rect 7016 -7747 7022 -7713
rect 7056 -7747 7062 -7713
rect 4853 -8273 5231 -8239
rect 5265 -8273 5643 -8239
rect 4853 -8311 5643 -8273
rect 5717 -8238 5913 -8228
rect 5717 -8290 5724 -8238
rect 5776 -8290 5788 -8238
rect 5840 -8290 5852 -8238
rect 5904 -8290 5913 -8238
rect 5717 -8298 5913 -8290
rect 6232 -8238 6428 -8228
rect 6232 -8290 6239 -8238
rect 6291 -8290 6303 -8238
rect 6355 -8290 6367 -8238
rect 6419 -8290 6428 -8238
rect 6232 -8298 6428 -8290
rect 6749 -8238 6945 -8228
rect 6749 -8290 6756 -8238
rect 6808 -8290 6820 -8238
rect 6872 -8290 6884 -8238
rect 6936 -8290 6945 -8238
rect 6749 -8298 6945 -8290
rect 4853 -8345 5231 -8311
rect 5265 -8345 5643 -8311
rect 4853 -8383 5643 -8345
rect 849 -8455 1285 -8417
rect 849 -8489 872 -8455
rect 906 -8489 1285 -8455
rect 2843 -8406 3039 -8396
rect 2843 -8458 2850 -8406
rect 2902 -8458 2914 -8406
rect 2966 -8458 2978 -8406
rect 3030 -8458 3039 -8406
rect 2843 -8466 3039 -8458
rect 3361 -8406 3557 -8396
rect 3361 -8458 3368 -8406
rect 3420 -8458 3432 -8406
rect 3484 -8458 3496 -8406
rect 3548 -8458 3557 -8406
rect 3361 -8466 3557 -8458
rect 4853 -8417 5231 -8383
rect 5265 -8417 5643 -8383
rect 7016 -8396 7062 -7747
rect 7274 -7641 7320 -7594
rect 7274 -7675 7280 -7641
rect 7314 -7675 7320 -7641
rect 7274 -7713 7320 -7675
rect 7274 -7747 7280 -7713
rect 7314 -7747 7320 -7713
rect 7274 -8065 7320 -7747
rect 7532 -7641 7578 -7594
rect 7532 -7675 7538 -7641
rect 7572 -7675 7578 -7641
rect 7532 -7713 7578 -7675
rect 7532 -7747 7538 -7713
rect 7572 -7747 7578 -7713
rect 7196 -8075 7392 -8065
rect 7196 -8127 7205 -8075
rect 7257 -8127 7269 -8075
rect 7321 -8127 7333 -8075
rect 7385 -8127 7392 -8075
rect 7196 -8135 7392 -8127
rect 7532 -8396 7578 -7747
rect 7790 -7641 7836 -7594
rect 7790 -7675 7796 -7641
rect 7830 -7675 7836 -7641
rect 7790 -7713 7836 -7675
rect 7790 -7747 7796 -7713
rect 7830 -7747 7836 -7713
rect 7790 -8065 7836 -7747
rect 7984 -7641 8030 -7594
rect 7984 -7675 7990 -7641
rect 8024 -7675 8030 -7641
rect 7984 -7713 8030 -7675
rect 7984 -7747 7990 -7713
rect 8024 -7747 8030 -7713
rect 7713 -8075 7909 -8065
rect 7713 -8127 7722 -8075
rect 7774 -8127 7786 -8075
rect 7838 -8127 7850 -8075
rect 7902 -8127 7909 -8075
rect 7713 -8135 7909 -8127
rect 7984 -8228 8030 -7747
rect 8242 -7641 8288 -7594
rect 8242 -7675 8248 -7641
rect 8282 -7675 8288 -7641
rect 8242 -7713 8288 -7675
rect 8242 -7747 8248 -7713
rect 8282 -7747 8288 -7713
rect 8242 -7896 8288 -7747
rect 8500 -7641 8546 -7594
rect 8500 -7675 8506 -7641
rect 8540 -7675 8546 -7641
rect 8500 -7713 8546 -7675
rect 8500 -7747 8506 -7713
rect 8540 -7747 8546 -7713
rect 8167 -7906 8363 -7896
rect 8167 -7958 8174 -7906
rect 8226 -7958 8238 -7906
rect 8290 -7958 8302 -7906
rect 8354 -7958 8363 -7906
rect 8167 -7966 8363 -7958
rect 8500 -8228 8546 -7747
rect 8758 -7641 8804 -7594
rect 8758 -7675 8764 -7641
rect 8798 -7675 8804 -7641
rect 8758 -7713 8804 -7675
rect 8758 -7747 8764 -7713
rect 8798 -7747 8804 -7713
rect 8758 -7896 8804 -7747
rect 9016 -7641 9062 -7594
rect 9016 -7675 9022 -7641
rect 9056 -7675 9062 -7641
rect 9016 -7713 9062 -7675
rect 9016 -7747 9022 -7713
rect 9056 -7747 9062 -7713
rect 8685 -7906 8881 -7896
rect 8685 -7958 8692 -7906
rect 8744 -7958 8756 -7906
rect 8808 -7958 8820 -7906
rect 8872 -7958 8881 -7906
rect 8685 -7966 8881 -7958
rect 9016 -8228 9062 -7747
rect 9210 -7625 9589 -7591
rect 9623 -7625 9646 -7591
rect 9210 -7641 9646 -7625
rect 9210 -7675 9216 -7641
rect 9250 -7675 9474 -7641
rect 9508 -7663 9646 -7641
rect 9508 -7675 9589 -7663
rect 9210 -7697 9589 -7675
rect 9623 -7697 9646 -7663
rect 9210 -7713 9646 -7697
rect 9210 -7747 9216 -7713
rect 9250 -7747 9474 -7713
rect 9508 -7735 9646 -7713
rect 9508 -7747 9589 -7735
rect 9210 -7769 9589 -7747
rect 9623 -7769 9646 -7735
rect 9210 -7807 9646 -7769
rect 9210 -7841 9589 -7807
rect 9623 -7841 9646 -7807
rect 9210 -7879 9646 -7841
rect 9210 -7913 9589 -7879
rect 9623 -7913 9646 -7879
rect 9210 -7951 9646 -7913
rect 9210 -7985 9589 -7951
rect 9623 -7985 9646 -7951
rect 9210 -8023 9646 -7985
rect 9210 -8057 9589 -8023
rect 9623 -8057 9646 -8023
rect 9210 -8095 9646 -8057
rect 9210 -8129 9589 -8095
rect 9623 -8129 9646 -8095
rect 9210 -8167 9646 -8129
rect 9210 -8201 9589 -8167
rect 9623 -8201 9646 -8167
rect 7910 -8238 8106 -8228
rect 7910 -8290 7917 -8238
rect 7969 -8290 7981 -8238
rect 8033 -8290 8045 -8238
rect 8097 -8290 8106 -8238
rect 7910 -8298 8106 -8290
rect 8427 -8238 8623 -8228
rect 8427 -8290 8434 -8238
rect 8486 -8290 8498 -8238
rect 8550 -8290 8562 -8238
rect 8614 -8290 8623 -8238
rect 8427 -8298 8623 -8290
rect 8944 -8238 9140 -8228
rect 8944 -8290 8951 -8238
rect 9003 -8290 9015 -8238
rect 9067 -8290 9079 -8238
rect 9131 -8290 9140 -8238
rect 8944 -8298 9140 -8290
rect 9210 -8239 9646 -8201
rect 9210 -8273 9589 -8239
rect 9623 -8273 9646 -8239
rect 9210 -8311 9646 -8273
rect 9210 -8345 9589 -8311
rect 9623 -8345 9646 -8311
rect 9210 -8383 9646 -8345
rect 4853 -8455 5643 -8417
rect 849 -8527 1285 -8489
rect 849 -8561 872 -8527
rect 906 -8561 1285 -8527
rect 4853 -8489 5231 -8455
rect 5265 -8489 5643 -8455
rect 6939 -8406 7135 -8396
rect 6939 -8458 6948 -8406
rect 7000 -8458 7012 -8406
rect 7064 -8458 7076 -8406
rect 7128 -8458 7135 -8406
rect 6939 -8466 7135 -8458
rect 7456 -8406 7652 -8396
rect 7456 -8458 7465 -8406
rect 7517 -8458 7529 -8406
rect 7581 -8458 7593 -8406
rect 7645 -8458 7652 -8406
rect 7456 -8466 7652 -8458
rect 9210 -8417 9589 -8383
rect 9623 -8417 9646 -8383
rect 9210 -8455 9646 -8417
rect 4853 -8527 5643 -8489
rect 849 -8585 1285 -8561
rect 849 -8599 987 -8585
rect 849 -8633 872 -8599
rect 906 -8619 987 -8599
rect 1021 -8619 1245 -8585
rect 1279 -8619 1285 -8585
rect 906 -8633 1285 -8619
rect 849 -8657 1285 -8633
rect 849 -8671 987 -8657
rect 849 -8705 872 -8671
rect 906 -8691 987 -8671
rect 1021 -8691 1245 -8657
rect 1279 -8691 1285 -8657
rect 906 -8705 1285 -8691
rect 849 -8743 1285 -8705
rect 849 -8777 872 -8743
rect 906 -8777 1285 -8743
rect 849 -8779 1285 -8777
rect 1433 -8585 1479 -8538
rect 1433 -8619 1439 -8585
rect 1473 -8619 1479 -8585
rect 1433 -8657 1479 -8619
rect 1433 -8691 1439 -8657
rect 1473 -8691 1479 -8657
rect 1433 -8779 1479 -8691
rect 1691 -8585 1737 -8538
rect 1691 -8619 1697 -8585
rect 1731 -8619 1737 -8585
rect 1691 -8657 1737 -8619
rect 1691 -8691 1697 -8657
rect 1731 -8691 1737 -8657
rect 1691 -8779 1737 -8691
rect 1949 -8585 1995 -8538
rect 1949 -8619 1955 -8585
rect 1989 -8619 1995 -8585
rect 1949 -8657 1995 -8619
rect 1949 -8691 1955 -8657
rect 1989 -8691 1995 -8657
rect 1949 -8779 1995 -8691
rect 2207 -8585 2253 -8538
rect 2207 -8619 2213 -8585
rect 2247 -8619 2253 -8585
rect 2207 -8657 2253 -8619
rect 2207 -8691 2213 -8657
rect 2247 -8691 2253 -8657
rect 2207 -8779 2253 -8691
rect 2465 -8585 2511 -8538
rect 2465 -8619 2471 -8585
rect 2505 -8619 2511 -8585
rect 2465 -8657 2511 -8619
rect 2465 -8691 2471 -8657
rect 2505 -8691 2511 -8657
rect 2465 -8779 2511 -8691
rect 2659 -8585 2705 -8538
rect 2659 -8619 2665 -8585
rect 2699 -8619 2705 -8585
rect 2659 -8657 2705 -8619
rect 2659 -8691 2665 -8657
rect 2699 -8691 2705 -8657
rect 2659 -8779 2705 -8691
rect 2917 -8585 2963 -8538
rect 2917 -8619 2923 -8585
rect 2957 -8619 2963 -8585
rect 2917 -8657 2963 -8619
rect 2917 -8691 2923 -8657
rect 2957 -8691 2963 -8657
rect 2917 -8779 2963 -8691
rect 3175 -8585 3221 -8538
rect 3175 -8619 3181 -8585
rect 3215 -8619 3221 -8585
rect 3175 -8657 3221 -8619
rect 3175 -8691 3181 -8657
rect 3215 -8691 3221 -8657
rect 3175 -8779 3221 -8691
rect 3433 -8585 3479 -8538
rect 3433 -8619 3439 -8585
rect 3473 -8619 3479 -8585
rect 3433 -8657 3479 -8619
rect 3433 -8691 3439 -8657
rect 3473 -8691 3479 -8657
rect 3433 -8779 3479 -8691
rect 3627 -8585 3673 -8538
rect 3627 -8619 3633 -8585
rect 3667 -8619 3673 -8585
rect 3627 -8657 3673 -8619
rect 3627 -8691 3633 -8657
rect 3667 -8691 3673 -8657
rect 3627 -8779 3673 -8691
rect 3885 -8585 3931 -8538
rect 3885 -8619 3891 -8585
rect 3925 -8619 3931 -8585
rect 3885 -8657 3931 -8619
rect 3885 -8691 3891 -8657
rect 3925 -8691 3931 -8657
rect 3885 -8779 3931 -8691
rect 4143 -8585 4189 -8538
rect 4143 -8619 4149 -8585
rect 4183 -8619 4189 -8585
rect 4143 -8657 4189 -8619
rect 4143 -8691 4149 -8657
rect 4183 -8691 4189 -8657
rect 4143 -8779 4189 -8691
rect 4401 -8585 4447 -8538
rect 4401 -8619 4407 -8585
rect 4441 -8619 4447 -8585
rect 4401 -8657 4447 -8619
rect 4401 -8691 4407 -8657
rect 4441 -8691 4447 -8657
rect 4401 -8779 4447 -8691
rect 4659 -8585 4705 -8538
rect 4659 -8619 4665 -8585
rect 4699 -8619 4705 -8585
rect 4659 -8657 4705 -8619
rect 4659 -8691 4665 -8657
rect 4699 -8691 4705 -8657
rect 4659 -8779 4705 -8691
rect 4853 -8561 5231 -8527
rect 5265 -8561 5643 -8527
rect 9210 -8489 9589 -8455
rect 9623 -8489 9646 -8455
rect 9210 -8527 9646 -8489
rect 4853 -8585 5643 -8561
rect 4853 -8619 4859 -8585
rect 4893 -8619 5117 -8585
rect 5151 -8599 5345 -8585
rect 5151 -8619 5231 -8599
rect 4853 -8633 5231 -8619
rect 5265 -8619 5345 -8599
rect 5379 -8619 5603 -8585
rect 5637 -8619 5643 -8585
rect 5265 -8633 5643 -8619
rect 4853 -8657 5643 -8633
rect 4853 -8691 4859 -8657
rect 4893 -8691 5117 -8657
rect 5151 -8671 5345 -8657
rect 5151 -8691 5231 -8671
rect 4853 -8705 5231 -8691
rect 5265 -8691 5345 -8671
rect 5379 -8691 5603 -8657
rect 5637 -8691 5643 -8657
rect 5265 -8705 5643 -8691
rect 4853 -8743 5643 -8705
rect 4853 -8777 5231 -8743
rect 5265 -8777 5643 -8743
rect 4853 -8779 5643 -8777
rect 5790 -8585 5836 -8538
rect 5790 -8619 5796 -8585
rect 5830 -8619 5836 -8585
rect 5790 -8657 5836 -8619
rect 5790 -8691 5796 -8657
rect 5830 -8691 5836 -8657
rect 5790 -8779 5836 -8691
rect 6048 -8585 6094 -8538
rect 6048 -8619 6054 -8585
rect 6088 -8619 6094 -8585
rect 6048 -8657 6094 -8619
rect 6048 -8691 6054 -8657
rect 6088 -8691 6094 -8657
rect 6048 -8779 6094 -8691
rect 6306 -8585 6352 -8538
rect 6306 -8619 6312 -8585
rect 6346 -8619 6352 -8585
rect 6306 -8657 6352 -8619
rect 6306 -8691 6312 -8657
rect 6346 -8691 6352 -8657
rect 6306 -8779 6352 -8691
rect 6564 -8585 6610 -8538
rect 6564 -8619 6570 -8585
rect 6604 -8619 6610 -8585
rect 6564 -8657 6610 -8619
rect 6564 -8691 6570 -8657
rect 6604 -8691 6610 -8657
rect 6564 -8779 6610 -8691
rect 6822 -8585 6868 -8538
rect 6822 -8619 6828 -8585
rect 6862 -8619 6868 -8585
rect 6822 -8657 6868 -8619
rect 6822 -8691 6828 -8657
rect 6862 -8691 6868 -8657
rect 6822 -8779 6868 -8691
rect 7016 -8585 7062 -8538
rect 7016 -8619 7022 -8585
rect 7056 -8619 7062 -8585
rect 7016 -8657 7062 -8619
rect 7016 -8691 7022 -8657
rect 7056 -8691 7062 -8657
rect 7016 -8779 7062 -8691
rect 7274 -8585 7320 -8538
rect 7274 -8619 7280 -8585
rect 7314 -8619 7320 -8585
rect 7274 -8657 7320 -8619
rect 7274 -8691 7280 -8657
rect 7314 -8691 7320 -8657
rect 7274 -8779 7320 -8691
rect 7532 -8585 7578 -8538
rect 7532 -8619 7538 -8585
rect 7572 -8619 7578 -8585
rect 7532 -8657 7578 -8619
rect 7532 -8691 7538 -8657
rect 7572 -8691 7578 -8657
rect 7532 -8779 7578 -8691
rect 7790 -8585 7836 -8538
rect 7790 -8619 7796 -8585
rect 7830 -8619 7836 -8585
rect 7790 -8657 7836 -8619
rect 7790 -8691 7796 -8657
rect 7830 -8691 7836 -8657
rect 7790 -8779 7836 -8691
rect 7984 -8585 8030 -8538
rect 7984 -8619 7990 -8585
rect 8024 -8619 8030 -8585
rect 7984 -8657 8030 -8619
rect 7984 -8691 7990 -8657
rect 8024 -8691 8030 -8657
rect 7984 -8779 8030 -8691
rect 8242 -8585 8288 -8538
rect 8242 -8619 8248 -8585
rect 8282 -8619 8288 -8585
rect 8242 -8657 8288 -8619
rect 8242 -8691 8248 -8657
rect 8282 -8691 8288 -8657
rect 8242 -8779 8288 -8691
rect 8500 -8585 8546 -8538
rect 8500 -8619 8506 -8585
rect 8540 -8619 8546 -8585
rect 8500 -8657 8546 -8619
rect 8500 -8691 8506 -8657
rect 8540 -8691 8546 -8657
rect 8500 -8779 8546 -8691
rect 8758 -8585 8804 -8538
rect 8758 -8619 8764 -8585
rect 8798 -8619 8804 -8585
rect 8758 -8657 8804 -8619
rect 8758 -8691 8764 -8657
rect 8798 -8691 8804 -8657
rect 8758 -8779 8804 -8691
rect 9016 -8585 9062 -8538
rect 9016 -8619 9022 -8585
rect 9056 -8619 9062 -8585
rect 9016 -8657 9062 -8619
rect 9016 -8691 9022 -8657
rect 9056 -8691 9062 -8657
rect 9016 -8779 9062 -8691
rect 9210 -8561 9589 -8527
rect 9623 -8561 9646 -8527
rect 9210 -8585 9646 -8561
rect 9210 -8619 9216 -8585
rect 9250 -8619 9474 -8585
rect 9508 -8599 9646 -8585
rect 9508 -8619 9589 -8599
rect 9210 -8633 9589 -8619
rect 9623 -8633 9646 -8599
rect 9210 -8657 9646 -8633
rect 9210 -8691 9216 -8657
rect 9250 -8691 9474 -8657
rect 9508 -8671 9646 -8657
rect 9508 -8691 9589 -8671
rect 9210 -8705 9589 -8691
rect 9623 -8705 9646 -8671
rect 9210 -8743 9646 -8705
rect 9210 -8777 9589 -8743
rect 9623 -8777 9646 -8743
rect 9210 -8779 9646 -8777
rect 847 -8785 9648 -8779
rect 847 -8819 1080 -8785
rect 1114 -8819 1152 -8785
rect 1186 -8819 1532 -8785
rect 1566 -8819 1604 -8785
rect 1638 -8819 1790 -8785
rect 1824 -8819 1862 -8785
rect 1896 -8819 2048 -8785
rect 2082 -8819 2120 -8785
rect 2154 -8819 2306 -8785
rect 2340 -8819 2378 -8785
rect 2412 -8819 2758 -8785
rect 2792 -8819 2830 -8785
rect 2864 -8819 3016 -8785
rect 3050 -8819 3088 -8785
rect 3122 -8819 3274 -8785
rect 3308 -8819 3346 -8785
rect 3380 -8819 3726 -8785
rect 3760 -8819 3798 -8785
rect 3832 -8819 3984 -8785
rect 4018 -8819 4056 -8785
rect 4090 -8819 4242 -8785
rect 4276 -8819 4314 -8785
rect 4348 -8819 4500 -8785
rect 4534 -8819 4572 -8785
rect 4606 -8819 4952 -8785
rect 4986 -8819 5024 -8785
rect 5058 -8819 5438 -8785
rect 5472 -8819 5510 -8785
rect 5544 -8819 5889 -8785
rect 5923 -8819 5961 -8785
rect 5995 -8819 6147 -8785
rect 6181 -8819 6219 -8785
rect 6253 -8819 6405 -8785
rect 6439 -8819 6477 -8785
rect 6511 -8819 6663 -8785
rect 6697 -8819 6735 -8785
rect 6769 -8819 7115 -8785
rect 7149 -8819 7187 -8785
rect 7221 -8819 7373 -8785
rect 7407 -8819 7445 -8785
rect 7479 -8819 7631 -8785
rect 7665 -8819 7703 -8785
rect 7737 -8819 8083 -8785
rect 8117 -8819 8155 -8785
rect 8189 -8819 8341 -8785
rect 8375 -8819 8413 -8785
rect 8447 -8819 8599 -8785
rect 8633 -8819 8671 -8785
rect 8705 -8819 8857 -8785
rect 8891 -8819 8929 -8785
rect 8963 -8819 9309 -8785
rect 9343 -8819 9381 -8785
rect 9415 -8819 9648 -8785
rect 847 -8899 9648 -8819
rect 847 -8933 946 -8899
rect 980 -8933 1018 -8899
rect 1052 -8933 1090 -8899
rect 1124 -8933 1162 -8899
rect 1196 -8933 1234 -8899
rect 1268 -8933 1306 -8899
rect 1340 -8933 1378 -8899
rect 1412 -8933 1450 -8899
rect 1484 -8933 1522 -8899
rect 1556 -8933 1594 -8899
rect 1628 -8933 1666 -8899
rect 1700 -8933 1738 -8899
rect 1772 -8933 1810 -8899
rect 1844 -8933 1882 -8899
rect 1916 -8933 1954 -8899
rect 1988 -8933 2026 -8899
rect 2060 -8933 2098 -8899
rect 2132 -8933 2170 -8899
rect 2204 -8933 2242 -8899
rect 2276 -8933 2314 -8899
rect 2348 -8933 2386 -8899
rect 2420 -8933 2458 -8899
rect 2492 -8933 2530 -8899
rect 2564 -8933 2602 -8899
rect 2636 -8933 2674 -8899
rect 2708 -8933 2746 -8899
rect 2780 -8933 2818 -8899
rect 2852 -8933 2890 -8899
rect 2924 -8933 2962 -8899
rect 2996 -8933 3034 -8899
rect 3068 -8933 3106 -8899
rect 3140 -8933 3178 -8899
rect 3212 -8933 3250 -8899
rect 3284 -8933 3322 -8899
rect 3356 -8933 3394 -8899
rect 3428 -8933 3466 -8899
rect 3500 -8933 3538 -8899
rect 3572 -8933 3610 -8899
rect 3644 -8933 3682 -8899
rect 3716 -8933 3754 -8899
rect 3788 -8933 3826 -8899
rect 3860 -8933 3898 -8899
rect 3932 -8933 3970 -8899
rect 4004 -8933 4042 -8899
rect 4076 -8933 4114 -8899
rect 4148 -8933 4186 -8899
rect 4220 -8933 4258 -8899
rect 4292 -8933 4330 -8899
rect 4364 -8933 4402 -8899
rect 4436 -8933 4474 -8899
rect 4508 -8933 4546 -8899
rect 4580 -8933 4618 -8899
rect 4652 -8933 4690 -8899
rect 4724 -8933 4762 -8899
rect 4796 -8933 4834 -8899
rect 4868 -8933 4906 -8899
rect 4940 -8933 4978 -8899
rect 5012 -8933 5050 -8899
rect 5084 -8933 5122 -8899
rect 5156 -8933 5339 -8899
rect 5373 -8933 5411 -8899
rect 5445 -8933 5483 -8899
rect 5517 -8933 5555 -8899
rect 5589 -8933 5627 -8899
rect 5661 -8933 5699 -8899
rect 5733 -8933 5771 -8899
rect 5805 -8933 5843 -8899
rect 5877 -8933 5915 -8899
rect 5949 -8933 5987 -8899
rect 6021 -8933 6059 -8899
rect 6093 -8933 6131 -8899
rect 6165 -8933 6203 -8899
rect 6237 -8933 6275 -8899
rect 6309 -8933 6347 -8899
rect 6381 -8933 6419 -8899
rect 6453 -8933 6491 -8899
rect 6525 -8933 6563 -8899
rect 6597 -8933 6635 -8899
rect 6669 -8933 6707 -8899
rect 6741 -8933 6779 -8899
rect 6813 -8933 6851 -8899
rect 6885 -8933 6923 -8899
rect 6957 -8933 6995 -8899
rect 7029 -8933 7067 -8899
rect 7101 -8933 7139 -8899
rect 7173 -8933 7211 -8899
rect 7245 -8933 7283 -8899
rect 7317 -8933 7355 -8899
rect 7389 -8933 7427 -8899
rect 7461 -8933 7499 -8899
rect 7533 -8933 7571 -8899
rect 7605 -8933 7643 -8899
rect 7677 -8933 7715 -8899
rect 7749 -8933 7787 -8899
rect 7821 -8933 7859 -8899
rect 7893 -8933 7931 -8899
rect 7965 -8933 8003 -8899
rect 8037 -8933 8075 -8899
rect 8109 -8933 8147 -8899
rect 8181 -8933 8219 -8899
rect 8253 -8933 8291 -8899
rect 8325 -8933 8363 -8899
rect 8397 -8933 8435 -8899
rect 8469 -8933 8507 -8899
rect 8541 -8933 8579 -8899
rect 8613 -8933 8651 -8899
rect 8685 -8933 8723 -8899
rect 8757 -8933 8795 -8899
rect 8829 -8933 8867 -8899
rect 8901 -8933 8939 -8899
rect 8973 -8933 9011 -8899
rect 9045 -8933 9083 -8899
rect 9117 -8933 9155 -8899
rect 9189 -8933 9227 -8899
rect 9261 -8933 9299 -8899
rect 9333 -8933 9371 -8899
rect 9405 -8933 9443 -8899
rect 9477 -8933 9515 -8899
rect 9549 -8933 9648 -8899
rect 847 -8958 9648 -8933
<< via1 >>
rect 2850 229 2902 281
rect 2914 229 2966 281
rect 2978 229 3030 281
rect 3368 229 3420 281
rect 3432 229 3484 281
rect 3496 229 3548 281
rect 1364 60 1416 112
rect 1428 60 1480 112
rect 1492 60 1544 112
rect 1882 60 1934 112
rect 1946 60 1998 112
rect 2010 60 2062 112
rect 2398 60 2450 112
rect 2462 60 2514 112
rect 2526 60 2578 112
rect 1624 -271 1676 -219
rect 1688 -271 1740 -219
rect 1752 -271 1804 -219
rect 2141 -271 2193 -219
rect 2205 -271 2257 -219
rect 2269 -271 2321 -219
rect 2593 -103 2645 -51
rect 2657 -103 2709 -51
rect 2721 -103 2773 -51
rect 3110 -103 3162 -51
rect 3174 -103 3226 -51
rect 3238 -103 3290 -51
rect 6948 229 7000 281
rect 7012 229 7064 281
rect 7076 229 7128 281
rect 7465 229 7517 281
rect 7529 229 7581 281
rect 7593 229 7645 281
rect 3559 60 3611 112
rect 3623 60 3675 112
rect 3687 60 3739 112
rect 4076 60 4128 112
rect 4140 60 4192 112
rect 4204 60 4256 112
rect 4591 60 4643 112
rect 4655 60 4707 112
rect 4719 60 4771 112
rect 3818 -271 3870 -219
rect 3882 -271 3934 -219
rect 3946 -271 3998 -219
rect 4335 -271 4387 -219
rect 4399 -271 4451 -219
rect 4463 -271 4515 -219
rect 5724 60 5776 112
rect 5788 60 5840 112
rect 5852 60 5904 112
rect 6239 60 6291 112
rect 6303 60 6355 112
rect 6367 60 6419 112
rect 6756 60 6808 112
rect 6820 60 6872 112
rect 6884 60 6936 112
rect 5980 -271 6032 -219
rect 6044 -271 6096 -219
rect 6108 -271 6160 -219
rect 6497 -271 6549 -219
rect 6561 -271 6613 -219
rect 6625 -271 6677 -219
rect 7205 -103 7257 -51
rect 7269 -103 7321 -51
rect 7333 -103 7385 -51
rect 7917 60 7969 112
rect 7981 60 8033 112
rect 8045 60 8097 112
rect 8434 60 8486 112
rect 8498 60 8550 112
rect 8562 60 8614 112
rect 8951 60 9003 112
rect 9015 60 9067 112
rect 9079 60 9131 112
rect 7722 -103 7774 -51
rect 7786 -103 7838 -51
rect 7850 -103 7902 -51
rect 8174 -271 8226 -219
rect 8238 -271 8290 -219
rect 8302 -271 8354 -219
rect 8692 -271 8744 -219
rect 8756 -271 8808 -219
rect 8820 -271 8872 -219
rect 1539 -664 1566 -643
rect 1566 -664 1591 -643
rect 1539 -695 1591 -664
rect 1603 -664 1604 -643
rect 1604 -664 1638 -643
rect 1638 -664 1655 -643
rect 1603 -695 1655 -664
rect 1667 -695 1719 -643
rect 1735 -695 1787 -643
rect 1799 -664 1824 -643
rect 1824 -664 1851 -643
rect 1863 -664 1896 -643
rect 1896 -664 1915 -643
rect 1799 -695 1851 -664
rect 1863 -695 1915 -664
rect 2025 -664 2048 -643
rect 2048 -664 2077 -643
rect 2089 -664 2120 -643
rect 2120 -664 2141 -643
rect 2153 -664 2154 -643
rect 2154 -664 2205 -643
rect 2025 -695 2077 -664
rect 2089 -695 2141 -664
rect 2153 -695 2205 -664
rect 2221 -695 2273 -643
rect 2285 -664 2306 -643
rect 2306 -664 2337 -643
rect 2349 -664 2378 -643
rect 2378 -664 2401 -643
rect 2285 -695 2337 -664
rect 2349 -695 2401 -664
rect 1539 -833 1591 -781
rect 1603 -833 1655 -781
rect 1667 -833 1719 -781
rect 1735 -833 1787 -781
rect 1799 -833 1851 -781
rect 1863 -833 1915 -781
rect 2025 -833 2077 -781
rect 2089 -833 2141 -781
rect 2153 -833 2205 -781
rect 2221 -833 2273 -781
rect 2285 -833 2337 -781
rect 2349 -833 2401 -781
rect 1539 -993 1591 -959
rect 1539 -1011 1566 -993
rect 1566 -1011 1591 -993
rect 1603 -993 1655 -959
rect 1603 -1011 1604 -993
rect 1604 -1011 1638 -993
rect 1638 -1011 1655 -993
rect 1667 -1011 1719 -959
rect 1735 -1011 1787 -959
rect 1799 -993 1851 -959
rect 1863 -993 1915 -959
rect 1799 -1011 1824 -993
rect 1824 -1011 1851 -993
rect 1863 -1011 1896 -993
rect 1896 -1011 1915 -993
rect 2025 -993 2077 -959
rect 2089 -993 2141 -959
rect 2153 -993 2205 -959
rect 2025 -1011 2048 -993
rect 2048 -1011 2077 -993
rect 2089 -1011 2120 -993
rect 2120 -1011 2141 -993
rect 2153 -1011 2154 -993
rect 2154 -1011 2205 -993
rect 2221 -1011 2273 -959
rect 2285 -993 2337 -959
rect 2349 -993 2401 -959
rect 2285 -1011 2306 -993
rect 2306 -1011 2337 -993
rect 2349 -1011 2378 -993
rect 2378 -1011 2401 -993
rect 2749 -833 2801 -781
rect 2813 -833 2865 -781
rect 2877 -833 2929 -781
rect 2945 -833 2997 -781
rect 3009 -833 3061 -781
rect 3073 -833 3125 -781
rect 3137 -833 3189 -781
rect 3205 -833 3257 -781
rect 3269 -833 3321 -781
rect 3333 -833 3385 -781
rect 3737 -664 3760 -643
rect 3760 -664 3789 -643
rect 3801 -664 3832 -643
rect 3832 -664 3853 -643
rect 3737 -695 3789 -664
rect 3801 -695 3853 -664
rect 3865 -695 3917 -643
rect 3933 -664 3984 -643
rect 3984 -664 3985 -643
rect 3997 -664 4018 -643
rect 4018 -664 4049 -643
rect 4061 -664 4090 -643
rect 4090 -664 4113 -643
rect 3933 -695 3985 -664
rect 3997 -695 4049 -664
rect 4061 -695 4113 -664
rect 4223 -664 4242 -643
rect 4242 -664 4275 -643
rect 4287 -664 4314 -643
rect 4314 -664 4339 -643
rect 4223 -695 4275 -664
rect 4287 -695 4339 -664
rect 4351 -695 4403 -643
rect 4419 -695 4471 -643
rect 4483 -664 4500 -643
rect 4500 -664 4534 -643
rect 4534 -664 4535 -643
rect 4483 -695 4535 -664
rect 4547 -664 4572 -643
rect 4572 -664 4599 -643
rect 4547 -695 4599 -664
rect 5896 -664 5923 -643
rect 5923 -664 5948 -643
rect 5896 -695 5948 -664
rect 5960 -664 5961 -643
rect 5961 -664 5995 -643
rect 5995 -664 6012 -643
rect 5960 -695 6012 -664
rect 6024 -695 6076 -643
rect 6092 -695 6144 -643
rect 6156 -664 6181 -643
rect 6181 -664 6208 -643
rect 6220 -664 6253 -643
rect 6253 -664 6272 -643
rect 6156 -695 6208 -664
rect 6220 -695 6272 -664
rect 6382 -664 6405 -643
rect 6405 -664 6434 -643
rect 6446 -664 6477 -643
rect 6477 -664 6498 -643
rect 6510 -664 6511 -643
rect 6511 -664 6562 -643
rect 6382 -695 6434 -664
rect 6446 -695 6498 -664
rect 6510 -695 6562 -664
rect 6578 -695 6630 -643
rect 6642 -664 6663 -643
rect 6663 -664 6694 -643
rect 6706 -664 6735 -643
rect 6735 -664 6758 -643
rect 6642 -695 6694 -664
rect 6706 -695 6758 -664
rect 3737 -833 3789 -781
rect 3801 -833 3853 -781
rect 3865 -833 3917 -781
rect 3933 -833 3985 -781
rect 3997 -833 4049 -781
rect 4061 -833 4113 -781
rect 4223 -833 4275 -781
rect 4287 -833 4339 -781
rect 4351 -833 4403 -781
rect 4419 -833 4471 -781
rect 4483 -833 4535 -781
rect 4547 -833 4599 -781
rect 3737 -993 3789 -959
rect 3801 -993 3853 -959
rect 3737 -1011 3760 -993
rect 3760 -1011 3789 -993
rect 3801 -1011 3832 -993
rect 3832 -1011 3853 -993
rect 3865 -1011 3917 -959
rect 3933 -993 3985 -959
rect 3997 -993 4049 -959
rect 4061 -993 4113 -959
rect 3933 -1011 3984 -993
rect 3984 -1011 3985 -993
rect 3997 -1011 4018 -993
rect 4018 -1011 4049 -993
rect 4061 -1011 4090 -993
rect 4090 -1011 4113 -993
rect 4223 -993 4275 -959
rect 4287 -993 4339 -959
rect 4223 -1011 4242 -993
rect 4242 -1011 4275 -993
rect 4287 -1011 4314 -993
rect 4314 -1011 4339 -993
rect 4351 -1011 4403 -959
rect 4419 -1011 4471 -959
rect 4483 -993 4535 -959
rect 4483 -1011 4500 -993
rect 4500 -1011 4534 -993
rect 4534 -1011 4535 -993
rect 4547 -993 4599 -959
rect 4547 -1011 4572 -993
rect 4572 -1011 4599 -993
rect 5896 -833 5948 -781
rect 5960 -833 6012 -781
rect 6024 -833 6076 -781
rect 6092 -833 6144 -781
rect 6156 -833 6208 -781
rect 6220 -833 6272 -781
rect 6382 -833 6434 -781
rect 6446 -833 6498 -781
rect 6510 -833 6562 -781
rect 6578 -833 6630 -781
rect 6642 -833 6694 -781
rect 6706 -833 6758 -781
rect 5896 -993 5948 -959
rect 5896 -1011 5923 -993
rect 5923 -1011 5948 -993
rect 5960 -993 6012 -959
rect 5960 -1011 5961 -993
rect 5961 -1011 5995 -993
rect 5995 -1011 6012 -993
rect 6024 -1011 6076 -959
rect 6092 -1011 6144 -959
rect 6156 -993 6208 -959
rect 6220 -993 6272 -959
rect 6156 -1011 6181 -993
rect 6181 -1011 6208 -993
rect 6220 -1011 6253 -993
rect 6253 -1011 6272 -993
rect 6382 -993 6434 -959
rect 6446 -993 6498 -959
rect 6510 -993 6562 -959
rect 6382 -1011 6405 -993
rect 6405 -1011 6434 -993
rect 6446 -1011 6477 -993
rect 6477 -1011 6498 -993
rect 6510 -1011 6511 -993
rect 6511 -1011 6562 -993
rect 6578 -1011 6630 -959
rect 6642 -993 6694 -959
rect 6706 -993 6758 -959
rect 6642 -1011 6663 -993
rect 6663 -1011 6694 -993
rect 6706 -1011 6735 -993
rect 6735 -1011 6758 -993
rect 7110 -833 7162 -781
rect 7174 -833 7226 -781
rect 7238 -833 7290 -781
rect 7306 -833 7358 -781
rect 7370 -833 7422 -781
rect 7434 -833 7486 -781
rect 7498 -833 7550 -781
rect 7566 -833 7618 -781
rect 7630 -833 7682 -781
rect 7694 -833 7746 -781
rect 8094 -664 8117 -643
rect 8117 -664 8146 -643
rect 8158 -664 8189 -643
rect 8189 -664 8210 -643
rect 8094 -695 8146 -664
rect 8158 -695 8210 -664
rect 8222 -695 8274 -643
rect 8290 -664 8341 -643
rect 8341 -664 8342 -643
rect 8354 -664 8375 -643
rect 8375 -664 8406 -643
rect 8418 -664 8447 -643
rect 8447 -664 8470 -643
rect 8290 -695 8342 -664
rect 8354 -695 8406 -664
rect 8418 -695 8470 -664
rect 8580 -664 8599 -643
rect 8599 -664 8632 -643
rect 8644 -664 8671 -643
rect 8671 -664 8696 -643
rect 8580 -695 8632 -664
rect 8644 -695 8696 -664
rect 8708 -695 8760 -643
rect 8776 -695 8828 -643
rect 8840 -664 8857 -643
rect 8857 -664 8891 -643
rect 8891 -664 8892 -643
rect 8840 -695 8892 -664
rect 8904 -664 8929 -643
rect 8929 -664 8956 -643
rect 8904 -695 8956 -664
rect 8094 -833 8146 -781
rect 8158 -833 8210 -781
rect 8222 -833 8274 -781
rect 8290 -833 8342 -781
rect 8354 -833 8406 -781
rect 8418 -833 8470 -781
rect 8580 -833 8632 -781
rect 8644 -833 8696 -781
rect 8708 -833 8760 -781
rect 8776 -833 8828 -781
rect 8840 -833 8892 -781
rect 8904 -833 8956 -781
rect 8094 -993 8146 -959
rect 8158 -993 8210 -959
rect 8094 -1011 8117 -993
rect 8117 -1011 8146 -993
rect 8158 -1011 8189 -993
rect 8189 -1011 8210 -993
rect 8222 -1011 8274 -959
rect 8290 -993 8342 -959
rect 8354 -993 8406 -959
rect 8418 -993 8470 -959
rect 8290 -1011 8341 -993
rect 8341 -1011 8342 -993
rect 8354 -1011 8375 -993
rect 8375 -1011 8406 -993
rect 8418 -1011 8447 -993
rect 8447 -1011 8470 -993
rect 8580 -993 8632 -959
rect 8644 -993 8696 -959
rect 8580 -1011 8599 -993
rect 8599 -1011 8632 -993
rect 8644 -1011 8671 -993
rect 8671 -1011 8696 -993
rect 8708 -1011 8760 -959
rect 8776 -1011 8828 -959
rect 8840 -993 8892 -959
rect 8840 -1011 8857 -993
rect 8857 -1011 8891 -993
rect 8891 -1011 8892 -993
rect 8904 -993 8956 -959
rect 8904 -1011 8929 -993
rect 8929 -1011 8956 -993
rect 1367 -1461 1419 -1409
rect 1431 -1461 1483 -1409
rect 1495 -1461 1547 -1409
rect 1882 -1461 1934 -1409
rect 1946 -1461 1998 -1409
rect 2010 -1461 2062 -1409
rect 1625 -1762 1677 -1710
rect 1689 -1762 1741 -1710
rect 1753 -1762 1805 -1710
rect 2399 -1461 2451 -1409
rect 2463 -1461 2515 -1409
rect 2527 -1461 2579 -1409
rect 2142 -1762 2194 -1710
rect 2206 -1762 2258 -1710
rect 2270 -1762 2322 -1710
rect 2849 -1601 2901 -1549
rect 2913 -1601 2965 -1549
rect 2977 -1601 3029 -1549
rect 2591 -1906 2643 -1854
rect 2655 -1906 2707 -1854
rect 2719 -1906 2771 -1854
rect 3559 -1461 3611 -1409
rect 3623 -1461 3675 -1409
rect 3687 -1461 3739 -1409
rect 3366 -1601 3418 -1549
rect 3430 -1601 3482 -1549
rect 3494 -1601 3546 -1549
rect 3108 -1906 3160 -1854
rect 3172 -1906 3224 -1854
rect 3236 -1906 3288 -1854
rect 4076 -1461 4128 -1409
rect 4140 -1461 4192 -1409
rect 4204 -1461 4256 -1409
rect 3819 -1762 3871 -1710
rect 3883 -1762 3935 -1710
rect 3947 -1762 3999 -1710
rect 4593 -1461 4645 -1409
rect 4657 -1461 4709 -1409
rect 4721 -1461 4773 -1409
rect 4336 -1762 4388 -1710
rect 4400 -1762 4452 -1710
rect 4464 -1762 4516 -1710
rect 5722 -1461 5774 -1409
rect 5786 -1461 5838 -1409
rect 5850 -1461 5902 -1409
rect 6239 -1461 6291 -1409
rect 6303 -1461 6355 -1409
rect 6367 -1461 6419 -1409
rect 5979 -1762 6031 -1710
rect 6043 -1762 6095 -1710
rect 6107 -1762 6159 -1710
rect 6756 -1461 6808 -1409
rect 6820 -1461 6872 -1409
rect 6884 -1461 6936 -1409
rect 6496 -1762 6548 -1710
rect 6560 -1762 6612 -1710
rect 6624 -1762 6676 -1710
rect 6949 -1601 7001 -1549
rect 7013 -1601 7065 -1549
rect 7077 -1601 7129 -1549
rect 7466 -1601 7518 -1549
rect 7530 -1601 7582 -1549
rect 7594 -1601 7646 -1549
rect 7207 -1906 7259 -1854
rect 7271 -1906 7323 -1854
rect 7335 -1906 7387 -1854
rect 7916 -1461 7968 -1409
rect 7980 -1461 8032 -1409
rect 8044 -1461 8096 -1409
rect 7724 -1906 7776 -1854
rect 7788 -1906 7840 -1854
rect 7852 -1906 7904 -1854
rect 8434 -1461 8486 -1409
rect 8498 -1461 8550 -1409
rect 8562 -1461 8614 -1409
rect 8173 -1762 8225 -1710
rect 8237 -1762 8289 -1710
rect 8301 -1762 8353 -1710
rect 8949 -1461 9001 -1409
rect 9013 -1461 9065 -1409
rect 9077 -1461 9129 -1409
rect 8691 -1762 8743 -1710
rect 8755 -1762 8807 -1710
rect 8819 -1762 8871 -1710
rect 1539 -2311 1566 -2290
rect 1566 -2311 1591 -2290
rect 1539 -2342 1591 -2311
rect 1603 -2311 1604 -2290
rect 1604 -2311 1638 -2290
rect 1638 -2311 1655 -2290
rect 1603 -2342 1655 -2311
rect 1667 -2342 1719 -2290
rect 1735 -2342 1787 -2290
rect 1799 -2311 1824 -2290
rect 1824 -2311 1851 -2290
rect 1863 -2311 1896 -2290
rect 1896 -2311 1915 -2290
rect 1799 -2342 1851 -2311
rect 1863 -2342 1915 -2311
rect 2025 -2311 2048 -2290
rect 2048 -2311 2077 -2290
rect 2089 -2311 2120 -2290
rect 2120 -2311 2141 -2290
rect 2153 -2311 2154 -2290
rect 2154 -2311 2205 -2290
rect 2025 -2342 2077 -2311
rect 2089 -2342 2141 -2311
rect 2153 -2342 2205 -2311
rect 2221 -2342 2273 -2290
rect 2285 -2311 2306 -2290
rect 2306 -2311 2337 -2290
rect 2349 -2311 2378 -2290
rect 2378 -2311 2401 -2290
rect 2285 -2342 2337 -2311
rect 2349 -2342 2401 -2311
rect 1539 -2480 1591 -2428
rect 1603 -2480 1655 -2428
rect 1667 -2480 1719 -2428
rect 1735 -2480 1787 -2428
rect 1799 -2480 1851 -2428
rect 1863 -2480 1915 -2428
rect 2025 -2480 2077 -2428
rect 2089 -2480 2141 -2428
rect 2153 -2480 2205 -2428
rect 2221 -2480 2273 -2428
rect 2285 -2480 2337 -2428
rect 2349 -2480 2401 -2428
rect 1539 -2640 1591 -2606
rect 1539 -2658 1566 -2640
rect 1566 -2658 1591 -2640
rect 1603 -2640 1655 -2606
rect 1603 -2658 1604 -2640
rect 1604 -2658 1638 -2640
rect 1638 -2658 1655 -2640
rect 1667 -2658 1719 -2606
rect 1735 -2658 1787 -2606
rect 1799 -2640 1851 -2606
rect 1863 -2640 1915 -2606
rect 1799 -2658 1824 -2640
rect 1824 -2658 1851 -2640
rect 1863 -2658 1896 -2640
rect 1896 -2658 1915 -2640
rect 2025 -2640 2077 -2606
rect 2089 -2640 2141 -2606
rect 2153 -2640 2205 -2606
rect 2025 -2658 2048 -2640
rect 2048 -2658 2077 -2640
rect 2089 -2658 2120 -2640
rect 2120 -2658 2141 -2640
rect 2153 -2658 2154 -2640
rect 2154 -2658 2205 -2640
rect 2221 -2658 2273 -2606
rect 2285 -2640 2337 -2606
rect 2349 -2640 2401 -2606
rect 2285 -2658 2306 -2640
rect 2306 -2658 2337 -2640
rect 2349 -2658 2378 -2640
rect 2378 -2658 2401 -2640
rect 2749 -2480 2801 -2428
rect 2813 -2480 2865 -2428
rect 2877 -2480 2929 -2428
rect 2945 -2480 2997 -2428
rect 3009 -2480 3061 -2428
rect 3073 -2480 3125 -2428
rect 3137 -2480 3189 -2428
rect 3205 -2480 3257 -2428
rect 3269 -2480 3321 -2428
rect 3333 -2480 3385 -2428
rect 3737 -2311 3760 -2290
rect 3760 -2311 3789 -2290
rect 3801 -2311 3832 -2290
rect 3832 -2311 3853 -2290
rect 3737 -2342 3789 -2311
rect 3801 -2342 3853 -2311
rect 3865 -2342 3917 -2290
rect 3933 -2311 3984 -2290
rect 3984 -2311 3985 -2290
rect 3997 -2311 4018 -2290
rect 4018 -2311 4049 -2290
rect 4061 -2311 4090 -2290
rect 4090 -2311 4113 -2290
rect 3933 -2342 3985 -2311
rect 3997 -2342 4049 -2311
rect 4061 -2342 4113 -2311
rect 4223 -2311 4242 -2290
rect 4242 -2311 4275 -2290
rect 4287 -2311 4314 -2290
rect 4314 -2311 4339 -2290
rect 4223 -2342 4275 -2311
rect 4287 -2342 4339 -2311
rect 4351 -2342 4403 -2290
rect 4419 -2342 4471 -2290
rect 4483 -2311 4500 -2290
rect 4500 -2311 4534 -2290
rect 4534 -2311 4535 -2290
rect 4483 -2342 4535 -2311
rect 4547 -2311 4572 -2290
rect 4572 -2311 4599 -2290
rect 4547 -2342 4599 -2311
rect 5896 -2311 5923 -2290
rect 5923 -2311 5948 -2290
rect 5896 -2342 5948 -2311
rect 5960 -2311 5961 -2290
rect 5961 -2311 5995 -2290
rect 5995 -2311 6012 -2290
rect 5960 -2342 6012 -2311
rect 6024 -2342 6076 -2290
rect 6092 -2342 6144 -2290
rect 6156 -2311 6181 -2290
rect 6181 -2311 6208 -2290
rect 6220 -2311 6253 -2290
rect 6253 -2311 6272 -2290
rect 6156 -2342 6208 -2311
rect 6220 -2342 6272 -2311
rect 6382 -2311 6405 -2290
rect 6405 -2311 6434 -2290
rect 6446 -2311 6477 -2290
rect 6477 -2311 6498 -2290
rect 6510 -2311 6511 -2290
rect 6511 -2311 6562 -2290
rect 6382 -2342 6434 -2311
rect 6446 -2342 6498 -2311
rect 6510 -2342 6562 -2311
rect 6578 -2342 6630 -2290
rect 6642 -2311 6663 -2290
rect 6663 -2311 6694 -2290
rect 6706 -2311 6735 -2290
rect 6735 -2311 6758 -2290
rect 6642 -2342 6694 -2311
rect 6706 -2342 6758 -2311
rect 3737 -2480 3789 -2428
rect 3801 -2480 3853 -2428
rect 3865 -2480 3917 -2428
rect 3933 -2480 3985 -2428
rect 3997 -2480 4049 -2428
rect 4061 -2480 4113 -2428
rect 4223 -2480 4275 -2428
rect 4287 -2480 4339 -2428
rect 4351 -2480 4403 -2428
rect 4419 -2480 4471 -2428
rect 4483 -2480 4535 -2428
rect 4547 -2480 4599 -2428
rect 3737 -2640 3789 -2606
rect 3801 -2640 3853 -2606
rect 3737 -2658 3760 -2640
rect 3760 -2658 3789 -2640
rect 3801 -2658 3832 -2640
rect 3832 -2658 3853 -2640
rect 3865 -2658 3917 -2606
rect 3933 -2640 3985 -2606
rect 3997 -2640 4049 -2606
rect 4061 -2640 4113 -2606
rect 3933 -2658 3984 -2640
rect 3984 -2658 3985 -2640
rect 3997 -2658 4018 -2640
rect 4018 -2658 4049 -2640
rect 4061 -2658 4090 -2640
rect 4090 -2658 4113 -2640
rect 4223 -2640 4275 -2606
rect 4287 -2640 4339 -2606
rect 4223 -2658 4242 -2640
rect 4242 -2658 4275 -2640
rect 4287 -2658 4314 -2640
rect 4314 -2658 4339 -2640
rect 4351 -2658 4403 -2606
rect 4419 -2658 4471 -2606
rect 4483 -2640 4535 -2606
rect 4483 -2658 4500 -2640
rect 4500 -2658 4534 -2640
rect 4534 -2658 4535 -2640
rect 4547 -2640 4599 -2606
rect 4547 -2658 4572 -2640
rect 4572 -2658 4599 -2640
rect 5896 -2480 5948 -2428
rect 5960 -2480 6012 -2428
rect 6024 -2480 6076 -2428
rect 6092 -2480 6144 -2428
rect 6156 -2480 6208 -2428
rect 6220 -2480 6272 -2428
rect 6382 -2480 6434 -2428
rect 6446 -2480 6498 -2428
rect 6510 -2480 6562 -2428
rect 6578 -2480 6630 -2428
rect 6642 -2480 6694 -2428
rect 6706 -2480 6758 -2428
rect 5896 -2640 5948 -2606
rect 5896 -2658 5923 -2640
rect 5923 -2658 5948 -2640
rect 5960 -2640 6012 -2606
rect 5960 -2658 5961 -2640
rect 5961 -2658 5995 -2640
rect 5995 -2658 6012 -2640
rect 6024 -2658 6076 -2606
rect 6092 -2658 6144 -2606
rect 6156 -2640 6208 -2606
rect 6220 -2640 6272 -2606
rect 6156 -2658 6181 -2640
rect 6181 -2658 6208 -2640
rect 6220 -2658 6253 -2640
rect 6253 -2658 6272 -2640
rect 6382 -2640 6434 -2606
rect 6446 -2640 6498 -2606
rect 6510 -2640 6562 -2606
rect 6382 -2658 6405 -2640
rect 6405 -2658 6434 -2640
rect 6446 -2658 6477 -2640
rect 6477 -2658 6498 -2640
rect 6510 -2658 6511 -2640
rect 6511 -2658 6562 -2640
rect 6578 -2658 6630 -2606
rect 6642 -2640 6694 -2606
rect 6706 -2640 6758 -2606
rect 6642 -2658 6663 -2640
rect 6663 -2658 6694 -2640
rect 6706 -2658 6735 -2640
rect 6735 -2658 6758 -2640
rect 7110 -2480 7162 -2428
rect 7174 -2480 7226 -2428
rect 7238 -2480 7290 -2428
rect 7306 -2480 7358 -2428
rect 7370 -2480 7422 -2428
rect 7434 -2480 7486 -2428
rect 7498 -2480 7550 -2428
rect 7566 -2480 7618 -2428
rect 7630 -2480 7682 -2428
rect 7694 -2480 7746 -2428
rect 8094 -2311 8117 -2290
rect 8117 -2311 8146 -2290
rect 8158 -2311 8189 -2290
rect 8189 -2311 8210 -2290
rect 8094 -2342 8146 -2311
rect 8158 -2342 8210 -2311
rect 8222 -2342 8274 -2290
rect 8290 -2311 8341 -2290
rect 8341 -2311 8342 -2290
rect 8354 -2311 8375 -2290
rect 8375 -2311 8406 -2290
rect 8418 -2311 8447 -2290
rect 8447 -2311 8470 -2290
rect 8290 -2342 8342 -2311
rect 8354 -2342 8406 -2311
rect 8418 -2342 8470 -2311
rect 8580 -2311 8599 -2290
rect 8599 -2311 8632 -2290
rect 8644 -2311 8671 -2290
rect 8671 -2311 8696 -2290
rect 8580 -2342 8632 -2311
rect 8644 -2342 8696 -2311
rect 8708 -2342 8760 -2290
rect 8776 -2342 8828 -2290
rect 8840 -2311 8857 -2290
rect 8857 -2311 8891 -2290
rect 8891 -2311 8892 -2290
rect 8840 -2342 8892 -2311
rect 8904 -2311 8929 -2290
rect 8929 -2311 8956 -2290
rect 8904 -2342 8956 -2311
rect 8094 -2480 8146 -2428
rect 8158 -2480 8210 -2428
rect 8222 -2480 8274 -2428
rect 8290 -2480 8342 -2428
rect 8354 -2480 8406 -2428
rect 8418 -2480 8470 -2428
rect 8580 -2480 8632 -2428
rect 8644 -2480 8696 -2428
rect 8708 -2480 8760 -2428
rect 8776 -2480 8828 -2428
rect 8840 -2480 8892 -2428
rect 8904 -2480 8956 -2428
rect 8094 -2640 8146 -2606
rect 8158 -2640 8210 -2606
rect 8094 -2658 8117 -2640
rect 8117 -2658 8146 -2640
rect 8158 -2658 8189 -2640
rect 8189 -2658 8210 -2640
rect 8222 -2658 8274 -2606
rect 8290 -2640 8342 -2606
rect 8354 -2640 8406 -2606
rect 8418 -2640 8470 -2606
rect 8290 -2658 8341 -2640
rect 8341 -2658 8342 -2640
rect 8354 -2658 8375 -2640
rect 8375 -2658 8406 -2640
rect 8418 -2658 8447 -2640
rect 8447 -2658 8470 -2640
rect 8580 -2640 8632 -2606
rect 8644 -2640 8696 -2606
rect 8580 -2658 8599 -2640
rect 8599 -2658 8632 -2640
rect 8644 -2658 8671 -2640
rect 8671 -2658 8696 -2640
rect 8708 -2658 8760 -2606
rect 8776 -2658 8828 -2606
rect 8840 -2640 8892 -2606
rect 8840 -2658 8857 -2640
rect 8857 -2658 8891 -2640
rect 8891 -2658 8892 -2640
rect 8904 -2640 8956 -2606
rect 8904 -2658 8929 -2640
rect 8929 -2658 8956 -2640
rect 1624 -3085 1676 -3033
rect 1688 -3085 1740 -3033
rect 1752 -3085 1804 -3033
rect 2141 -3085 2193 -3033
rect 2205 -3085 2257 -3033
rect 2269 -3085 2321 -3033
rect 2593 -3254 2645 -3202
rect 2657 -3254 2709 -3202
rect 2721 -3254 2773 -3202
rect 1364 -3416 1416 -3364
rect 1428 -3416 1480 -3364
rect 1492 -3416 1544 -3364
rect 1882 -3416 1934 -3364
rect 1946 -3416 1998 -3364
rect 2010 -3416 2062 -3364
rect 2398 -3416 2450 -3364
rect 2462 -3416 2514 -3364
rect 2526 -3416 2578 -3364
rect 3110 -3254 3162 -3202
rect 3174 -3254 3226 -3202
rect 3238 -3254 3290 -3202
rect 3818 -3085 3870 -3033
rect 3882 -3085 3934 -3033
rect 3946 -3085 3998 -3033
rect 4335 -3085 4387 -3033
rect 4399 -3085 4451 -3033
rect 4463 -3085 4515 -3033
rect 3559 -3416 3611 -3364
rect 3623 -3416 3675 -3364
rect 3687 -3416 3739 -3364
rect 4076 -3416 4128 -3364
rect 4140 -3416 4192 -3364
rect 4204 -3416 4256 -3364
rect 4591 -3416 4643 -3364
rect 4655 -3416 4707 -3364
rect 4719 -3416 4771 -3364
rect 5980 -3085 6032 -3033
rect 6044 -3085 6096 -3033
rect 6108 -3085 6160 -3033
rect 6497 -3085 6549 -3033
rect 6561 -3085 6613 -3033
rect 6625 -3085 6677 -3033
rect 5724 -3416 5776 -3364
rect 5788 -3416 5840 -3364
rect 5852 -3416 5904 -3364
rect 6239 -3416 6291 -3364
rect 6303 -3416 6355 -3364
rect 6367 -3416 6419 -3364
rect 6756 -3416 6808 -3364
rect 6820 -3416 6872 -3364
rect 6884 -3416 6936 -3364
rect 2850 -3585 2902 -3533
rect 2914 -3585 2966 -3533
rect 2978 -3585 3030 -3533
rect 3368 -3585 3420 -3533
rect 3432 -3585 3484 -3533
rect 3496 -3585 3548 -3533
rect 7205 -3254 7257 -3202
rect 7269 -3254 7321 -3202
rect 7333 -3254 7385 -3202
rect 7722 -3254 7774 -3202
rect 7786 -3254 7838 -3202
rect 7850 -3254 7902 -3202
rect 8174 -3085 8226 -3033
rect 8238 -3085 8290 -3033
rect 8302 -3085 8354 -3033
rect 8692 -3085 8744 -3033
rect 8756 -3085 8808 -3033
rect 8820 -3085 8872 -3033
rect 7917 -3416 7969 -3364
rect 7981 -3416 8033 -3364
rect 8045 -3416 8097 -3364
rect 8434 -3416 8486 -3364
rect 8498 -3416 8550 -3364
rect 8562 -3416 8614 -3364
rect 8951 -3416 9003 -3364
rect 9015 -3416 9067 -3364
rect 9079 -3416 9131 -3364
rect 6948 -3585 7000 -3533
rect 7012 -3585 7064 -3533
rect 7076 -3585 7128 -3533
rect 7465 -3585 7517 -3533
rect 7529 -3585 7581 -3533
rect 7593 -3585 7645 -3533
rect 2850 -4644 2902 -4592
rect 2914 -4644 2966 -4592
rect 2978 -4644 3030 -4592
rect 3368 -4644 3420 -4592
rect 3432 -4644 3484 -4592
rect 3496 -4644 3548 -4592
rect 1364 -4813 1416 -4761
rect 1428 -4813 1480 -4761
rect 1492 -4813 1544 -4761
rect 1882 -4813 1934 -4761
rect 1946 -4813 1998 -4761
rect 2010 -4813 2062 -4761
rect 2398 -4813 2450 -4761
rect 2462 -4813 2514 -4761
rect 2526 -4813 2578 -4761
rect 1624 -5145 1676 -5093
rect 1688 -5145 1740 -5093
rect 1752 -5145 1804 -5093
rect 2141 -5145 2193 -5093
rect 2205 -5145 2257 -5093
rect 2269 -5145 2321 -5093
rect 2593 -4976 2645 -4924
rect 2657 -4976 2709 -4924
rect 2721 -4976 2773 -4924
rect 3110 -4976 3162 -4924
rect 3174 -4976 3226 -4924
rect 3238 -4976 3290 -4924
rect 6948 -4644 7000 -4592
rect 7012 -4644 7064 -4592
rect 7076 -4644 7128 -4592
rect 7465 -4644 7517 -4592
rect 7529 -4644 7581 -4592
rect 7593 -4644 7645 -4592
rect 3559 -4813 3611 -4761
rect 3623 -4813 3675 -4761
rect 3687 -4813 3739 -4761
rect 4076 -4813 4128 -4761
rect 4140 -4813 4192 -4761
rect 4204 -4813 4256 -4761
rect 4591 -4813 4643 -4761
rect 4655 -4813 4707 -4761
rect 4719 -4813 4771 -4761
rect 3818 -5145 3870 -5093
rect 3882 -5145 3934 -5093
rect 3946 -5145 3998 -5093
rect 4335 -5145 4387 -5093
rect 4399 -5145 4451 -5093
rect 4463 -5145 4515 -5093
rect 5724 -4813 5776 -4761
rect 5788 -4813 5840 -4761
rect 5852 -4813 5904 -4761
rect 6239 -4813 6291 -4761
rect 6303 -4813 6355 -4761
rect 6367 -4813 6419 -4761
rect 6756 -4813 6808 -4761
rect 6820 -4813 6872 -4761
rect 6884 -4813 6936 -4761
rect 5980 -5145 6032 -5093
rect 6044 -5145 6096 -5093
rect 6108 -5145 6160 -5093
rect 6497 -5145 6549 -5093
rect 6561 -5145 6613 -5093
rect 6625 -5145 6677 -5093
rect 7205 -4976 7257 -4924
rect 7269 -4976 7321 -4924
rect 7333 -4976 7385 -4924
rect 7917 -4813 7969 -4761
rect 7981 -4813 8033 -4761
rect 8045 -4813 8097 -4761
rect 8434 -4813 8486 -4761
rect 8498 -4813 8550 -4761
rect 8562 -4813 8614 -4761
rect 8951 -4813 9003 -4761
rect 9015 -4813 9067 -4761
rect 9079 -4813 9131 -4761
rect 7722 -4976 7774 -4924
rect 7786 -4976 7838 -4924
rect 7850 -4976 7902 -4924
rect 8174 -5145 8226 -5093
rect 8238 -5145 8290 -5093
rect 8302 -5145 8354 -5093
rect 8692 -5145 8744 -5093
rect 8756 -5145 8808 -5093
rect 8820 -5145 8872 -5093
rect 1539 -5538 1566 -5519
rect 1566 -5538 1591 -5519
rect 1539 -5571 1591 -5538
rect 1603 -5538 1604 -5519
rect 1604 -5538 1638 -5519
rect 1638 -5538 1655 -5519
rect 1603 -5571 1655 -5538
rect 1667 -5571 1719 -5519
rect 1735 -5571 1787 -5519
rect 1799 -5538 1824 -5519
rect 1824 -5538 1851 -5519
rect 1863 -5538 1896 -5519
rect 1896 -5538 1915 -5519
rect 1799 -5571 1851 -5538
rect 1863 -5571 1915 -5538
rect 2025 -5538 2048 -5519
rect 2048 -5538 2077 -5519
rect 2089 -5538 2120 -5519
rect 2120 -5538 2141 -5519
rect 2153 -5538 2154 -5519
rect 2154 -5538 2205 -5519
rect 2025 -5571 2077 -5538
rect 2089 -5571 2141 -5538
rect 2153 -5571 2205 -5538
rect 2221 -5571 2273 -5519
rect 2285 -5538 2306 -5519
rect 2306 -5538 2337 -5519
rect 2349 -5538 2378 -5519
rect 2378 -5538 2401 -5519
rect 2285 -5571 2337 -5538
rect 2349 -5571 2401 -5538
rect 1539 -5749 1591 -5697
rect 1603 -5749 1655 -5697
rect 1667 -5749 1719 -5697
rect 1735 -5749 1787 -5697
rect 1799 -5749 1851 -5697
rect 1863 -5749 1915 -5697
rect 2025 -5749 2077 -5697
rect 2089 -5749 2141 -5697
rect 2153 -5749 2205 -5697
rect 2221 -5749 2273 -5697
rect 2285 -5749 2337 -5697
rect 2349 -5749 2401 -5697
rect 1539 -5866 1591 -5836
rect 1539 -5888 1566 -5866
rect 1566 -5888 1591 -5866
rect 1603 -5866 1655 -5836
rect 1603 -5888 1604 -5866
rect 1604 -5888 1638 -5866
rect 1638 -5888 1655 -5866
rect 1667 -5888 1719 -5836
rect 1735 -5888 1787 -5836
rect 1799 -5866 1851 -5836
rect 1863 -5866 1915 -5836
rect 1799 -5888 1824 -5866
rect 1824 -5888 1851 -5866
rect 1863 -5888 1896 -5866
rect 1896 -5888 1915 -5866
rect 2025 -5866 2077 -5836
rect 2089 -5866 2141 -5836
rect 2153 -5866 2205 -5836
rect 2025 -5888 2048 -5866
rect 2048 -5888 2077 -5866
rect 2089 -5888 2120 -5866
rect 2120 -5888 2141 -5866
rect 2153 -5888 2154 -5866
rect 2154 -5888 2205 -5866
rect 2221 -5888 2273 -5836
rect 2285 -5866 2337 -5836
rect 2349 -5866 2401 -5836
rect 2285 -5888 2306 -5866
rect 2306 -5888 2337 -5866
rect 2349 -5888 2378 -5866
rect 2378 -5888 2401 -5866
rect 2749 -5749 2801 -5697
rect 2813 -5749 2865 -5697
rect 2877 -5749 2929 -5697
rect 2945 -5749 2997 -5697
rect 3009 -5749 3061 -5697
rect 3073 -5749 3125 -5697
rect 3137 -5749 3189 -5697
rect 3205 -5749 3257 -5697
rect 3269 -5749 3321 -5697
rect 3333 -5749 3385 -5697
rect 3737 -5538 3760 -5519
rect 3760 -5538 3789 -5519
rect 3801 -5538 3832 -5519
rect 3832 -5538 3853 -5519
rect 3737 -5571 3789 -5538
rect 3801 -5571 3853 -5538
rect 3865 -5571 3917 -5519
rect 3933 -5538 3984 -5519
rect 3984 -5538 3985 -5519
rect 3997 -5538 4018 -5519
rect 4018 -5538 4049 -5519
rect 4061 -5538 4090 -5519
rect 4090 -5538 4113 -5519
rect 3933 -5571 3985 -5538
rect 3997 -5571 4049 -5538
rect 4061 -5571 4113 -5538
rect 4223 -5538 4242 -5519
rect 4242 -5538 4275 -5519
rect 4287 -5538 4314 -5519
rect 4314 -5538 4339 -5519
rect 4223 -5571 4275 -5538
rect 4287 -5571 4339 -5538
rect 4351 -5571 4403 -5519
rect 4419 -5571 4471 -5519
rect 4483 -5538 4500 -5519
rect 4500 -5538 4534 -5519
rect 4534 -5538 4535 -5519
rect 4483 -5571 4535 -5538
rect 4547 -5538 4572 -5519
rect 4572 -5538 4599 -5519
rect 4547 -5571 4599 -5538
rect 3737 -5749 3789 -5697
rect 3801 -5749 3853 -5697
rect 3865 -5749 3917 -5697
rect 3933 -5749 3985 -5697
rect 3997 -5749 4049 -5697
rect 4061 -5749 4113 -5697
rect 4223 -5749 4275 -5697
rect 4287 -5749 4339 -5697
rect 4351 -5749 4403 -5697
rect 4419 -5749 4471 -5697
rect 4483 -5749 4535 -5697
rect 4547 -5749 4599 -5697
rect 5896 -5538 5923 -5519
rect 5923 -5538 5948 -5519
rect 5896 -5571 5948 -5538
rect 5960 -5538 5961 -5519
rect 5961 -5538 5995 -5519
rect 5995 -5538 6012 -5519
rect 5960 -5571 6012 -5538
rect 6024 -5571 6076 -5519
rect 6092 -5571 6144 -5519
rect 6156 -5538 6181 -5519
rect 6181 -5538 6208 -5519
rect 6220 -5538 6253 -5519
rect 6253 -5538 6272 -5519
rect 6156 -5571 6208 -5538
rect 6220 -5571 6272 -5538
rect 6382 -5538 6405 -5519
rect 6405 -5538 6434 -5519
rect 6446 -5538 6477 -5519
rect 6477 -5538 6498 -5519
rect 6510 -5538 6511 -5519
rect 6511 -5538 6562 -5519
rect 6382 -5571 6434 -5538
rect 6446 -5571 6498 -5538
rect 6510 -5571 6562 -5538
rect 6578 -5571 6630 -5519
rect 6642 -5538 6663 -5519
rect 6663 -5538 6694 -5519
rect 6706 -5538 6735 -5519
rect 6735 -5538 6758 -5519
rect 6642 -5571 6694 -5538
rect 6706 -5571 6758 -5538
rect 5896 -5749 5948 -5697
rect 5960 -5749 6012 -5697
rect 6024 -5749 6076 -5697
rect 6092 -5749 6144 -5697
rect 6156 -5749 6208 -5697
rect 6220 -5749 6272 -5697
rect 6382 -5749 6434 -5697
rect 6446 -5749 6498 -5697
rect 6510 -5749 6562 -5697
rect 6578 -5749 6630 -5697
rect 6642 -5749 6694 -5697
rect 6706 -5749 6758 -5697
rect 3737 -5866 3789 -5836
rect 3801 -5866 3853 -5836
rect 3737 -5888 3760 -5866
rect 3760 -5888 3789 -5866
rect 3801 -5888 3832 -5866
rect 3832 -5888 3853 -5866
rect 3865 -5888 3917 -5836
rect 3933 -5866 3985 -5836
rect 3997 -5866 4049 -5836
rect 4061 -5866 4113 -5836
rect 3933 -5888 3984 -5866
rect 3984 -5888 3985 -5866
rect 3997 -5888 4018 -5866
rect 4018 -5888 4049 -5866
rect 4061 -5888 4090 -5866
rect 4090 -5888 4113 -5866
rect 4223 -5866 4275 -5836
rect 4287 -5866 4339 -5836
rect 4223 -5888 4242 -5866
rect 4242 -5888 4275 -5866
rect 4287 -5888 4314 -5866
rect 4314 -5888 4339 -5866
rect 4351 -5888 4403 -5836
rect 4419 -5888 4471 -5836
rect 4483 -5866 4535 -5836
rect 4483 -5888 4500 -5866
rect 4500 -5888 4534 -5866
rect 4534 -5888 4535 -5866
rect 4547 -5866 4599 -5836
rect 4547 -5888 4572 -5866
rect 4572 -5888 4599 -5866
rect 5896 -5866 5948 -5836
rect 5896 -5888 5923 -5866
rect 5923 -5888 5948 -5866
rect 5960 -5866 6012 -5836
rect 5960 -5888 5961 -5866
rect 5961 -5888 5995 -5866
rect 5995 -5888 6012 -5866
rect 6024 -5888 6076 -5836
rect 6092 -5888 6144 -5836
rect 6156 -5866 6208 -5836
rect 6220 -5866 6272 -5836
rect 6156 -5888 6181 -5866
rect 6181 -5888 6208 -5866
rect 6220 -5888 6253 -5866
rect 6253 -5888 6272 -5866
rect 6382 -5866 6434 -5836
rect 6446 -5866 6498 -5836
rect 6510 -5866 6562 -5836
rect 6382 -5888 6405 -5866
rect 6405 -5888 6434 -5866
rect 6446 -5888 6477 -5866
rect 6477 -5888 6498 -5866
rect 6510 -5888 6511 -5866
rect 6511 -5888 6562 -5866
rect 6578 -5888 6630 -5836
rect 6642 -5866 6694 -5836
rect 6706 -5866 6758 -5836
rect 6642 -5888 6663 -5866
rect 6663 -5888 6694 -5866
rect 6706 -5888 6735 -5866
rect 6735 -5888 6758 -5866
rect 7110 -5749 7162 -5697
rect 7174 -5749 7226 -5697
rect 7238 -5749 7290 -5697
rect 7306 -5749 7358 -5697
rect 7370 -5749 7422 -5697
rect 7434 -5749 7486 -5697
rect 7498 -5749 7550 -5697
rect 7566 -5749 7618 -5697
rect 7630 -5749 7682 -5697
rect 7694 -5749 7746 -5697
rect 8094 -5538 8117 -5519
rect 8117 -5538 8146 -5519
rect 8158 -5538 8189 -5519
rect 8189 -5538 8210 -5519
rect 8094 -5571 8146 -5538
rect 8158 -5571 8210 -5538
rect 8222 -5571 8274 -5519
rect 8290 -5538 8341 -5519
rect 8341 -5538 8342 -5519
rect 8354 -5538 8375 -5519
rect 8375 -5538 8406 -5519
rect 8418 -5538 8447 -5519
rect 8447 -5538 8470 -5519
rect 8290 -5571 8342 -5538
rect 8354 -5571 8406 -5538
rect 8418 -5571 8470 -5538
rect 8580 -5538 8599 -5519
rect 8599 -5538 8632 -5519
rect 8644 -5538 8671 -5519
rect 8671 -5538 8696 -5519
rect 8580 -5571 8632 -5538
rect 8644 -5571 8696 -5538
rect 8708 -5571 8760 -5519
rect 8776 -5571 8828 -5519
rect 8840 -5538 8857 -5519
rect 8857 -5538 8891 -5519
rect 8891 -5538 8892 -5519
rect 8840 -5571 8892 -5538
rect 8904 -5538 8929 -5519
rect 8929 -5538 8956 -5519
rect 8904 -5571 8956 -5538
rect 8094 -5749 8146 -5697
rect 8158 -5749 8210 -5697
rect 8222 -5749 8274 -5697
rect 8290 -5749 8342 -5697
rect 8354 -5749 8406 -5697
rect 8418 -5749 8470 -5697
rect 8580 -5749 8632 -5697
rect 8644 -5749 8696 -5697
rect 8708 -5749 8760 -5697
rect 8776 -5749 8828 -5697
rect 8840 -5749 8892 -5697
rect 8904 -5749 8956 -5697
rect 8094 -5866 8146 -5836
rect 8158 -5866 8210 -5836
rect 8094 -5888 8117 -5866
rect 8117 -5888 8146 -5866
rect 8158 -5888 8189 -5866
rect 8189 -5888 8210 -5866
rect 8222 -5888 8274 -5836
rect 8290 -5866 8342 -5836
rect 8354 -5866 8406 -5836
rect 8418 -5866 8470 -5836
rect 8290 -5888 8341 -5866
rect 8341 -5888 8342 -5866
rect 8354 -5888 8375 -5866
rect 8375 -5888 8406 -5866
rect 8418 -5888 8447 -5866
rect 8447 -5888 8470 -5866
rect 8580 -5866 8632 -5836
rect 8644 -5866 8696 -5836
rect 8580 -5888 8599 -5866
rect 8599 -5888 8632 -5866
rect 8644 -5888 8671 -5866
rect 8671 -5888 8696 -5866
rect 8708 -5888 8760 -5836
rect 8776 -5888 8828 -5836
rect 8840 -5866 8892 -5836
rect 8840 -5888 8857 -5866
rect 8857 -5888 8891 -5866
rect 8891 -5888 8892 -5866
rect 8904 -5866 8956 -5836
rect 8904 -5888 8929 -5866
rect 8929 -5888 8956 -5866
rect 1625 -6468 1677 -6416
rect 1689 -6468 1741 -6416
rect 1753 -6468 1805 -6416
rect 1367 -6769 1419 -6717
rect 1431 -6769 1483 -6717
rect 1495 -6769 1547 -6717
rect 2142 -6468 2194 -6416
rect 2206 -6468 2258 -6416
rect 2270 -6468 2322 -6416
rect 1882 -6769 1934 -6717
rect 1946 -6769 1998 -6717
rect 2010 -6769 2062 -6717
rect 2591 -6323 2643 -6271
rect 2655 -6323 2707 -6271
rect 2719 -6323 2771 -6271
rect 2399 -6769 2451 -6717
rect 2463 -6769 2515 -6717
rect 2527 -6769 2579 -6717
rect 3108 -6323 3160 -6271
rect 3172 -6323 3224 -6271
rect 3236 -6323 3288 -6271
rect 2849 -6629 2901 -6577
rect 2913 -6629 2965 -6577
rect 2977 -6629 3029 -6577
rect 3366 -6629 3418 -6577
rect 3430 -6629 3482 -6577
rect 3494 -6629 3546 -6577
rect 3819 -6468 3871 -6416
rect 3883 -6468 3935 -6416
rect 3947 -6468 3999 -6416
rect 3559 -6769 3611 -6717
rect 3623 -6769 3675 -6717
rect 3687 -6769 3739 -6717
rect 4336 -6468 4388 -6416
rect 4400 -6468 4452 -6416
rect 4464 -6468 4516 -6416
rect 4076 -6769 4128 -6717
rect 4140 -6769 4192 -6717
rect 4204 -6769 4256 -6717
rect 4593 -6769 4645 -6717
rect 4657 -6769 4709 -6717
rect 4721 -6769 4773 -6717
rect 5979 -6468 6031 -6416
rect 6043 -6468 6095 -6416
rect 6107 -6468 6159 -6416
rect 5722 -6769 5774 -6717
rect 5786 -6769 5838 -6717
rect 5850 -6769 5902 -6717
rect 6496 -6468 6548 -6416
rect 6560 -6468 6612 -6416
rect 6624 -6468 6676 -6416
rect 6239 -6769 6291 -6717
rect 6303 -6769 6355 -6717
rect 6367 -6769 6419 -6717
rect 7207 -6323 7259 -6271
rect 7271 -6323 7323 -6271
rect 7335 -6323 7387 -6271
rect 6949 -6629 7001 -6577
rect 7013 -6629 7065 -6577
rect 7077 -6629 7129 -6577
rect 6756 -6769 6808 -6717
rect 6820 -6769 6872 -6717
rect 6884 -6769 6936 -6717
rect 7724 -6323 7776 -6271
rect 7788 -6323 7840 -6271
rect 7852 -6323 7904 -6271
rect 7466 -6629 7518 -6577
rect 7530 -6629 7582 -6577
rect 7594 -6629 7646 -6577
rect 8173 -6468 8225 -6416
rect 8237 -6468 8289 -6416
rect 8301 -6468 8353 -6416
rect 7916 -6769 7968 -6717
rect 7980 -6769 8032 -6717
rect 8044 -6769 8096 -6717
rect 8691 -6468 8743 -6416
rect 8755 -6468 8807 -6416
rect 8819 -6468 8871 -6416
rect 8434 -6769 8486 -6717
rect 8498 -6769 8550 -6717
rect 8562 -6769 8614 -6717
rect 8949 -6769 9001 -6717
rect 9013 -6769 9065 -6717
rect 9077 -6769 9129 -6717
rect 1539 -7185 1566 -7166
rect 1566 -7185 1591 -7166
rect 1539 -7218 1591 -7185
rect 1603 -7185 1604 -7166
rect 1604 -7185 1638 -7166
rect 1638 -7185 1655 -7166
rect 1603 -7218 1655 -7185
rect 1667 -7218 1719 -7166
rect 1735 -7218 1787 -7166
rect 1799 -7185 1824 -7166
rect 1824 -7185 1851 -7166
rect 1863 -7185 1896 -7166
rect 1896 -7185 1915 -7166
rect 1799 -7218 1851 -7185
rect 1863 -7218 1915 -7185
rect 2025 -7185 2048 -7166
rect 2048 -7185 2077 -7166
rect 2089 -7185 2120 -7166
rect 2120 -7185 2141 -7166
rect 2153 -7185 2154 -7166
rect 2154 -7185 2205 -7166
rect 2025 -7218 2077 -7185
rect 2089 -7218 2141 -7185
rect 2153 -7218 2205 -7185
rect 2221 -7218 2273 -7166
rect 2285 -7185 2306 -7166
rect 2306 -7185 2337 -7166
rect 2349 -7185 2378 -7166
rect 2378 -7185 2401 -7166
rect 2285 -7218 2337 -7185
rect 2349 -7218 2401 -7185
rect 1539 -7396 1591 -7344
rect 1603 -7396 1655 -7344
rect 1667 -7396 1719 -7344
rect 1735 -7396 1787 -7344
rect 1799 -7396 1851 -7344
rect 1863 -7396 1915 -7344
rect 2025 -7396 2077 -7344
rect 2089 -7396 2141 -7344
rect 2153 -7396 2205 -7344
rect 2221 -7396 2273 -7344
rect 2285 -7396 2337 -7344
rect 2349 -7396 2401 -7344
rect 1539 -7513 1591 -7483
rect 1539 -7535 1566 -7513
rect 1566 -7535 1591 -7513
rect 1603 -7513 1655 -7483
rect 1603 -7535 1604 -7513
rect 1604 -7535 1638 -7513
rect 1638 -7535 1655 -7513
rect 1667 -7535 1719 -7483
rect 1735 -7535 1787 -7483
rect 1799 -7513 1851 -7483
rect 1863 -7513 1915 -7483
rect 1799 -7535 1824 -7513
rect 1824 -7535 1851 -7513
rect 1863 -7535 1896 -7513
rect 1896 -7535 1915 -7513
rect 2025 -7513 2077 -7483
rect 2089 -7513 2141 -7483
rect 2153 -7513 2205 -7483
rect 2025 -7535 2048 -7513
rect 2048 -7535 2077 -7513
rect 2089 -7535 2120 -7513
rect 2120 -7535 2141 -7513
rect 2153 -7535 2154 -7513
rect 2154 -7535 2205 -7513
rect 2221 -7535 2273 -7483
rect 2285 -7513 2337 -7483
rect 2349 -7513 2401 -7483
rect 2285 -7535 2306 -7513
rect 2306 -7535 2337 -7513
rect 2349 -7535 2378 -7513
rect 2378 -7535 2401 -7513
rect 2749 -7396 2801 -7344
rect 2813 -7396 2865 -7344
rect 2877 -7396 2929 -7344
rect 2945 -7396 2997 -7344
rect 3009 -7396 3061 -7344
rect 3073 -7396 3125 -7344
rect 3137 -7396 3189 -7344
rect 3205 -7396 3257 -7344
rect 3269 -7396 3321 -7344
rect 3333 -7396 3385 -7344
rect 3737 -7185 3760 -7166
rect 3760 -7185 3789 -7166
rect 3801 -7185 3832 -7166
rect 3832 -7185 3853 -7166
rect 3737 -7218 3789 -7185
rect 3801 -7218 3853 -7185
rect 3865 -7218 3917 -7166
rect 3933 -7185 3984 -7166
rect 3984 -7185 3985 -7166
rect 3997 -7185 4018 -7166
rect 4018 -7185 4049 -7166
rect 4061 -7185 4090 -7166
rect 4090 -7185 4113 -7166
rect 3933 -7218 3985 -7185
rect 3997 -7218 4049 -7185
rect 4061 -7218 4113 -7185
rect 4223 -7185 4242 -7166
rect 4242 -7185 4275 -7166
rect 4287 -7185 4314 -7166
rect 4314 -7185 4339 -7166
rect 4223 -7218 4275 -7185
rect 4287 -7218 4339 -7185
rect 4351 -7218 4403 -7166
rect 4419 -7218 4471 -7166
rect 4483 -7185 4500 -7166
rect 4500 -7185 4534 -7166
rect 4534 -7185 4535 -7166
rect 4483 -7218 4535 -7185
rect 4547 -7185 4572 -7166
rect 4572 -7185 4599 -7166
rect 4547 -7218 4599 -7185
rect 3737 -7396 3789 -7344
rect 3801 -7396 3853 -7344
rect 3865 -7396 3917 -7344
rect 3933 -7396 3985 -7344
rect 3997 -7396 4049 -7344
rect 4061 -7396 4113 -7344
rect 4223 -7396 4275 -7344
rect 4287 -7396 4339 -7344
rect 4351 -7396 4403 -7344
rect 4419 -7396 4471 -7344
rect 4483 -7396 4535 -7344
rect 4547 -7396 4599 -7344
rect 5896 -7185 5923 -7166
rect 5923 -7185 5948 -7166
rect 5896 -7218 5948 -7185
rect 5960 -7185 5961 -7166
rect 5961 -7185 5995 -7166
rect 5995 -7185 6012 -7166
rect 5960 -7218 6012 -7185
rect 6024 -7218 6076 -7166
rect 6092 -7218 6144 -7166
rect 6156 -7185 6181 -7166
rect 6181 -7185 6208 -7166
rect 6220 -7185 6253 -7166
rect 6253 -7185 6272 -7166
rect 6156 -7218 6208 -7185
rect 6220 -7218 6272 -7185
rect 6382 -7185 6405 -7166
rect 6405 -7185 6434 -7166
rect 6446 -7185 6477 -7166
rect 6477 -7185 6498 -7166
rect 6510 -7185 6511 -7166
rect 6511 -7185 6562 -7166
rect 6382 -7218 6434 -7185
rect 6446 -7218 6498 -7185
rect 6510 -7218 6562 -7185
rect 6578 -7218 6630 -7166
rect 6642 -7185 6663 -7166
rect 6663 -7185 6694 -7166
rect 6706 -7185 6735 -7166
rect 6735 -7185 6758 -7166
rect 6642 -7218 6694 -7185
rect 6706 -7218 6758 -7185
rect 5896 -7396 5948 -7344
rect 5960 -7396 6012 -7344
rect 6024 -7396 6076 -7344
rect 6092 -7396 6144 -7344
rect 6156 -7396 6208 -7344
rect 6220 -7396 6272 -7344
rect 6382 -7396 6434 -7344
rect 6446 -7396 6498 -7344
rect 6510 -7396 6562 -7344
rect 6578 -7396 6630 -7344
rect 6642 -7396 6694 -7344
rect 6706 -7396 6758 -7344
rect 3737 -7513 3789 -7483
rect 3801 -7513 3853 -7483
rect 3737 -7535 3760 -7513
rect 3760 -7535 3789 -7513
rect 3801 -7535 3832 -7513
rect 3832 -7535 3853 -7513
rect 3865 -7535 3917 -7483
rect 3933 -7513 3985 -7483
rect 3997 -7513 4049 -7483
rect 4061 -7513 4113 -7483
rect 3933 -7535 3984 -7513
rect 3984 -7535 3985 -7513
rect 3997 -7535 4018 -7513
rect 4018 -7535 4049 -7513
rect 4061 -7535 4090 -7513
rect 4090 -7535 4113 -7513
rect 4223 -7513 4275 -7483
rect 4287 -7513 4339 -7483
rect 4223 -7535 4242 -7513
rect 4242 -7535 4275 -7513
rect 4287 -7535 4314 -7513
rect 4314 -7535 4339 -7513
rect 4351 -7535 4403 -7483
rect 4419 -7535 4471 -7483
rect 4483 -7513 4535 -7483
rect 4483 -7535 4500 -7513
rect 4500 -7535 4534 -7513
rect 4534 -7535 4535 -7513
rect 4547 -7513 4599 -7483
rect 4547 -7535 4572 -7513
rect 4572 -7535 4599 -7513
rect 5896 -7513 5948 -7483
rect 5896 -7535 5923 -7513
rect 5923 -7535 5948 -7513
rect 5960 -7513 6012 -7483
rect 5960 -7535 5961 -7513
rect 5961 -7535 5995 -7513
rect 5995 -7535 6012 -7513
rect 6024 -7535 6076 -7483
rect 6092 -7535 6144 -7483
rect 6156 -7513 6208 -7483
rect 6220 -7513 6272 -7483
rect 6156 -7535 6181 -7513
rect 6181 -7535 6208 -7513
rect 6220 -7535 6253 -7513
rect 6253 -7535 6272 -7513
rect 6382 -7513 6434 -7483
rect 6446 -7513 6498 -7483
rect 6510 -7513 6562 -7483
rect 6382 -7535 6405 -7513
rect 6405 -7535 6434 -7513
rect 6446 -7535 6477 -7513
rect 6477 -7535 6498 -7513
rect 6510 -7535 6511 -7513
rect 6511 -7535 6562 -7513
rect 6578 -7535 6630 -7483
rect 6642 -7513 6694 -7483
rect 6706 -7513 6758 -7483
rect 6642 -7535 6663 -7513
rect 6663 -7535 6694 -7513
rect 6706 -7535 6735 -7513
rect 6735 -7535 6758 -7513
rect 7110 -7396 7162 -7344
rect 7174 -7396 7226 -7344
rect 7238 -7396 7290 -7344
rect 7306 -7396 7358 -7344
rect 7370 -7396 7422 -7344
rect 7434 -7396 7486 -7344
rect 7498 -7396 7550 -7344
rect 7566 -7396 7618 -7344
rect 7630 -7396 7682 -7344
rect 7694 -7396 7746 -7344
rect 8094 -7185 8117 -7166
rect 8117 -7185 8146 -7166
rect 8158 -7185 8189 -7166
rect 8189 -7185 8210 -7166
rect 8094 -7218 8146 -7185
rect 8158 -7218 8210 -7185
rect 8222 -7218 8274 -7166
rect 8290 -7185 8341 -7166
rect 8341 -7185 8342 -7166
rect 8354 -7185 8375 -7166
rect 8375 -7185 8406 -7166
rect 8418 -7185 8447 -7166
rect 8447 -7185 8470 -7166
rect 8290 -7218 8342 -7185
rect 8354 -7218 8406 -7185
rect 8418 -7218 8470 -7185
rect 8580 -7185 8599 -7166
rect 8599 -7185 8632 -7166
rect 8644 -7185 8671 -7166
rect 8671 -7185 8696 -7166
rect 8580 -7218 8632 -7185
rect 8644 -7218 8696 -7185
rect 8708 -7218 8760 -7166
rect 8776 -7218 8828 -7166
rect 8840 -7185 8857 -7166
rect 8857 -7185 8891 -7166
rect 8891 -7185 8892 -7166
rect 8840 -7218 8892 -7185
rect 8904 -7185 8929 -7166
rect 8929 -7185 8956 -7166
rect 8904 -7218 8956 -7185
rect 8094 -7396 8146 -7344
rect 8158 -7396 8210 -7344
rect 8222 -7396 8274 -7344
rect 8290 -7396 8342 -7344
rect 8354 -7396 8406 -7344
rect 8418 -7396 8470 -7344
rect 8580 -7396 8632 -7344
rect 8644 -7396 8696 -7344
rect 8708 -7396 8760 -7344
rect 8776 -7396 8828 -7344
rect 8840 -7396 8892 -7344
rect 8904 -7396 8956 -7344
rect 8094 -7513 8146 -7483
rect 8158 -7513 8210 -7483
rect 8094 -7535 8117 -7513
rect 8117 -7535 8146 -7513
rect 8158 -7535 8189 -7513
rect 8189 -7535 8210 -7513
rect 8222 -7535 8274 -7483
rect 8290 -7513 8342 -7483
rect 8354 -7513 8406 -7483
rect 8418 -7513 8470 -7483
rect 8290 -7535 8341 -7513
rect 8341 -7535 8342 -7513
rect 8354 -7535 8375 -7513
rect 8375 -7535 8406 -7513
rect 8418 -7535 8447 -7513
rect 8447 -7535 8470 -7513
rect 8580 -7513 8632 -7483
rect 8644 -7513 8696 -7483
rect 8580 -7535 8599 -7513
rect 8599 -7535 8632 -7513
rect 8644 -7535 8671 -7513
rect 8671 -7535 8696 -7513
rect 8708 -7535 8760 -7483
rect 8776 -7535 8828 -7483
rect 8840 -7513 8892 -7483
rect 8840 -7535 8857 -7513
rect 8857 -7535 8891 -7513
rect 8891 -7535 8892 -7513
rect 8904 -7513 8956 -7483
rect 8904 -7535 8929 -7513
rect 8929 -7535 8956 -7513
rect 1624 -7958 1676 -7906
rect 1688 -7958 1740 -7906
rect 1752 -7958 1804 -7906
rect 2141 -7958 2193 -7906
rect 2205 -7958 2257 -7906
rect 2269 -7958 2321 -7906
rect 2593 -8127 2645 -8075
rect 2657 -8127 2709 -8075
rect 2721 -8127 2773 -8075
rect 1364 -8290 1416 -8238
rect 1428 -8290 1480 -8238
rect 1492 -8290 1544 -8238
rect 1882 -8290 1934 -8238
rect 1946 -8290 1998 -8238
rect 2010 -8290 2062 -8238
rect 2398 -8290 2450 -8238
rect 2462 -8290 2514 -8238
rect 2526 -8290 2578 -8238
rect 3110 -8127 3162 -8075
rect 3174 -8127 3226 -8075
rect 3238 -8127 3290 -8075
rect 3818 -7958 3870 -7906
rect 3882 -7958 3934 -7906
rect 3946 -7958 3998 -7906
rect 4335 -7958 4387 -7906
rect 4399 -7958 4451 -7906
rect 4463 -7958 4515 -7906
rect 3559 -8290 3611 -8238
rect 3623 -8290 3675 -8238
rect 3687 -8290 3739 -8238
rect 4076 -8290 4128 -8238
rect 4140 -8290 4192 -8238
rect 4204 -8290 4256 -8238
rect 4591 -8290 4643 -8238
rect 4655 -8290 4707 -8238
rect 4719 -8290 4771 -8238
rect 5980 -7958 6032 -7906
rect 6044 -7958 6096 -7906
rect 6108 -7958 6160 -7906
rect 6497 -7958 6549 -7906
rect 6561 -7958 6613 -7906
rect 6625 -7958 6677 -7906
rect 5724 -8290 5776 -8238
rect 5788 -8290 5840 -8238
rect 5852 -8290 5904 -8238
rect 6239 -8290 6291 -8238
rect 6303 -8290 6355 -8238
rect 6367 -8290 6419 -8238
rect 6756 -8290 6808 -8238
rect 6820 -8290 6872 -8238
rect 6884 -8290 6936 -8238
rect 2850 -8458 2902 -8406
rect 2914 -8458 2966 -8406
rect 2978 -8458 3030 -8406
rect 3368 -8458 3420 -8406
rect 3432 -8458 3484 -8406
rect 3496 -8458 3548 -8406
rect 7205 -8127 7257 -8075
rect 7269 -8127 7321 -8075
rect 7333 -8127 7385 -8075
rect 7722 -8127 7774 -8075
rect 7786 -8127 7838 -8075
rect 7850 -8127 7902 -8075
rect 8174 -7958 8226 -7906
rect 8238 -7958 8290 -7906
rect 8302 -7958 8354 -7906
rect 8692 -7958 8744 -7906
rect 8756 -7958 8808 -7906
rect 8820 -7958 8872 -7906
rect 7917 -8290 7969 -8238
rect 7981 -8290 8033 -8238
rect 8045 -8290 8097 -8238
rect 8434 -8290 8486 -8238
rect 8498 -8290 8550 -8238
rect 8562 -8290 8614 -8238
rect 8951 -8290 9003 -8238
rect 9015 -8290 9067 -8238
rect 9079 -8290 9131 -8238
rect 6948 -8458 7000 -8406
rect 7012 -8458 7064 -8406
rect 7076 -8458 7128 -8406
rect 7465 -8458 7517 -8406
rect 7529 -8458 7581 -8406
rect 7593 -8458 7645 -8406
<< metal2 >>
rect 2843 297 7652 319
rect 2843 281 5001 297
rect 2843 229 2850 281
rect 2902 229 2914 281
rect 2966 229 2978 281
rect 3030 229 3368 281
rect 3420 229 3432 281
rect 3484 229 3496 281
rect 3548 241 5001 281
rect 5057 241 5081 297
rect 5137 241 5161 297
rect 5217 241 5278 297
rect 5334 241 5358 297
rect 5414 241 5438 297
rect 5494 281 7652 297
rect 5494 241 6948 281
rect 3548 229 6948 241
rect 7000 229 7012 281
rect 7064 229 7076 281
rect 7128 229 7465 281
rect 7517 229 7529 281
rect 7581 229 7593 281
rect 7645 229 7652 281
rect 2843 219 7652 229
rect 892 128 9603 150
rect 892 72 932 128
rect 988 72 1012 128
rect 1068 72 1092 128
rect 1148 112 9347 128
rect 1148 72 1364 112
rect 892 60 1364 72
rect 1416 60 1428 112
rect 1480 60 1492 112
rect 1544 60 1882 112
rect 1934 60 1946 112
rect 1998 60 2010 112
rect 2062 60 2398 112
rect 2450 60 2462 112
rect 2514 60 2526 112
rect 2578 60 3559 112
rect 3611 60 3623 112
rect 3675 60 3687 112
rect 3739 60 4076 112
rect 4128 60 4140 112
rect 4192 60 4204 112
rect 4256 60 4591 112
rect 4643 60 4655 112
rect 4707 60 4719 112
rect 4771 60 5724 112
rect 5776 60 5788 112
rect 5840 60 5852 112
rect 5904 60 6239 112
rect 6291 60 6303 112
rect 6355 60 6367 112
rect 6419 60 6756 112
rect 6808 60 6820 112
rect 6872 60 6884 112
rect 6936 60 7917 112
rect 7969 60 7981 112
rect 8033 60 8045 112
rect 8097 60 8434 112
rect 8486 60 8498 112
rect 8550 60 8562 112
rect 8614 60 8951 112
rect 9003 60 9015 112
rect 9067 60 9079 112
rect 9131 72 9347 112
rect 9403 72 9427 128
rect 9483 72 9507 128
rect 9563 72 9603 128
rect 9131 60 9603 72
rect 892 50 9603 60
rect 2586 -35 7909 -13
rect 2586 -51 4566 -35
rect 2586 -103 2593 -51
rect 2645 -103 2657 -51
rect 2709 -103 2721 -51
rect 2773 -103 3110 -51
rect 3162 -103 3174 -51
rect 3226 -103 3238 -51
rect 3290 -91 4566 -51
rect 4622 -91 4646 -35
rect 4702 -91 4726 -35
rect 4782 -91 5713 -35
rect 5769 -91 5793 -35
rect 5849 -91 5873 -35
rect 5929 -51 7909 -35
rect 5929 -91 7205 -51
rect 3290 -103 7205 -91
rect 7257 -103 7269 -51
rect 7321 -103 7333 -51
rect 7385 -103 7722 -51
rect 7774 -103 7786 -51
rect 7838 -103 7850 -51
rect 7902 -103 7909 -51
rect 2586 -113 7909 -103
rect 1315 -203 9181 -181
rect 1315 -259 1355 -203
rect 1411 -259 1435 -203
rect 1491 -259 1515 -203
rect 1571 -219 8925 -203
rect 1571 -259 1624 -219
rect 1315 -271 1624 -259
rect 1676 -271 1688 -219
rect 1740 -271 1752 -219
rect 1804 -271 2141 -219
rect 2193 -271 2205 -219
rect 2257 -271 2269 -219
rect 2321 -271 3818 -219
rect 3870 -271 3882 -219
rect 3934 -271 3946 -219
rect 3998 -271 4335 -219
rect 4387 -271 4399 -219
rect 4451 -271 4463 -219
rect 4515 -271 5980 -219
rect 6032 -271 6044 -219
rect 6096 -271 6108 -219
rect 6160 -271 6497 -219
rect 6549 -271 6561 -219
rect 6613 -271 6625 -219
rect 6677 -271 8174 -219
rect 8226 -271 8238 -219
rect 8290 -271 8302 -219
rect 8354 -271 8692 -219
rect 8744 -271 8756 -219
rect 8808 -271 8820 -219
rect 8872 -259 8925 -219
rect 8981 -259 9005 -203
rect 9061 -259 9085 -203
rect 9141 -259 9181 -203
rect 8872 -271 9181 -259
rect 1315 -281 9181 -271
rect 2441 -624 2741 -613
rect 7754 -624 8054 -613
rect 1489 -635 9006 -624
rect 1489 -643 2481 -635
rect 1489 -695 1539 -643
rect 1591 -695 1603 -643
rect 1655 -695 1667 -643
rect 1719 -695 1735 -643
rect 1787 -695 1799 -643
rect 1851 -695 1863 -643
rect 1915 -695 2025 -643
rect 2077 -695 2089 -643
rect 2141 -695 2153 -643
rect 2205 -695 2221 -643
rect 2273 -695 2285 -643
rect 2337 -695 2349 -643
rect 2401 -691 2481 -643
rect 2537 -691 2561 -635
rect 2617 -691 2641 -635
rect 2697 -643 7798 -635
rect 2697 -691 3737 -643
rect 2401 -695 3737 -691
rect 3789 -695 3801 -643
rect 3853 -695 3865 -643
rect 3917 -695 3933 -643
rect 3985 -695 3997 -643
rect 4049 -695 4061 -643
rect 4113 -695 4223 -643
rect 4275 -695 4287 -643
rect 4339 -695 4351 -643
rect 4403 -695 4419 -643
rect 4471 -695 4483 -643
rect 4535 -695 4547 -643
rect 4599 -695 5896 -643
rect 5948 -695 5960 -643
rect 6012 -695 6024 -643
rect 6076 -695 6092 -643
rect 6144 -695 6156 -643
rect 6208 -695 6220 -643
rect 6272 -695 6382 -643
rect 6434 -695 6446 -643
rect 6498 -695 6510 -643
rect 6562 -695 6578 -643
rect 6630 -695 6642 -643
rect 6694 -695 6706 -643
rect 6758 -691 7798 -643
rect 7854 -691 7878 -635
rect 7934 -691 7958 -635
rect 8014 -643 9006 -635
rect 8014 -691 8094 -643
rect 6758 -695 8094 -691
rect 8146 -695 8158 -643
rect 8210 -695 8222 -643
rect 8274 -695 8290 -643
rect 8342 -695 8354 -643
rect 8406 -695 8418 -643
rect 8470 -695 8580 -643
rect 8632 -695 8644 -643
rect 8696 -695 8708 -643
rect 8760 -695 8776 -643
rect 8828 -695 8840 -643
rect 8892 -695 8904 -643
rect 8956 -695 9006 -643
rect 1489 -713 9006 -695
rect 1489 -781 9006 -763
rect 1489 -833 1539 -781
rect 1591 -833 1603 -781
rect 1655 -833 1667 -781
rect 1719 -833 1735 -781
rect 1787 -833 1799 -781
rect 1851 -833 1863 -781
rect 1915 -833 2025 -781
rect 2077 -833 2089 -781
rect 2141 -833 2153 -781
rect 2205 -833 2221 -781
rect 2273 -833 2285 -781
rect 2337 -833 2349 -781
rect 2401 -833 2749 -781
rect 2801 -833 2813 -781
rect 2865 -833 2877 -781
rect 2929 -833 2945 -781
rect 2997 -833 3009 -781
rect 3061 -833 3073 -781
rect 3125 -833 3137 -781
rect 3189 -833 3205 -781
rect 3257 -833 3269 -781
rect 3321 -833 3333 -781
rect 3385 -833 3737 -781
rect 3789 -833 3801 -781
rect 3853 -833 3865 -781
rect 3917 -833 3933 -781
rect 3985 -833 3997 -781
rect 4049 -833 4061 -781
rect 4113 -833 4223 -781
rect 4275 -833 4287 -781
rect 4339 -833 4351 -781
rect 4403 -833 4419 -781
rect 4471 -833 4483 -781
rect 4535 -833 4547 -781
rect 4599 -833 5896 -781
rect 5948 -833 5960 -781
rect 6012 -833 6024 -781
rect 6076 -833 6092 -781
rect 6144 -833 6156 -781
rect 6208 -833 6220 -781
rect 6272 -833 6382 -781
rect 6434 -833 6446 -781
rect 6498 -833 6510 -781
rect 6562 -833 6578 -781
rect 6630 -833 6642 -781
rect 6694 -833 6706 -781
rect 6758 -833 7110 -781
rect 7162 -833 7174 -781
rect 7226 -833 7238 -781
rect 7290 -833 7306 -781
rect 7358 -833 7370 -781
rect 7422 -833 7434 -781
rect 7486 -833 7498 -781
rect 7550 -833 7566 -781
rect 7618 -833 7630 -781
rect 7682 -833 7694 -781
rect 7746 -833 8094 -781
rect 8146 -833 8158 -781
rect 8210 -833 8222 -781
rect 8274 -833 8290 -781
rect 8342 -833 8354 -781
rect 8406 -833 8418 -781
rect 8470 -833 8580 -781
rect 8632 -833 8644 -781
rect 8696 -833 8708 -781
rect 8760 -833 8776 -781
rect 8828 -833 8840 -781
rect 8892 -833 8904 -781
rect 8956 -833 9006 -781
rect 1489 -851 9006 -833
rect 3409 -945 3709 -933
rect 6786 -945 7086 -933
rect 1489 -955 9006 -945
rect 1489 -959 3449 -955
rect 1489 -1011 1539 -959
rect 1591 -1011 1603 -959
rect 1655 -1011 1667 -959
rect 1719 -1011 1735 -959
rect 1787 -1011 1799 -959
rect 1851 -1011 1863 -959
rect 1915 -1011 2025 -959
rect 2077 -1011 2089 -959
rect 2141 -1011 2153 -959
rect 2205 -1011 2221 -959
rect 2273 -1011 2285 -959
rect 2337 -1011 2349 -959
rect 2401 -1011 3449 -959
rect 3505 -1011 3529 -955
rect 3585 -1011 3609 -955
rect 3665 -959 6830 -955
rect 3665 -1011 3737 -959
rect 3789 -1011 3801 -959
rect 3853 -1011 3865 -959
rect 3917 -1011 3933 -959
rect 3985 -1011 3997 -959
rect 4049 -1011 4061 -959
rect 4113 -1011 4223 -959
rect 4275 -1011 4287 -959
rect 4339 -1011 4351 -959
rect 4403 -1011 4419 -959
rect 4471 -1011 4483 -959
rect 4535 -1011 4547 -959
rect 4599 -1011 5896 -959
rect 5948 -1011 5960 -959
rect 6012 -1011 6024 -959
rect 6076 -1011 6092 -959
rect 6144 -1011 6156 -959
rect 6208 -1011 6220 -959
rect 6272 -1011 6382 -959
rect 6434 -1011 6446 -959
rect 6498 -1011 6510 -959
rect 6562 -1011 6578 -959
rect 6630 -1011 6642 -959
rect 6694 -1011 6706 -959
rect 6758 -1011 6830 -959
rect 6886 -1011 6910 -955
rect 6966 -1011 6990 -955
rect 7046 -959 9006 -955
rect 7046 -1011 8094 -959
rect 8146 -1011 8158 -959
rect 8210 -1011 8222 -959
rect 8274 -1011 8290 -959
rect 8342 -1011 8354 -959
rect 8406 -1011 8418 -959
rect 8470 -1011 8580 -959
rect 8632 -1011 8644 -959
rect 8696 -1011 8708 -959
rect 8760 -1011 8776 -959
rect 8828 -1011 8840 -959
rect 8892 -1011 8904 -959
rect 8956 -1011 9006 -959
rect 1489 -1033 9006 -1011
rect 1360 -1393 9136 -1371
rect 1360 -1409 5001 -1393
rect 1360 -1461 1367 -1409
rect 1419 -1461 1431 -1409
rect 1483 -1461 1495 -1409
rect 1547 -1461 1882 -1409
rect 1934 -1461 1946 -1409
rect 1998 -1461 2010 -1409
rect 2062 -1461 2399 -1409
rect 2451 -1461 2463 -1409
rect 2515 -1461 2527 -1409
rect 2579 -1461 3559 -1409
rect 3611 -1461 3623 -1409
rect 3675 -1461 3687 -1409
rect 3739 -1461 4076 -1409
rect 4128 -1461 4140 -1409
rect 4192 -1461 4204 -1409
rect 4256 -1461 4593 -1409
rect 4645 -1461 4657 -1409
rect 4709 -1461 4721 -1409
rect 4773 -1449 5001 -1409
rect 5057 -1449 5081 -1393
rect 5137 -1449 5161 -1393
rect 5217 -1449 5278 -1393
rect 5334 -1449 5358 -1393
rect 5414 -1449 5438 -1393
rect 5494 -1409 9136 -1393
rect 5494 -1449 5722 -1409
rect 4773 -1461 5722 -1449
rect 5774 -1461 5786 -1409
rect 5838 -1461 5850 -1409
rect 5902 -1461 6239 -1409
rect 6291 -1461 6303 -1409
rect 6355 -1461 6367 -1409
rect 6419 -1461 6756 -1409
rect 6808 -1461 6820 -1409
rect 6872 -1461 6884 -1409
rect 6936 -1461 7916 -1409
rect 7968 -1461 7980 -1409
rect 8032 -1461 8044 -1409
rect 8096 -1461 8434 -1409
rect 8486 -1461 8498 -1409
rect 8550 -1461 8562 -1409
rect 8614 -1461 8949 -1409
rect 9001 -1461 9013 -1409
rect 9065 -1461 9077 -1409
rect 9129 -1461 9136 -1409
rect 1360 -1471 9136 -1461
rect 1315 -1533 9181 -1511
rect 1315 -1589 1355 -1533
rect 1411 -1589 1435 -1533
rect 1491 -1589 1515 -1533
rect 1571 -1549 8925 -1533
rect 1571 -1589 2849 -1549
rect 1315 -1601 2849 -1589
rect 2901 -1601 2913 -1549
rect 2965 -1601 2977 -1549
rect 3029 -1601 3366 -1549
rect 3418 -1601 3430 -1549
rect 3482 -1601 3494 -1549
rect 3546 -1601 6949 -1549
rect 7001 -1601 7013 -1549
rect 7065 -1601 7077 -1549
rect 7129 -1601 7466 -1549
rect 7518 -1601 7530 -1549
rect 7582 -1601 7594 -1549
rect 7646 -1589 8925 -1549
rect 8981 -1589 9005 -1533
rect 9061 -1589 9085 -1533
rect 9141 -1589 9181 -1533
rect 7646 -1601 9181 -1589
rect 1315 -1611 9181 -1601
rect 1618 -1694 8878 -1672
rect 1618 -1710 4566 -1694
rect 1618 -1762 1625 -1710
rect 1677 -1762 1689 -1710
rect 1741 -1762 1753 -1710
rect 1805 -1762 2142 -1710
rect 2194 -1762 2206 -1710
rect 2258 -1762 2270 -1710
rect 2322 -1762 3819 -1710
rect 3871 -1762 3883 -1710
rect 3935 -1762 3947 -1710
rect 3999 -1762 4336 -1710
rect 4388 -1762 4400 -1710
rect 4452 -1762 4464 -1710
rect 4516 -1750 4566 -1710
rect 4622 -1750 4646 -1694
rect 4702 -1750 4726 -1694
rect 4782 -1750 5713 -1694
rect 5769 -1750 5793 -1694
rect 5849 -1750 5873 -1694
rect 5929 -1710 8878 -1694
rect 5929 -1750 5979 -1710
rect 4516 -1762 5979 -1750
rect 6031 -1762 6043 -1710
rect 6095 -1762 6107 -1710
rect 6159 -1762 6496 -1710
rect 6548 -1762 6560 -1710
rect 6612 -1762 6624 -1710
rect 6676 -1762 8173 -1710
rect 8225 -1762 8237 -1710
rect 8289 -1762 8301 -1710
rect 8353 -1762 8691 -1710
rect 8743 -1762 8755 -1710
rect 8807 -1762 8819 -1710
rect 8871 -1762 8878 -1710
rect 1618 -1772 8878 -1762
rect 881 -1838 9614 -1816
rect 881 -1894 932 -1838
rect 988 -1894 1012 -1838
rect 1068 -1894 1092 -1838
rect 1148 -1854 9347 -1838
rect 1148 -1894 2591 -1854
rect 881 -1906 2591 -1894
rect 2643 -1906 2655 -1854
rect 2707 -1906 2719 -1854
rect 2771 -1906 3108 -1854
rect 3160 -1906 3172 -1854
rect 3224 -1906 3236 -1854
rect 3288 -1906 7207 -1854
rect 7259 -1906 7271 -1854
rect 7323 -1906 7335 -1854
rect 7387 -1906 7724 -1854
rect 7776 -1906 7788 -1854
rect 7840 -1906 7852 -1854
rect 7904 -1894 9347 -1854
rect 9403 -1894 9427 -1838
rect 9483 -1894 9507 -1838
rect 9563 -1894 9614 -1838
rect 7904 -1906 9614 -1894
rect 881 -1916 9614 -1906
rect 3409 -2271 3709 -2260
rect 1489 -2282 9006 -2271
rect 1489 -2290 3449 -2282
rect 1489 -2342 1539 -2290
rect 1591 -2342 1603 -2290
rect 1655 -2342 1667 -2290
rect 1719 -2342 1735 -2290
rect 1787 -2342 1799 -2290
rect 1851 -2342 1863 -2290
rect 1915 -2342 2025 -2290
rect 2077 -2342 2089 -2290
rect 2141 -2342 2153 -2290
rect 2205 -2342 2221 -2290
rect 2273 -2342 2285 -2290
rect 2337 -2342 2349 -2290
rect 2401 -2338 3449 -2290
rect 3505 -2338 3529 -2282
rect 3585 -2338 3609 -2282
rect 3665 -2290 9006 -2282
rect 3665 -2338 3737 -2290
rect 2401 -2342 3737 -2338
rect 3789 -2342 3801 -2290
rect 3853 -2342 3865 -2290
rect 3917 -2342 3933 -2290
rect 3985 -2342 3997 -2290
rect 4049 -2342 4061 -2290
rect 4113 -2342 4223 -2290
rect 4275 -2342 4287 -2290
rect 4339 -2342 4351 -2290
rect 4403 -2342 4419 -2290
rect 4471 -2342 4483 -2290
rect 4535 -2342 4547 -2290
rect 4599 -2342 5896 -2290
rect 5948 -2342 5960 -2290
rect 6012 -2342 6024 -2290
rect 6076 -2342 6092 -2290
rect 6144 -2342 6156 -2290
rect 6208 -2342 6220 -2290
rect 6272 -2342 6382 -2290
rect 6434 -2342 6446 -2290
rect 6498 -2342 6510 -2290
rect 6562 -2342 6578 -2290
rect 6630 -2342 6642 -2290
rect 6694 -2342 6706 -2290
rect 6758 -2293 8094 -2290
rect 6758 -2342 6830 -2293
rect 1489 -2349 6830 -2342
rect 6886 -2349 6910 -2293
rect 6966 -2349 6990 -2293
rect 7046 -2342 8094 -2293
rect 8146 -2342 8158 -2290
rect 8210 -2342 8222 -2290
rect 8274 -2342 8290 -2290
rect 8342 -2342 8354 -2290
rect 8406 -2342 8418 -2290
rect 8470 -2342 8580 -2290
rect 8632 -2342 8644 -2290
rect 8696 -2342 8708 -2290
rect 8760 -2342 8776 -2290
rect 8828 -2342 8840 -2290
rect 8892 -2342 8904 -2290
rect 8956 -2342 9006 -2290
rect 7046 -2349 9006 -2342
rect 1489 -2360 9006 -2349
rect 6786 -2371 7086 -2360
rect 1489 -2428 9006 -2410
rect 1489 -2480 1539 -2428
rect 1591 -2480 1603 -2428
rect 1655 -2480 1667 -2428
rect 1719 -2480 1735 -2428
rect 1787 -2480 1799 -2428
rect 1851 -2480 1863 -2428
rect 1915 -2480 2025 -2428
rect 2077 -2480 2089 -2428
rect 2141 -2480 2153 -2428
rect 2205 -2480 2221 -2428
rect 2273 -2480 2285 -2428
rect 2337 -2480 2349 -2428
rect 2401 -2480 2749 -2428
rect 2801 -2480 2813 -2428
rect 2865 -2480 2877 -2428
rect 2929 -2480 2945 -2428
rect 2997 -2480 3009 -2428
rect 3061 -2480 3073 -2428
rect 3125 -2480 3137 -2428
rect 3189 -2480 3205 -2428
rect 3257 -2480 3269 -2428
rect 3321 -2480 3333 -2428
rect 3385 -2480 3737 -2428
rect 3789 -2480 3801 -2428
rect 3853 -2480 3865 -2428
rect 3917 -2480 3933 -2428
rect 3985 -2480 3997 -2428
rect 4049 -2480 4061 -2428
rect 4113 -2480 4223 -2428
rect 4275 -2480 4287 -2428
rect 4339 -2480 4351 -2428
rect 4403 -2480 4419 -2428
rect 4471 -2480 4483 -2428
rect 4535 -2480 4547 -2428
rect 4599 -2480 5896 -2428
rect 5948 -2480 5960 -2428
rect 6012 -2480 6024 -2428
rect 6076 -2480 6092 -2428
rect 6144 -2480 6156 -2428
rect 6208 -2480 6220 -2428
rect 6272 -2480 6382 -2428
rect 6434 -2480 6446 -2428
rect 6498 -2480 6510 -2428
rect 6562 -2480 6578 -2428
rect 6630 -2480 6642 -2428
rect 6694 -2480 6706 -2428
rect 6758 -2480 7110 -2428
rect 7162 -2480 7174 -2428
rect 7226 -2480 7238 -2428
rect 7290 -2480 7306 -2428
rect 7358 -2480 7370 -2428
rect 7422 -2480 7434 -2428
rect 7486 -2480 7498 -2428
rect 7550 -2480 7566 -2428
rect 7618 -2480 7630 -2428
rect 7682 -2480 7694 -2428
rect 7746 -2480 8094 -2428
rect 8146 -2480 8158 -2428
rect 8210 -2480 8222 -2428
rect 8274 -2480 8290 -2428
rect 8342 -2480 8354 -2428
rect 8406 -2480 8418 -2428
rect 8470 -2480 8580 -2428
rect 8632 -2480 8644 -2428
rect 8696 -2480 8708 -2428
rect 8760 -2480 8776 -2428
rect 8828 -2480 8840 -2428
rect 8892 -2480 8904 -2428
rect 8956 -2480 9006 -2428
rect 1489 -2498 9006 -2480
rect 1489 -2606 9006 -2592
rect 1489 -2658 1539 -2606
rect 1591 -2658 1603 -2606
rect 1655 -2658 1667 -2606
rect 1719 -2658 1735 -2606
rect 1787 -2658 1799 -2606
rect 1851 -2658 1863 -2606
rect 1915 -2658 2025 -2606
rect 2077 -2658 2089 -2606
rect 2141 -2658 2153 -2606
rect 2205 -2658 2221 -2606
rect 2273 -2658 2285 -2606
rect 2337 -2658 2349 -2606
rect 2401 -2614 3737 -2606
rect 2401 -2658 2481 -2614
rect 1489 -2670 2481 -2658
rect 2537 -2670 2561 -2614
rect 2617 -2670 2641 -2614
rect 2697 -2658 3737 -2614
rect 3789 -2658 3801 -2606
rect 3853 -2658 3865 -2606
rect 3917 -2658 3933 -2606
rect 3985 -2658 3997 -2606
rect 4049 -2658 4061 -2606
rect 4113 -2658 4223 -2606
rect 4275 -2658 4287 -2606
rect 4339 -2658 4351 -2606
rect 4403 -2658 4419 -2606
rect 4471 -2658 4483 -2606
rect 4535 -2658 4547 -2606
rect 4599 -2658 5896 -2606
rect 5948 -2658 5960 -2606
rect 6012 -2658 6024 -2606
rect 6076 -2658 6092 -2606
rect 6144 -2658 6156 -2606
rect 6208 -2658 6220 -2606
rect 6272 -2658 6382 -2606
rect 6434 -2658 6446 -2606
rect 6498 -2658 6510 -2606
rect 6562 -2658 6578 -2606
rect 6630 -2658 6642 -2606
rect 6694 -2658 6706 -2606
rect 6758 -2614 8094 -2606
rect 6758 -2658 7798 -2614
rect 2697 -2670 7798 -2658
rect 7854 -2670 7878 -2614
rect 7934 -2670 7958 -2614
rect 8014 -2658 8094 -2614
rect 8146 -2658 8158 -2606
rect 8210 -2658 8222 -2606
rect 8274 -2658 8290 -2606
rect 8342 -2658 8354 -2606
rect 8406 -2658 8418 -2606
rect 8470 -2658 8580 -2606
rect 8632 -2658 8644 -2606
rect 8696 -2658 8708 -2606
rect 8760 -2658 8776 -2606
rect 8828 -2658 8840 -2606
rect 8892 -2658 8904 -2606
rect 8956 -2658 9006 -2606
rect 8014 -2670 9006 -2658
rect 1489 -2680 9006 -2670
rect 2441 -2692 2741 -2680
rect 7754 -2692 8054 -2680
rect 1315 -3033 9181 -3023
rect 1315 -3045 1624 -3033
rect 1315 -3101 1355 -3045
rect 1411 -3101 1435 -3045
rect 1491 -3101 1515 -3045
rect 1571 -3085 1624 -3045
rect 1676 -3085 1688 -3033
rect 1740 -3085 1752 -3033
rect 1804 -3085 2141 -3033
rect 2193 -3085 2205 -3033
rect 2257 -3085 2269 -3033
rect 2321 -3085 3818 -3033
rect 3870 -3085 3882 -3033
rect 3934 -3085 3946 -3033
rect 3998 -3085 4335 -3033
rect 4387 -3085 4399 -3033
rect 4451 -3085 4463 -3033
rect 4515 -3085 5980 -3033
rect 6032 -3085 6044 -3033
rect 6096 -3085 6108 -3033
rect 6160 -3085 6497 -3033
rect 6549 -3085 6561 -3033
rect 6613 -3085 6625 -3033
rect 6677 -3085 8174 -3033
rect 8226 -3085 8238 -3033
rect 8290 -3085 8302 -3033
rect 8354 -3085 8692 -3033
rect 8744 -3085 8756 -3033
rect 8808 -3085 8820 -3033
rect 8872 -3045 9181 -3033
rect 8872 -3085 8925 -3045
rect 1571 -3101 8925 -3085
rect 8981 -3101 9005 -3045
rect 9061 -3101 9085 -3045
rect 9141 -3101 9181 -3045
rect 1315 -3123 9181 -3101
rect 2586 -3202 7909 -3192
rect 2586 -3254 2593 -3202
rect 2645 -3254 2657 -3202
rect 2709 -3254 2721 -3202
rect 2773 -3254 3110 -3202
rect 3162 -3254 3174 -3202
rect 3226 -3254 3238 -3202
rect 3290 -3214 7205 -3202
rect 3290 -3254 4566 -3214
rect 2586 -3270 4566 -3254
rect 4622 -3270 4646 -3214
rect 4702 -3270 4726 -3214
rect 4782 -3270 5713 -3214
rect 5769 -3270 5793 -3214
rect 5849 -3270 5873 -3214
rect 5929 -3254 7205 -3214
rect 7257 -3254 7269 -3202
rect 7321 -3254 7333 -3202
rect 7385 -3254 7722 -3202
rect 7774 -3254 7786 -3202
rect 7838 -3254 7850 -3202
rect 7902 -3254 7909 -3202
rect 5929 -3270 7909 -3254
rect 2586 -3292 7909 -3270
rect 892 -3364 9603 -3354
rect 892 -3376 1364 -3364
rect 892 -3432 932 -3376
rect 988 -3432 1012 -3376
rect 1068 -3432 1092 -3376
rect 1148 -3416 1364 -3376
rect 1416 -3416 1428 -3364
rect 1480 -3416 1492 -3364
rect 1544 -3416 1882 -3364
rect 1934 -3416 1946 -3364
rect 1998 -3416 2010 -3364
rect 2062 -3416 2398 -3364
rect 2450 -3416 2462 -3364
rect 2514 -3416 2526 -3364
rect 2578 -3416 3559 -3364
rect 3611 -3416 3623 -3364
rect 3675 -3416 3687 -3364
rect 3739 -3416 4076 -3364
rect 4128 -3416 4140 -3364
rect 4192 -3416 4204 -3364
rect 4256 -3416 4591 -3364
rect 4643 -3416 4655 -3364
rect 4707 -3416 4719 -3364
rect 4771 -3416 5724 -3364
rect 5776 -3416 5788 -3364
rect 5840 -3416 5852 -3364
rect 5904 -3416 6239 -3364
rect 6291 -3416 6303 -3364
rect 6355 -3416 6367 -3364
rect 6419 -3416 6756 -3364
rect 6808 -3416 6820 -3364
rect 6872 -3416 6884 -3364
rect 6936 -3416 7917 -3364
rect 7969 -3416 7981 -3364
rect 8033 -3416 8045 -3364
rect 8097 -3416 8434 -3364
rect 8486 -3416 8498 -3364
rect 8550 -3416 8562 -3364
rect 8614 -3416 8951 -3364
rect 9003 -3416 9015 -3364
rect 9067 -3416 9079 -3364
rect 9131 -3376 9603 -3364
rect 9131 -3416 9347 -3376
rect 1148 -3432 9347 -3416
rect 9403 -3432 9427 -3376
rect 9483 -3432 9507 -3376
rect 9563 -3432 9603 -3376
rect 892 -3454 9603 -3432
rect 2843 -3533 7652 -3523
rect 2843 -3585 2850 -3533
rect 2902 -3585 2914 -3533
rect 2966 -3585 2978 -3533
rect 3030 -3585 3368 -3533
rect 3420 -3585 3432 -3533
rect 3484 -3585 3496 -3533
rect 3548 -3545 6948 -3533
rect 3548 -3585 5001 -3545
rect 2843 -3601 5001 -3585
rect 5057 -3601 5081 -3545
rect 5137 -3601 5161 -3545
rect 5217 -3601 5278 -3545
rect 5334 -3601 5358 -3545
rect 5414 -3601 5438 -3545
rect 5494 -3585 6948 -3545
rect 7000 -3585 7012 -3533
rect 7064 -3585 7076 -3533
rect 7128 -3585 7465 -3533
rect 7517 -3585 7529 -3533
rect 7581 -3585 7593 -3533
rect 7645 -3585 7652 -3533
rect 5494 -3601 7652 -3585
rect 2843 -3623 7652 -3601
rect 2843 -4576 7652 -4554
rect 2843 -4592 5001 -4576
rect 2843 -4644 2850 -4592
rect 2902 -4644 2914 -4592
rect 2966 -4644 2978 -4592
rect 3030 -4644 3368 -4592
rect 3420 -4644 3432 -4592
rect 3484 -4644 3496 -4592
rect 3548 -4632 5001 -4592
rect 5057 -4632 5081 -4576
rect 5137 -4632 5161 -4576
rect 5217 -4632 5278 -4576
rect 5334 -4632 5358 -4576
rect 5414 -4632 5438 -4576
rect 5494 -4592 7652 -4576
rect 5494 -4632 6948 -4592
rect 3548 -4644 6948 -4632
rect 7000 -4644 7012 -4592
rect 7064 -4644 7076 -4592
rect 7128 -4644 7465 -4592
rect 7517 -4644 7529 -4592
rect 7581 -4644 7593 -4592
rect 7645 -4644 7652 -4592
rect 2843 -4654 7652 -4644
rect 892 -4745 9603 -4723
rect 892 -4801 932 -4745
rect 988 -4801 1012 -4745
rect 1068 -4801 1092 -4745
rect 1148 -4761 9347 -4745
rect 1148 -4801 1364 -4761
rect 892 -4813 1364 -4801
rect 1416 -4813 1428 -4761
rect 1480 -4813 1492 -4761
rect 1544 -4813 1882 -4761
rect 1934 -4813 1946 -4761
rect 1998 -4813 2010 -4761
rect 2062 -4813 2398 -4761
rect 2450 -4813 2462 -4761
rect 2514 -4813 2526 -4761
rect 2578 -4813 3559 -4761
rect 3611 -4813 3623 -4761
rect 3675 -4813 3687 -4761
rect 3739 -4813 4076 -4761
rect 4128 -4813 4140 -4761
rect 4192 -4813 4204 -4761
rect 4256 -4813 4591 -4761
rect 4643 -4813 4655 -4761
rect 4707 -4813 4719 -4761
rect 4771 -4813 5724 -4761
rect 5776 -4813 5788 -4761
rect 5840 -4813 5852 -4761
rect 5904 -4813 6239 -4761
rect 6291 -4813 6303 -4761
rect 6355 -4813 6367 -4761
rect 6419 -4813 6756 -4761
rect 6808 -4813 6820 -4761
rect 6872 -4813 6884 -4761
rect 6936 -4813 7917 -4761
rect 7969 -4813 7981 -4761
rect 8033 -4813 8045 -4761
rect 8097 -4813 8434 -4761
rect 8486 -4813 8498 -4761
rect 8550 -4813 8562 -4761
rect 8614 -4813 8951 -4761
rect 9003 -4813 9015 -4761
rect 9067 -4813 9079 -4761
rect 9131 -4801 9347 -4761
rect 9403 -4801 9427 -4745
rect 9483 -4801 9507 -4745
rect 9563 -4801 9603 -4745
rect 9131 -4813 9603 -4801
rect 892 -4823 9603 -4813
rect 2586 -4908 7909 -4886
rect 2586 -4924 4566 -4908
rect 2586 -4976 2593 -4924
rect 2645 -4976 2657 -4924
rect 2709 -4976 2721 -4924
rect 2773 -4976 3110 -4924
rect 3162 -4976 3174 -4924
rect 3226 -4976 3238 -4924
rect 3290 -4964 4566 -4924
rect 4622 -4964 4646 -4908
rect 4702 -4964 4726 -4908
rect 4782 -4964 5713 -4908
rect 5769 -4964 5793 -4908
rect 5849 -4964 5873 -4908
rect 5929 -4924 7909 -4908
rect 5929 -4964 7205 -4924
rect 3290 -4976 7205 -4964
rect 7257 -4976 7269 -4924
rect 7321 -4976 7333 -4924
rect 7385 -4976 7722 -4924
rect 7774 -4976 7786 -4924
rect 7838 -4976 7850 -4924
rect 7902 -4976 7909 -4924
rect 2586 -4986 7909 -4976
rect 1315 -5077 9181 -5055
rect 1315 -5133 1355 -5077
rect 1411 -5133 1435 -5077
rect 1491 -5133 1515 -5077
rect 1571 -5093 8925 -5077
rect 1571 -5133 1624 -5093
rect 1315 -5145 1624 -5133
rect 1676 -5145 1688 -5093
rect 1740 -5145 1752 -5093
rect 1804 -5145 2141 -5093
rect 2193 -5145 2205 -5093
rect 2257 -5145 2269 -5093
rect 2321 -5145 3818 -5093
rect 3870 -5145 3882 -5093
rect 3934 -5145 3946 -5093
rect 3998 -5145 4335 -5093
rect 4387 -5145 4399 -5093
rect 4451 -5145 4463 -5093
rect 4515 -5145 5980 -5093
rect 6032 -5145 6044 -5093
rect 6096 -5145 6108 -5093
rect 6160 -5145 6497 -5093
rect 6549 -5145 6561 -5093
rect 6613 -5145 6625 -5093
rect 6677 -5145 8174 -5093
rect 8226 -5145 8238 -5093
rect 8290 -5145 8302 -5093
rect 8354 -5145 8692 -5093
rect 8744 -5145 8756 -5093
rect 8808 -5145 8820 -5093
rect 8872 -5133 8925 -5093
rect 8981 -5133 9005 -5077
rect 9061 -5133 9085 -5077
rect 9141 -5133 9181 -5077
rect 8872 -5145 9181 -5133
rect 1315 -5155 9181 -5145
rect 2441 -5498 2741 -5486
rect 7754 -5498 8054 -5486
rect 1489 -5508 9006 -5498
rect 1489 -5519 2481 -5508
rect 1489 -5571 1539 -5519
rect 1591 -5571 1603 -5519
rect 1655 -5571 1667 -5519
rect 1719 -5571 1735 -5519
rect 1787 -5571 1799 -5519
rect 1851 -5571 1863 -5519
rect 1915 -5571 2025 -5519
rect 2077 -5571 2089 -5519
rect 2141 -5571 2153 -5519
rect 2205 -5571 2221 -5519
rect 2273 -5571 2285 -5519
rect 2337 -5571 2349 -5519
rect 2401 -5564 2481 -5519
rect 2537 -5564 2561 -5508
rect 2617 -5564 2641 -5508
rect 2697 -5519 7798 -5508
rect 2697 -5564 3737 -5519
rect 2401 -5571 3737 -5564
rect 3789 -5571 3801 -5519
rect 3853 -5571 3865 -5519
rect 3917 -5571 3933 -5519
rect 3985 -5571 3997 -5519
rect 4049 -5571 4061 -5519
rect 4113 -5571 4223 -5519
rect 4275 -5571 4287 -5519
rect 4339 -5571 4351 -5519
rect 4403 -5571 4419 -5519
rect 4471 -5571 4483 -5519
rect 4535 -5571 4547 -5519
rect 4599 -5571 5896 -5519
rect 5948 -5571 5960 -5519
rect 6012 -5571 6024 -5519
rect 6076 -5571 6092 -5519
rect 6144 -5571 6156 -5519
rect 6208 -5571 6220 -5519
rect 6272 -5571 6382 -5519
rect 6434 -5571 6446 -5519
rect 6498 -5571 6510 -5519
rect 6562 -5571 6578 -5519
rect 6630 -5571 6642 -5519
rect 6694 -5571 6706 -5519
rect 6758 -5564 7798 -5519
rect 7854 -5564 7878 -5508
rect 7934 -5564 7958 -5508
rect 8014 -5519 9006 -5508
rect 8014 -5564 8094 -5519
rect 6758 -5571 8094 -5564
rect 8146 -5571 8158 -5519
rect 8210 -5571 8222 -5519
rect 8274 -5571 8290 -5519
rect 8342 -5571 8354 -5519
rect 8406 -5571 8418 -5519
rect 8470 -5571 8580 -5519
rect 8632 -5571 8644 -5519
rect 8696 -5571 8708 -5519
rect 8760 -5571 8776 -5519
rect 8828 -5571 8840 -5519
rect 8892 -5571 8904 -5519
rect 8956 -5571 9006 -5519
rect 1489 -5586 9006 -5571
rect 1489 -5697 9006 -5680
rect 1489 -5749 1539 -5697
rect 1591 -5749 1603 -5697
rect 1655 -5749 1667 -5697
rect 1719 -5749 1735 -5697
rect 1787 -5749 1799 -5697
rect 1851 -5749 1863 -5697
rect 1915 -5749 2025 -5697
rect 2077 -5749 2089 -5697
rect 2141 -5749 2153 -5697
rect 2205 -5749 2221 -5697
rect 2273 -5749 2285 -5697
rect 2337 -5749 2349 -5697
rect 2401 -5749 2749 -5697
rect 2801 -5749 2813 -5697
rect 2865 -5749 2877 -5697
rect 2929 -5749 2945 -5697
rect 2997 -5749 3009 -5697
rect 3061 -5749 3073 -5697
rect 3125 -5749 3137 -5697
rect 3189 -5749 3205 -5697
rect 3257 -5749 3269 -5697
rect 3321 -5749 3333 -5697
rect 3385 -5749 3737 -5697
rect 3789 -5749 3801 -5697
rect 3853 -5749 3865 -5697
rect 3917 -5749 3933 -5697
rect 3985 -5749 3997 -5697
rect 4049 -5749 4061 -5697
rect 4113 -5749 4223 -5697
rect 4275 -5749 4287 -5697
rect 4339 -5749 4351 -5697
rect 4403 -5749 4419 -5697
rect 4471 -5749 4483 -5697
rect 4535 -5749 4547 -5697
rect 4599 -5749 5896 -5697
rect 5948 -5749 5960 -5697
rect 6012 -5749 6024 -5697
rect 6076 -5749 6092 -5697
rect 6144 -5749 6156 -5697
rect 6208 -5749 6220 -5697
rect 6272 -5749 6382 -5697
rect 6434 -5749 6446 -5697
rect 6498 -5749 6510 -5697
rect 6562 -5749 6578 -5697
rect 6630 -5749 6642 -5697
rect 6694 -5749 6706 -5697
rect 6758 -5749 7110 -5697
rect 7162 -5749 7174 -5697
rect 7226 -5749 7238 -5697
rect 7290 -5749 7306 -5697
rect 7358 -5749 7370 -5697
rect 7422 -5749 7434 -5697
rect 7486 -5749 7498 -5697
rect 7550 -5749 7566 -5697
rect 7618 -5749 7630 -5697
rect 7682 -5749 7694 -5697
rect 7746 -5749 8094 -5697
rect 8146 -5749 8158 -5697
rect 8210 -5749 8222 -5697
rect 8274 -5749 8290 -5697
rect 8342 -5749 8354 -5697
rect 8406 -5749 8418 -5697
rect 8470 -5749 8580 -5697
rect 8632 -5749 8644 -5697
rect 8696 -5749 8708 -5697
rect 8760 -5749 8776 -5697
rect 8828 -5749 8840 -5697
rect 8892 -5749 8904 -5697
rect 8956 -5749 9006 -5697
rect 1489 -5768 9006 -5749
rect 1489 -5836 9006 -5818
rect 1489 -5888 1539 -5836
rect 1591 -5888 1603 -5836
rect 1655 -5888 1667 -5836
rect 1719 -5888 1735 -5836
rect 1787 -5888 1799 -5836
rect 1851 -5888 1863 -5836
rect 1915 -5888 2025 -5836
rect 2077 -5888 2089 -5836
rect 2141 -5888 2153 -5836
rect 2205 -5888 2221 -5836
rect 2273 -5888 2285 -5836
rect 2337 -5888 2349 -5836
rect 2401 -5840 3737 -5836
rect 2401 -5888 3449 -5840
rect 1489 -5896 3449 -5888
rect 3505 -5896 3529 -5840
rect 3585 -5896 3609 -5840
rect 3665 -5888 3737 -5840
rect 3789 -5888 3801 -5836
rect 3853 -5888 3865 -5836
rect 3917 -5888 3933 -5836
rect 3985 -5888 3997 -5836
rect 4049 -5888 4061 -5836
rect 4113 -5888 4223 -5836
rect 4275 -5888 4287 -5836
rect 4339 -5888 4351 -5836
rect 4403 -5888 4419 -5836
rect 4471 -5888 4483 -5836
rect 4535 -5888 4547 -5836
rect 4599 -5888 5896 -5836
rect 5948 -5888 5960 -5836
rect 6012 -5888 6024 -5836
rect 6076 -5888 6092 -5836
rect 6144 -5888 6156 -5836
rect 6208 -5888 6220 -5836
rect 6272 -5888 6382 -5836
rect 6434 -5888 6446 -5836
rect 6498 -5888 6510 -5836
rect 6562 -5888 6578 -5836
rect 6630 -5888 6642 -5836
rect 6694 -5888 6706 -5836
rect 6758 -5840 8094 -5836
rect 6758 -5888 6830 -5840
rect 3665 -5896 6830 -5888
rect 6886 -5896 6910 -5840
rect 6966 -5896 6990 -5840
rect 7046 -5888 8094 -5840
rect 8146 -5888 8158 -5836
rect 8210 -5888 8222 -5836
rect 8274 -5888 8290 -5836
rect 8342 -5888 8354 -5836
rect 8406 -5888 8418 -5836
rect 8470 -5888 8580 -5836
rect 8632 -5888 8644 -5836
rect 8696 -5888 8708 -5836
rect 8760 -5888 8776 -5836
rect 8828 -5888 8840 -5836
rect 8892 -5888 8904 -5836
rect 8956 -5888 9006 -5836
rect 7046 -5896 9006 -5888
rect 1489 -5906 9006 -5896
rect 3409 -5918 3709 -5906
rect 6786 -5918 7086 -5906
rect 881 -6271 9614 -6261
rect 881 -6283 2591 -6271
rect 881 -6339 932 -6283
rect 988 -6339 1012 -6283
rect 1068 -6339 1092 -6283
rect 1148 -6323 2591 -6283
rect 2643 -6323 2655 -6271
rect 2707 -6323 2719 -6271
rect 2771 -6323 3108 -6271
rect 3160 -6323 3172 -6271
rect 3224 -6323 3236 -6271
rect 3288 -6323 7207 -6271
rect 7259 -6323 7271 -6271
rect 7323 -6323 7335 -6271
rect 7387 -6323 7724 -6271
rect 7776 -6323 7788 -6271
rect 7840 -6323 7852 -6271
rect 7904 -6283 9614 -6271
rect 7904 -6323 9347 -6283
rect 1148 -6339 9347 -6323
rect 9403 -6339 9427 -6283
rect 9483 -6339 9507 -6283
rect 9563 -6339 9614 -6283
rect 881 -6361 9614 -6339
rect 1618 -6416 8878 -6406
rect 1618 -6468 1625 -6416
rect 1677 -6468 1689 -6416
rect 1741 -6468 1753 -6416
rect 1805 -6468 2142 -6416
rect 2194 -6468 2206 -6416
rect 2258 -6468 2270 -6416
rect 2322 -6468 3819 -6416
rect 3871 -6468 3883 -6416
rect 3935 -6468 3947 -6416
rect 3999 -6468 4336 -6416
rect 4388 -6468 4400 -6416
rect 4452 -6468 4464 -6416
rect 4516 -6428 5979 -6416
rect 4516 -6468 4566 -6428
rect 1618 -6484 4566 -6468
rect 4622 -6484 4646 -6428
rect 4702 -6484 4726 -6428
rect 4782 -6484 5713 -6428
rect 5769 -6484 5793 -6428
rect 5849 -6484 5873 -6428
rect 5929 -6468 5979 -6428
rect 6031 -6468 6043 -6416
rect 6095 -6468 6107 -6416
rect 6159 -6468 6496 -6416
rect 6548 -6468 6560 -6416
rect 6612 -6468 6624 -6416
rect 6676 -6468 8173 -6416
rect 8225 -6468 8237 -6416
rect 8289 -6468 8301 -6416
rect 8353 -6468 8691 -6416
rect 8743 -6468 8755 -6416
rect 8807 -6468 8819 -6416
rect 8871 -6468 8878 -6416
rect 5929 -6484 8878 -6468
rect 1618 -6506 8878 -6484
rect 1315 -6577 9181 -6567
rect 1315 -6589 2849 -6577
rect 1315 -6645 1355 -6589
rect 1411 -6645 1435 -6589
rect 1491 -6645 1515 -6589
rect 1571 -6629 2849 -6589
rect 2901 -6629 2913 -6577
rect 2965 -6629 2977 -6577
rect 3029 -6629 3366 -6577
rect 3418 -6629 3430 -6577
rect 3482 -6629 3494 -6577
rect 3546 -6629 6949 -6577
rect 7001 -6629 7013 -6577
rect 7065 -6629 7077 -6577
rect 7129 -6629 7466 -6577
rect 7518 -6629 7530 -6577
rect 7582 -6629 7594 -6577
rect 7646 -6589 9181 -6577
rect 7646 -6629 8925 -6589
rect 1571 -6645 8925 -6629
rect 8981 -6645 9005 -6589
rect 9061 -6645 9085 -6589
rect 9141 -6645 9181 -6589
rect 1315 -6667 9181 -6645
rect 1360 -6717 9136 -6707
rect 1360 -6769 1367 -6717
rect 1419 -6769 1431 -6717
rect 1483 -6769 1495 -6717
rect 1547 -6769 1882 -6717
rect 1934 -6769 1946 -6717
rect 1998 -6769 2010 -6717
rect 2062 -6769 2399 -6717
rect 2451 -6769 2463 -6717
rect 2515 -6769 2527 -6717
rect 2579 -6769 3559 -6717
rect 3611 -6769 3623 -6717
rect 3675 -6769 3687 -6717
rect 3739 -6769 4076 -6717
rect 4128 -6769 4140 -6717
rect 4192 -6769 4204 -6717
rect 4256 -6769 4593 -6717
rect 4645 -6769 4657 -6717
rect 4709 -6769 4721 -6717
rect 4773 -6729 5722 -6717
rect 4773 -6769 5001 -6729
rect 1360 -6785 5001 -6769
rect 5057 -6785 5081 -6729
rect 5137 -6785 5161 -6729
rect 5217 -6785 5278 -6729
rect 5334 -6785 5358 -6729
rect 5414 -6785 5438 -6729
rect 5494 -6769 5722 -6729
rect 5774 -6769 5786 -6717
rect 5838 -6769 5850 -6717
rect 5902 -6769 6239 -6717
rect 6291 -6769 6303 -6717
rect 6355 -6769 6367 -6717
rect 6419 -6769 6756 -6717
rect 6808 -6769 6820 -6717
rect 6872 -6769 6884 -6717
rect 6936 -6769 7916 -6717
rect 7968 -6769 7980 -6717
rect 8032 -6769 8044 -6717
rect 8096 -6769 8434 -6717
rect 8486 -6769 8498 -6717
rect 8550 -6769 8562 -6717
rect 8614 -6769 8949 -6717
rect 9001 -6769 9013 -6717
rect 9065 -6769 9077 -6717
rect 9129 -6769 9136 -6717
rect 5494 -6785 9136 -6769
rect 1360 -6807 9136 -6785
rect 1489 -7166 9006 -7145
rect 1489 -7218 1539 -7166
rect 1591 -7218 1603 -7166
rect 1655 -7218 1667 -7166
rect 1719 -7218 1735 -7166
rect 1787 -7218 1799 -7166
rect 1851 -7218 1863 -7166
rect 1915 -7218 2025 -7166
rect 2077 -7218 2089 -7166
rect 2141 -7218 2153 -7166
rect 2205 -7218 2221 -7166
rect 2273 -7218 2285 -7166
rect 2337 -7218 2349 -7166
rect 2401 -7167 3737 -7166
rect 2401 -7218 3449 -7167
rect 1489 -7223 3449 -7218
rect 3505 -7223 3529 -7167
rect 3585 -7223 3609 -7167
rect 3665 -7218 3737 -7167
rect 3789 -7218 3801 -7166
rect 3853 -7218 3865 -7166
rect 3917 -7218 3933 -7166
rect 3985 -7218 3997 -7166
rect 4049 -7218 4061 -7166
rect 4113 -7218 4223 -7166
rect 4275 -7218 4287 -7166
rect 4339 -7218 4351 -7166
rect 4403 -7218 4419 -7166
rect 4471 -7218 4483 -7166
rect 4535 -7218 4547 -7166
rect 4599 -7218 5896 -7166
rect 5948 -7218 5960 -7166
rect 6012 -7218 6024 -7166
rect 6076 -7218 6092 -7166
rect 6144 -7218 6156 -7166
rect 6208 -7218 6220 -7166
rect 6272 -7218 6382 -7166
rect 6434 -7218 6446 -7166
rect 6498 -7218 6510 -7166
rect 6562 -7218 6578 -7166
rect 6630 -7218 6642 -7166
rect 6694 -7218 6706 -7166
rect 6758 -7167 8094 -7166
rect 6758 -7218 6830 -7167
rect 3665 -7223 6830 -7218
rect 6886 -7223 6910 -7167
rect 6966 -7223 6990 -7167
rect 7046 -7218 8094 -7167
rect 8146 -7218 8158 -7166
rect 8210 -7218 8222 -7166
rect 8274 -7218 8290 -7166
rect 8342 -7218 8354 -7166
rect 8406 -7218 8418 -7166
rect 8470 -7218 8580 -7166
rect 8632 -7218 8644 -7166
rect 8696 -7218 8708 -7166
rect 8760 -7218 8776 -7166
rect 8828 -7218 8840 -7166
rect 8892 -7218 8904 -7166
rect 8956 -7218 9006 -7166
rect 7046 -7223 9006 -7218
rect 1489 -7233 9006 -7223
rect 3409 -7245 3709 -7233
rect 6786 -7245 7086 -7233
rect 1489 -7344 9006 -7327
rect 1489 -7396 1539 -7344
rect 1591 -7396 1603 -7344
rect 1655 -7396 1667 -7344
rect 1719 -7396 1735 -7344
rect 1787 -7396 1799 -7344
rect 1851 -7396 1863 -7344
rect 1915 -7396 2025 -7344
rect 2077 -7396 2089 -7344
rect 2141 -7396 2153 -7344
rect 2205 -7396 2221 -7344
rect 2273 -7396 2285 -7344
rect 2337 -7396 2349 -7344
rect 2401 -7396 2749 -7344
rect 2801 -7396 2813 -7344
rect 2865 -7396 2877 -7344
rect 2929 -7396 2945 -7344
rect 2997 -7396 3009 -7344
rect 3061 -7396 3073 -7344
rect 3125 -7396 3137 -7344
rect 3189 -7396 3205 -7344
rect 3257 -7396 3269 -7344
rect 3321 -7396 3333 -7344
rect 3385 -7396 3737 -7344
rect 3789 -7396 3801 -7344
rect 3853 -7396 3865 -7344
rect 3917 -7396 3933 -7344
rect 3985 -7396 3997 -7344
rect 4049 -7396 4061 -7344
rect 4113 -7396 4223 -7344
rect 4275 -7396 4287 -7344
rect 4339 -7396 4351 -7344
rect 4403 -7396 4419 -7344
rect 4471 -7396 4483 -7344
rect 4535 -7396 4547 -7344
rect 4599 -7396 5896 -7344
rect 5948 -7396 5960 -7344
rect 6012 -7396 6024 -7344
rect 6076 -7396 6092 -7344
rect 6144 -7396 6156 -7344
rect 6208 -7396 6220 -7344
rect 6272 -7396 6382 -7344
rect 6434 -7396 6446 -7344
rect 6498 -7396 6510 -7344
rect 6562 -7396 6578 -7344
rect 6630 -7396 6642 -7344
rect 6694 -7396 6706 -7344
rect 6758 -7396 7110 -7344
rect 7162 -7396 7174 -7344
rect 7226 -7396 7238 -7344
rect 7290 -7396 7306 -7344
rect 7358 -7396 7370 -7344
rect 7422 -7396 7434 -7344
rect 7486 -7396 7498 -7344
rect 7550 -7396 7566 -7344
rect 7618 -7396 7630 -7344
rect 7682 -7396 7694 -7344
rect 7746 -7396 8094 -7344
rect 8146 -7396 8158 -7344
rect 8210 -7396 8222 -7344
rect 8274 -7396 8290 -7344
rect 8342 -7396 8354 -7344
rect 8406 -7396 8418 -7344
rect 8470 -7396 8580 -7344
rect 8632 -7396 8644 -7344
rect 8696 -7396 8708 -7344
rect 8760 -7396 8776 -7344
rect 8828 -7396 8840 -7344
rect 8892 -7396 8904 -7344
rect 8956 -7396 9006 -7344
rect 1489 -7415 9006 -7396
rect 1489 -7483 9006 -7465
rect 1489 -7535 1539 -7483
rect 1591 -7535 1603 -7483
rect 1655 -7535 1667 -7483
rect 1719 -7535 1735 -7483
rect 1787 -7535 1799 -7483
rect 1851 -7535 1863 -7483
rect 1915 -7535 2025 -7483
rect 2077 -7535 2089 -7483
rect 2141 -7535 2153 -7483
rect 2205 -7535 2221 -7483
rect 2273 -7535 2285 -7483
rect 2337 -7535 2349 -7483
rect 2401 -7487 3737 -7483
rect 2401 -7535 2481 -7487
rect 1489 -7543 2481 -7535
rect 2537 -7543 2561 -7487
rect 2617 -7543 2641 -7487
rect 2697 -7535 3737 -7487
rect 3789 -7535 3801 -7483
rect 3853 -7535 3865 -7483
rect 3917 -7535 3933 -7483
rect 3985 -7535 3997 -7483
rect 4049 -7535 4061 -7483
rect 4113 -7535 4223 -7483
rect 4275 -7535 4287 -7483
rect 4339 -7535 4351 -7483
rect 4403 -7535 4419 -7483
rect 4471 -7535 4483 -7483
rect 4535 -7535 4547 -7483
rect 4599 -7535 5896 -7483
rect 5948 -7535 5960 -7483
rect 6012 -7535 6024 -7483
rect 6076 -7535 6092 -7483
rect 6144 -7535 6156 -7483
rect 6208 -7535 6220 -7483
rect 6272 -7535 6382 -7483
rect 6434 -7535 6446 -7483
rect 6498 -7535 6510 -7483
rect 6562 -7535 6578 -7483
rect 6630 -7535 6642 -7483
rect 6694 -7535 6706 -7483
rect 6758 -7487 8094 -7483
rect 6758 -7535 7798 -7487
rect 2697 -7543 7798 -7535
rect 7854 -7543 7878 -7487
rect 7934 -7543 7958 -7487
rect 8014 -7535 8094 -7487
rect 8146 -7535 8158 -7483
rect 8210 -7535 8222 -7483
rect 8274 -7535 8290 -7483
rect 8342 -7535 8354 -7483
rect 8406 -7535 8418 -7483
rect 8470 -7535 8580 -7483
rect 8632 -7535 8644 -7483
rect 8696 -7535 8708 -7483
rect 8760 -7535 8776 -7483
rect 8828 -7535 8840 -7483
rect 8892 -7535 8904 -7483
rect 8956 -7535 9006 -7483
rect 8014 -7543 9006 -7535
rect 1489 -7553 9006 -7543
rect 2441 -7565 2741 -7553
rect 7754 -7565 8054 -7553
rect 1315 -7906 9181 -7896
rect 1315 -7918 1624 -7906
rect 1315 -7974 1355 -7918
rect 1411 -7974 1435 -7918
rect 1491 -7974 1515 -7918
rect 1571 -7958 1624 -7918
rect 1676 -7958 1688 -7906
rect 1740 -7958 1752 -7906
rect 1804 -7958 2141 -7906
rect 2193 -7958 2205 -7906
rect 2257 -7958 2269 -7906
rect 2321 -7958 3818 -7906
rect 3870 -7958 3882 -7906
rect 3934 -7958 3946 -7906
rect 3998 -7958 4335 -7906
rect 4387 -7958 4399 -7906
rect 4451 -7958 4463 -7906
rect 4515 -7958 5980 -7906
rect 6032 -7958 6044 -7906
rect 6096 -7958 6108 -7906
rect 6160 -7958 6497 -7906
rect 6549 -7958 6561 -7906
rect 6613 -7958 6625 -7906
rect 6677 -7958 8174 -7906
rect 8226 -7958 8238 -7906
rect 8290 -7958 8302 -7906
rect 8354 -7958 8692 -7906
rect 8744 -7958 8756 -7906
rect 8808 -7958 8820 -7906
rect 8872 -7918 9181 -7906
rect 8872 -7958 8925 -7918
rect 1571 -7974 8925 -7958
rect 8981 -7974 9005 -7918
rect 9061 -7974 9085 -7918
rect 9141 -7974 9181 -7918
rect 1315 -7996 9181 -7974
rect 2586 -8075 7909 -8065
rect 2586 -8127 2593 -8075
rect 2645 -8127 2657 -8075
rect 2709 -8127 2721 -8075
rect 2773 -8127 3110 -8075
rect 3162 -8127 3174 -8075
rect 3226 -8127 3238 -8075
rect 3290 -8087 7205 -8075
rect 3290 -8127 4566 -8087
rect 2586 -8143 4566 -8127
rect 4622 -8143 4646 -8087
rect 4702 -8143 4726 -8087
rect 4782 -8143 5713 -8087
rect 5769 -8143 5793 -8087
rect 5849 -8143 5873 -8087
rect 5929 -8127 7205 -8087
rect 7257 -8127 7269 -8075
rect 7321 -8127 7333 -8075
rect 7385 -8127 7722 -8075
rect 7774 -8127 7786 -8075
rect 7838 -8127 7850 -8075
rect 7902 -8127 7909 -8075
rect 5929 -8143 7909 -8127
rect 2586 -8165 7909 -8143
rect 892 -8238 9603 -8228
rect 892 -8250 1364 -8238
rect 892 -8306 932 -8250
rect 988 -8306 1012 -8250
rect 1068 -8306 1092 -8250
rect 1148 -8290 1364 -8250
rect 1416 -8290 1428 -8238
rect 1480 -8290 1492 -8238
rect 1544 -8290 1882 -8238
rect 1934 -8290 1946 -8238
rect 1998 -8290 2010 -8238
rect 2062 -8290 2398 -8238
rect 2450 -8290 2462 -8238
rect 2514 -8290 2526 -8238
rect 2578 -8290 3559 -8238
rect 3611 -8290 3623 -8238
rect 3675 -8290 3687 -8238
rect 3739 -8290 4076 -8238
rect 4128 -8290 4140 -8238
rect 4192 -8290 4204 -8238
rect 4256 -8290 4591 -8238
rect 4643 -8290 4655 -8238
rect 4707 -8290 4719 -8238
rect 4771 -8290 5724 -8238
rect 5776 -8290 5788 -8238
rect 5840 -8290 5852 -8238
rect 5904 -8290 6239 -8238
rect 6291 -8290 6303 -8238
rect 6355 -8290 6367 -8238
rect 6419 -8290 6756 -8238
rect 6808 -8290 6820 -8238
rect 6872 -8290 6884 -8238
rect 6936 -8290 7917 -8238
rect 7969 -8290 7981 -8238
rect 8033 -8290 8045 -8238
rect 8097 -8290 8434 -8238
rect 8486 -8290 8498 -8238
rect 8550 -8290 8562 -8238
rect 8614 -8290 8951 -8238
rect 9003 -8290 9015 -8238
rect 9067 -8290 9079 -8238
rect 9131 -8250 9603 -8238
rect 9131 -8290 9347 -8250
rect 1148 -8306 9347 -8290
rect 9403 -8306 9427 -8250
rect 9483 -8306 9507 -8250
rect 9563 -8306 9603 -8250
rect 892 -8328 9603 -8306
rect 2843 -8406 7652 -8396
rect 2843 -8458 2850 -8406
rect 2902 -8458 2914 -8406
rect 2966 -8458 2978 -8406
rect 3030 -8458 3368 -8406
rect 3420 -8458 3432 -8406
rect 3484 -8458 3496 -8406
rect 3548 -8418 6948 -8406
rect 3548 -8458 5001 -8418
rect 2843 -8474 5001 -8458
rect 5057 -8474 5081 -8418
rect 5137 -8474 5161 -8418
rect 5217 -8474 5278 -8418
rect 5334 -8474 5358 -8418
rect 5414 -8474 5438 -8418
rect 5494 -8458 6948 -8418
rect 7000 -8458 7012 -8406
rect 7064 -8458 7076 -8406
rect 7128 -8458 7465 -8406
rect 7517 -8458 7529 -8406
rect 7581 -8458 7593 -8406
rect 7645 -8458 7652 -8406
rect 5494 -8474 7652 -8458
rect 2843 -8496 7652 -8474
<< via2 >>
rect 5001 241 5057 297
rect 5081 241 5137 297
rect 5161 241 5217 297
rect 5278 241 5334 297
rect 5358 241 5414 297
rect 5438 241 5494 297
rect 932 72 988 128
rect 1012 72 1068 128
rect 1092 72 1148 128
rect 9347 72 9403 128
rect 9427 72 9483 128
rect 9507 72 9563 128
rect 4566 -91 4622 -35
rect 4646 -91 4702 -35
rect 4726 -91 4782 -35
rect 5713 -91 5769 -35
rect 5793 -91 5849 -35
rect 5873 -91 5929 -35
rect 1355 -259 1411 -203
rect 1435 -259 1491 -203
rect 1515 -259 1571 -203
rect 8925 -259 8981 -203
rect 9005 -259 9061 -203
rect 9085 -259 9141 -203
rect 2481 -691 2537 -635
rect 2561 -691 2617 -635
rect 2641 -691 2697 -635
rect 7798 -691 7854 -635
rect 7878 -691 7934 -635
rect 7958 -691 8014 -635
rect 3449 -1011 3505 -955
rect 3529 -1011 3585 -955
rect 3609 -1011 3665 -955
rect 6830 -1011 6886 -955
rect 6910 -1011 6966 -955
rect 6990 -1011 7046 -955
rect 5001 -1449 5057 -1393
rect 5081 -1449 5137 -1393
rect 5161 -1449 5217 -1393
rect 5278 -1449 5334 -1393
rect 5358 -1449 5414 -1393
rect 5438 -1449 5494 -1393
rect 1355 -1589 1411 -1533
rect 1435 -1589 1491 -1533
rect 1515 -1589 1571 -1533
rect 8925 -1589 8981 -1533
rect 9005 -1589 9061 -1533
rect 9085 -1589 9141 -1533
rect 4566 -1750 4622 -1694
rect 4646 -1750 4702 -1694
rect 4726 -1750 4782 -1694
rect 5713 -1750 5769 -1694
rect 5793 -1750 5849 -1694
rect 5873 -1750 5929 -1694
rect 932 -1894 988 -1838
rect 1012 -1894 1068 -1838
rect 1092 -1894 1148 -1838
rect 9347 -1894 9403 -1838
rect 9427 -1894 9483 -1838
rect 9507 -1894 9563 -1838
rect 3449 -2338 3505 -2282
rect 3529 -2338 3585 -2282
rect 3609 -2338 3665 -2282
rect 6830 -2349 6886 -2293
rect 6910 -2349 6966 -2293
rect 6990 -2349 7046 -2293
rect 2481 -2670 2537 -2614
rect 2561 -2670 2617 -2614
rect 2641 -2670 2697 -2614
rect 7798 -2670 7854 -2614
rect 7878 -2670 7934 -2614
rect 7958 -2670 8014 -2614
rect 1355 -3101 1411 -3045
rect 1435 -3101 1491 -3045
rect 1515 -3101 1571 -3045
rect 8925 -3101 8981 -3045
rect 9005 -3101 9061 -3045
rect 9085 -3101 9141 -3045
rect 4566 -3270 4622 -3214
rect 4646 -3270 4702 -3214
rect 4726 -3270 4782 -3214
rect 5713 -3270 5769 -3214
rect 5793 -3270 5849 -3214
rect 5873 -3270 5929 -3214
rect 932 -3432 988 -3376
rect 1012 -3432 1068 -3376
rect 1092 -3432 1148 -3376
rect 9347 -3432 9403 -3376
rect 9427 -3432 9483 -3376
rect 9507 -3432 9563 -3376
rect 5001 -3601 5057 -3545
rect 5081 -3601 5137 -3545
rect 5161 -3601 5217 -3545
rect 5278 -3601 5334 -3545
rect 5358 -3601 5414 -3545
rect 5438 -3601 5494 -3545
rect 5001 -4632 5057 -4576
rect 5081 -4632 5137 -4576
rect 5161 -4632 5217 -4576
rect 5278 -4632 5334 -4576
rect 5358 -4632 5414 -4576
rect 5438 -4632 5494 -4576
rect 932 -4801 988 -4745
rect 1012 -4801 1068 -4745
rect 1092 -4801 1148 -4745
rect 9347 -4801 9403 -4745
rect 9427 -4801 9483 -4745
rect 9507 -4801 9563 -4745
rect 4566 -4964 4622 -4908
rect 4646 -4964 4702 -4908
rect 4726 -4964 4782 -4908
rect 5713 -4964 5769 -4908
rect 5793 -4964 5849 -4908
rect 5873 -4964 5929 -4908
rect 1355 -5133 1411 -5077
rect 1435 -5133 1491 -5077
rect 1515 -5133 1571 -5077
rect 8925 -5133 8981 -5077
rect 9005 -5133 9061 -5077
rect 9085 -5133 9141 -5077
rect 2481 -5564 2537 -5508
rect 2561 -5564 2617 -5508
rect 2641 -5564 2697 -5508
rect 7798 -5564 7854 -5508
rect 7878 -5564 7934 -5508
rect 7958 -5564 8014 -5508
rect 3449 -5896 3505 -5840
rect 3529 -5896 3585 -5840
rect 3609 -5896 3665 -5840
rect 6830 -5896 6886 -5840
rect 6910 -5896 6966 -5840
rect 6990 -5896 7046 -5840
rect 932 -6339 988 -6283
rect 1012 -6339 1068 -6283
rect 1092 -6339 1148 -6283
rect 9347 -6339 9403 -6283
rect 9427 -6339 9483 -6283
rect 9507 -6339 9563 -6283
rect 4566 -6484 4622 -6428
rect 4646 -6484 4702 -6428
rect 4726 -6484 4782 -6428
rect 5713 -6484 5769 -6428
rect 5793 -6484 5849 -6428
rect 5873 -6484 5929 -6428
rect 1355 -6645 1411 -6589
rect 1435 -6645 1491 -6589
rect 1515 -6645 1571 -6589
rect 8925 -6645 8981 -6589
rect 9005 -6645 9061 -6589
rect 9085 -6645 9141 -6589
rect 5001 -6785 5057 -6729
rect 5081 -6785 5137 -6729
rect 5161 -6785 5217 -6729
rect 5278 -6785 5334 -6729
rect 5358 -6785 5414 -6729
rect 5438 -6785 5494 -6729
rect 3449 -7223 3505 -7167
rect 3529 -7223 3585 -7167
rect 3609 -7223 3665 -7167
rect 6830 -7223 6886 -7167
rect 6910 -7223 6966 -7167
rect 6990 -7223 7046 -7167
rect 2481 -7543 2537 -7487
rect 2561 -7543 2617 -7487
rect 2641 -7543 2697 -7487
rect 7798 -7543 7854 -7487
rect 7878 -7543 7934 -7487
rect 7958 -7543 8014 -7487
rect 1355 -7974 1411 -7918
rect 1435 -7974 1491 -7918
rect 1515 -7974 1571 -7918
rect 8925 -7974 8981 -7918
rect 9005 -7974 9061 -7918
rect 9085 -7974 9141 -7918
rect 4566 -8143 4622 -8087
rect 4646 -8143 4702 -8087
rect 4726 -8143 4782 -8087
rect 5713 -8143 5769 -8087
rect 5793 -8143 5849 -8087
rect 5873 -8143 5929 -8087
rect 932 -8306 988 -8250
rect 1012 -8306 1068 -8250
rect 1092 -8306 1148 -8250
rect 9347 -8306 9403 -8250
rect 9427 -8306 9483 -8250
rect 9507 -8306 9563 -8250
rect 5001 -8474 5057 -8418
rect 5081 -8474 5137 -8418
rect 5161 -8474 5217 -8418
rect 5278 -8474 5334 -8418
rect 5358 -8474 5414 -8418
rect 5438 -8474 5494 -8418
<< metal3 >>
rect 4957 297 5538 319
rect 4957 241 5001 297
rect 5057 241 5081 297
rect 5137 241 5161 297
rect 5217 241 5278 297
rect 5334 241 5358 297
rect 5414 241 5438 297
rect 5494 241 5538 297
rect 892 128 1192 150
rect 892 72 932 128
rect 988 72 1012 128
rect 1068 72 1092 128
rect 1148 72 1192 128
rect 892 -1838 1192 72
rect 4522 -35 4822 -13
rect 4522 -91 4566 -35
rect 4622 -91 4646 -35
rect 4702 -91 4726 -35
rect 4782 -91 4822 -35
rect 892 -1894 932 -1838
rect 988 -1894 1012 -1838
rect 1068 -1894 1092 -1838
rect 1148 -1894 1192 -1838
rect 892 -3376 1192 -1894
rect 892 -3432 932 -3376
rect 988 -3432 1012 -3376
rect 1068 -3432 1092 -3376
rect 1148 -3432 1192 -3376
rect 892 -4745 1192 -3432
rect 892 -4801 932 -4745
rect 988 -4801 1012 -4745
rect 1068 -4801 1092 -4745
rect 1148 -4801 1192 -4745
rect 892 -6283 1192 -4801
rect 892 -6339 932 -6283
rect 988 -6339 1012 -6283
rect 1068 -6339 1092 -6283
rect 1148 -6339 1192 -6283
rect 892 -8250 1192 -6339
rect 1315 -203 1615 -181
rect 1315 -259 1355 -203
rect 1411 -259 1435 -203
rect 1491 -259 1515 -203
rect 1571 -259 1615 -203
rect 1315 -1533 1615 -259
rect 1315 -1589 1355 -1533
rect 1411 -1589 1435 -1533
rect 1491 -1589 1515 -1533
rect 1571 -1589 1615 -1533
rect 1315 -3045 1615 -1589
rect 1315 -3101 1355 -3045
rect 1411 -3101 1435 -3045
rect 1491 -3101 1515 -3045
rect 1571 -3101 1615 -3045
rect 1315 -5077 1615 -3101
rect 1315 -5133 1355 -5077
rect 1411 -5133 1435 -5077
rect 1491 -5133 1515 -5077
rect 1571 -5133 1615 -5077
rect 1315 -6589 1615 -5133
rect 1315 -6645 1355 -6589
rect 1411 -6645 1435 -6589
rect 1491 -6645 1515 -6589
rect 1571 -6645 1615 -6589
rect 1315 -7918 1615 -6645
rect 2441 -635 2741 -613
rect 2441 -691 2481 -635
rect 2537 -691 2561 -635
rect 2617 -691 2641 -635
rect 2697 -691 2741 -635
rect 2441 -2614 2741 -691
rect 2441 -2670 2481 -2614
rect 2537 -2670 2561 -2614
rect 2617 -2670 2641 -2614
rect 2697 -2670 2741 -2614
rect 2441 -5508 2741 -2670
rect 2441 -5564 2481 -5508
rect 2537 -5564 2561 -5508
rect 2617 -5564 2641 -5508
rect 2697 -5564 2741 -5508
rect 2441 -7487 2741 -5564
rect 3409 -955 3709 -933
rect 3409 -1011 3449 -955
rect 3505 -1011 3529 -955
rect 3585 -1011 3609 -955
rect 3665 -1011 3709 -955
rect 3409 -2282 3709 -1011
rect 3409 -2338 3449 -2282
rect 3505 -2338 3529 -2282
rect 3585 -2338 3609 -2282
rect 3665 -2338 3709 -2282
rect 3409 -5840 3709 -2338
rect 3409 -5896 3449 -5840
rect 3505 -5896 3529 -5840
rect 3585 -5896 3609 -5840
rect 3665 -5896 3709 -5840
rect 3409 -7167 3709 -5896
rect 3409 -7223 3449 -7167
rect 3505 -7223 3529 -7167
rect 3585 -7223 3609 -7167
rect 3665 -7223 3709 -7167
rect 3409 -7245 3709 -7223
rect 4522 -1694 4822 -91
rect 4522 -1750 4566 -1694
rect 4622 -1750 4646 -1694
rect 4702 -1750 4726 -1694
rect 4782 -1750 4822 -1694
rect 4522 -3214 4822 -1750
rect 4522 -3270 4566 -3214
rect 4622 -3270 4646 -3214
rect 4702 -3270 4726 -3214
rect 4782 -3270 4822 -3214
rect 4522 -4908 4822 -3270
rect 4522 -4964 4566 -4908
rect 4622 -4964 4646 -4908
rect 4702 -4964 4726 -4908
rect 4782 -4964 4822 -4908
rect 4522 -6428 4822 -4964
rect 4522 -6484 4566 -6428
rect 4622 -6484 4646 -6428
rect 4702 -6484 4726 -6428
rect 4782 -6484 4822 -6428
rect 2441 -7543 2481 -7487
rect 2537 -7543 2561 -7487
rect 2617 -7543 2641 -7487
rect 2697 -7543 2741 -7487
rect 2441 -7565 2741 -7543
rect 1315 -7974 1355 -7918
rect 1411 -7974 1435 -7918
rect 1491 -7974 1515 -7918
rect 1571 -7974 1615 -7918
rect 1315 -7996 1615 -7974
rect 4522 -8087 4822 -6484
rect 4522 -8143 4566 -8087
rect 4622 -8143 4646 -8087
rect 4702 -8143 4726 -8087
rect 4782 -8143 4822 -8087
rect 4522 -8165 4822 -8143
rect 4957 -1393 5538 241
rect 9303 128 9603 150
rect 9303 72 9347 128
rect 9403 72 9427 128
rect 9483 72 9507 128
rect 9563 72 9603 128
rect 4957 -1449 5001 -1393
rect 5057 -1449 5081 -1393
rect 5137 -1449 5161 -1393
rect 5217 -1449 5278 -1393
rect 5334 -1449 5358 -1393
rect 5414 -1449 5438 -1393
rect 5494 -1449 5538 -1393
rect 4957 -3545 5538 -1449
rect 4957 -3601 5001 -3545
rect 5057 -3601 5081 -3545
rect 5137 -3601 5161 -3545
rect 5217 -3601 5278 -3545
rect 5334 -3601 5358 -3545
rect 5414 -3601 5438 -3545
rect 5494 -3601 5538 -3545
rect 4957 -4576 5538 -3601
rect 4957 -4632 5001 -4576
rect 5057 -4632 5081 -4576
rect 5137 -4632 5161 -4576
rect 5217 -4632 5278 -4576
rect 5334 -4632 5358 -4576
rect 5414 -4632 5438 -4576
rect 5494 -4632 5538 -4576
rect 4957 -6729 5538 -4632
rect 4957 -6785 5001 -6729
rect 5057 -6785 5081 -6729
rect 5137 -6785 5161 -6729
rect 5217 -6785 5278 -6729
rect 5334 -6785 5358 -6729
rect 5414 -6785 5438 -6729
rect 5494 -6785 5538 -6729
rect 892 -8306 932 -8250
rect 988 -8306 1012 -8250
rect 1068 -8306 1092 -8250
rect 1148 -8306 1192 -8250
rect 892 -8328 1192 -8306
rect 4957 -8418 5538 -6785
rect 5673 -35 5973 -13
rect 5673 -91 5713 -35
rect 5769 -91 5793 -35
rect 5849 -91 5873 -35
rect 5929 -91 5973 -35
rect 5673 -1694 5973 -91
rect 8881 -203 9181 -181
rect 8881 -259 8925 -203
rect 8981 -259 9005 -203
rect 9061 -259 9085 -203
rect 9141 -259 9181 -203
rect 7754 -635 8054 -613
rect 7754 -691 7798 -635
rect 7854 -691 7878 -635
rect 7934 -691 7958 -635
rect 8014 -691 8054 -635
rect 5673 -1750 5713 -1694
rect 5769 -1750 5793 -1694
rect 5849 -1750 5873 -1694
rect 5929 -1750 5973 -1694
rect 5673 -3214 5973 -1750
rect 5673 -3270 5713 -3214
rect 5769 -3270 5793 -3214
rect 5849 -3270 5873 -3214
rect 5929 -3270 5973 -3214
rect 5673 -4908 5973 -3270
rect 5673 -4964 5713 -4908
rect 5769 -4964 5793 -4908
rect 5849 -4964 5873 -4908
rect 5929 -4964 5973 -4908
rect 5673 -6428 5973 -4964
rect 5673 -6484 5713 -6428
rect 5769 -6484 5793 -6428
rect 5849 -6484 5873 -6428
rect 5929 -6484 5973 -6428
rect 5673 -8087 5973 -6484
rect 6786 -955 7086 -933
rect 6786 -1011 6830 -955
rect 6886 -1011 6910 -955
rect 6966 -1011 6990 -955
rect 7046 -1011 7086 -955
rect 6786 -2293 7086 -1011
rect 6786 -2349 6830 -2293
rect 6886 -2349 6910 -2293
rect 6966 -2349 6990 -2293
rect 7046 -2349 7086 -2293
rect 6786 -5840 7086 -2349
rect 6786 -5896 6830 -5840
rect 6886 -5896 6910 -5840
rect 6966 -5896 6990 -5840
rect 7046 -5896 7086 -5840
rect 6786 -7167 7086 -5896
rect 6786 -7223 6830 -7167
rect 6886 -7223 6910 -7167
rect 6966 -7223 6990 -7167
rect 7046 -7223 7086 -7167
rect 6786 -7245 7086 -7223
rect 7754 -2614 8054 -691
rect 7754 -2670 7798 -2614
rect 7854 -2670 7878 -2614
rect 7934 -2670 7958 -2614
rect 8014 -2670 8054 -2614
rect 7754 -5508 8054 -2670
rect 7754 -5564 7798 -5508
rect 7854 -5564 7878 -5508
rect 7934 -5564 7958 -5508
rect 8014 -5564 8054 -5508
rect 7754 -7487 8054 -5564
rect 7754 -7543 7798 -7487
rect 7854 -7543 7878 -7487
rect 7934 -7543 7958 -7487
rect 8014 -7543 8054 -7487
rect 7754 -7565 8054 -7543
rect 8881 -1533 9181 -259
rect 8881 -1589 8925 -1533
rect 8981 -1589 9005 -1533
rect 9061 -1589 9085 -1533
rect 9141 -1589 9181 -1533
rect 8881 -3045 9181 -1589
rect 8881 -3101 8925 -3045
rect 8981 -3101 9005 -3045
rect 9061 -3101 9085 -3045
rect 9141 -3101 9181 -3045
rect 8881 -5077 9181 -3101
rect 8881 -5133 8925 -5077
rect 8981 -5133 9005 -5077
rect 9061 -5133 9085 -5077
rect 9141 -5133 9181 -5077
rect 8881 -6589 9181 -5133
rect 8881 -6645 8925 -6589
rect 8981 -6645 9005 -6589
rect 9061 -6645 9085 -6589
rect 9141 -6645 9181 -6589
rect 8881 -7918 9181 -6645
rect 8881 -7974 8925 -7918
rect 8981 -7974 9005 -7918
rect 9061 -7974 9085 -7918
rect 9141 -7974 9181 -7918
rect 8881 -7996 9181 -7974
rect 9303 -1838 9603 72
rect 9303 -1894 9347 -1838
rect 9403 -1894 9427 -1838
rect 9483 -1894 9507 -1838
rect 9563 -1894 9603 -1838
rect 9303 -3376 9603 -1894
rect 9303 -3432 9347 -3376
rect 9403 -3432 9427 -3376
rect 9483 -3432 9507 -3376
rect 9563 -3432 9603 -3376
rect 9303 -4745 9603 -3432
rect 9303 -4801 9347 -4745
rect 9403 -4801 9427 -4745
rect 9483 -4801 9507 -4745
rect 9563 -4801 9603 -4745
rect 9303 -6283 9603 -4801
rect 9303 -6339 9347 -6283
rect 9403 -6339 9427 -6283
rect 9483 -6339 9507 -6283
rect 9563 -6339 9603 -6283
rect 5673 -8143 5713 -8087
rect 5769 -8143 5793 -8087
rect 5849 -8143 5873 -8087
rect 5929 -8143 5973 -8087
rect 5673 -8165 5973 -8143
rect 9303 -8250 9603 -6339
rect 9303 -8306 9347 -8250
rect 9403 -8306 9427 -8250
rect 9483 -8306 9507 -8250
rect 9563 -8306 9603 -8250
rect 9303 -8328 9603 -8306
rect 4957 -8474 5001 -8418
rect 5057 -8474 5081 -8418
rect 5137 -8474 5161 -8418
rect 5217 -8474 5278 -8418
rect 5334 -8474 5358 -8418
rect 5414 -8474 5438 -8418
rect 5494 -8474 5538 -8418
rect 4957 -8496 5538 -8474
<< end >>
