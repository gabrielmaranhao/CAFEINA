magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< nwell >>
rect 6036 4621 11696 7504
<< metal1 >>
rect 6076 4628 9953 7484
rect 6953 -3612 8514 -3262
<< metal2 >>
rect 7266 -665 10510 -664
rect 4351 -734 10510 -665
rect 4351 -735 10509 -734
rect 6502 -837 10509 -735
rect 5858 -1097 9591 -1065
rect 5858 -1135 9296 -1097
rect 7196 -1153 9296 -1135
rect 9352 -1153 9376 -1097
rect 9432 -1153 9456 -1097
rect 9512 -1153 9591 -1097
rect 7196 -1197 9591 -1153
rect 7196 -1205 9296 -1197
rect 5858 -1253 9296 -1205
rect 9352 -1253 9376 -1197
rect 9432 -1253 9456 -1197
rect 9512 -1253 9591 -1197
rect 5858 -1275 9591 -1253
rect 12977 -1854 13277 -1832
rect 12977 -1910 13017 -1854
rect 13073 -1910 13097 -1854
rect 13153 -1910 13177 -1854
rect 13233 -1910 13277 -1854
rect 12977 -1954 13277 -1910
rect 12977 -2010 13017 -1954
rect 13073 -2010 13097 -1954
rect 13153 -2010 13177 -1954
rect 13233 -2010 13277 -1954
rect 12977 -2054 13277 -2010
rect 12977 -2110 13017 -2054
rect 13073 -2110 13097 -2054
rect 13153 -2110 13177 -2054
rect 13233 -2110 13277 -2054
rect 12977 -2132 13277 -2110
rect 4775 -3184 7041 -3114
<< via2 >>
rect 9296 -1153 9352 -1097
rect 9376 -1153 9432 -1097
rect 9456 -1153 9512 -1097
rect 9296 -1253 9352 -1197
rect 9376 -1253 9432 -1197
rect 9456 -1253 9512 -1197
rect 13017 -1910 13073 -1854
rect 13097 -1910 13153 -1854
rect 13177 -1910 13233 -1854
rect 13017 -2010 13073 -1954
rect 13097 -2010 13153 -1954
rect 13177 -2010 13233 -1954
rect 13017 -2110 13073 -2054
rect 13097 -2110 13153 -2054
rect 13177 -2110 13233 -2054
<< metal3 >>
rect 1001 4114 1301 6799
rect 2241 4990 2541 7675
rect 8438 598 8738 3494
rect 9256 -1097 9556 1576
rect 10141 -837 10441 2059
rect 11031 1215 11331 6706
rect 9256 -1153 9296 -1097
rect 9352 -1153 9376 -1097
rect 9432 -1153 9456 -1097
rect 9512 -1153 9556 -1097
rect 9256 -1197 9556 -1153
rect 9256 -1253 9296 -1197
rect 9352 -1253 9376 -1197
rect 9432 -1253 9456 -1197
rect 9512 -1253 9556 -1197
rect 9256 -1320 9556 -1253
rect 12977 -1854 13277 -1547
rect 12977 -1910 13017 -1854
rect 13073 -1910 13097 -1854
rect 13153 -1910 13177 -1854
rect 13233 -1910 13277 -1854
rect 12977 -1954 13277 -1910
rect 12977 -2010 13017 -1954
rect 13073 -2010 13097 -1954
rect 13153 -2010 13177 -1954
rect 13233 -2010 13277 -1954
rect 12977 -2054 13277 -2010
rect 12977 -2110 13017 -2054
rect 13073 -2110 13097 -2054
rect 13153 -2110 13177 -2054
rect 13233 -2110 13277 -2054
rect 12977 -2177 13277 -2110
use nbias_vb3  nbias_vb3_0
timestamp 1698888477
transform 1 0 9508 0 1 -1570
box 1048 -754 3305 562
use nbias_vb124  nbias_vb124_0
timestamp 1698888477
transform 1 0 9316 0 1 1285
box -2484 -1841 3567 2164
use pbias_vb4  pbias_vb4_0
timestamp 1698888477
transform 1 0 8850 0 1 6997
box 806 -2412 2846 508
use pbias_vb123  pbias_vb123_0
timestamp 1698888477
transform 1 0 0 0 1 1504
box 290 -5592 6219 6020
<< labels >>
flabel metal3 s 10169 -412 10399 225 2 FreeSans 3126 0 0 0 VB2
port 1 nsew
flabel metal3 s 8468 969 8713 1551 2 FreeSans 3126 0 0 0 IREF
port 2 nsew
flabel metal3 s 12995 -1843 13265 -1567 2 FreeSans 3126 0 0 0 VB3
port 3 nsew
flabel metal3 s 1023 5755 1288 6012 2 FreeSans 3126 0 0 0 AVDD
port 4 nsew
flabel metal3 s 11058 3695 11306 4379 2 FreeSans 3126 0 0 0 VB4
port 5 nsew
flabel metal3 s 2259 7400 2524 7657 2 FreeSans 3126 0 0 0 VB1
port 6 nsew
flabel metal1 s 6953 -3611 8514 -3262 2 FreeSans 3126 0 0 0 AVSS
port 7 nsew
<< end >>
