magic
tech sky130A
timestamp 1697634299
<< nwell >>
rect -745 -599 745 599
<< pwell >>
rect -835 599 835 689
rect -835 -599 -745 599
rect 745 -599 835 599
rect -835 -689 835 -599
<< mvpsubdiff >>
rect -817 665 817 671
rect -817 648 -763 665
rect 763 648 817 665
rect -817 642 817 648
rect -817 617 -788 642
rect -817 -617 -811 617
rect -794 -617 -788 617
rect 788 617 817 642
rect -817 -642 -788 -617
rect 788 -617 794 617
rect 811 -617 817 617
rect 788 -642 817 -617
rect -817 -648 817 -642
rect -817 -665 -763 -648
rect 763 -665 817 -648
rect -817 -671 817 -665
<< mvnsubdiff >>
rect -712 560 -480 566
rect -712 543 -658 560
rect -534 543 -480 560
rect -712 537 -480 543
rect -712 512 -683 537
rect -712 -512 -706 512
rect -689 -512 -683 512
rect -509 512 -480 537
rect -712 -537 -683 -512
rect -509 -512 -503 512
rect -486 -512 -480 512
rect -509 -537 -480 -512
rect -712 -543 -480 -537
rect -712 -560 -658 -543
rect -534 -560 -480 -543
rect -712 -566 -480 -560
rect -414 560 -182 566
rect -414 543 -360 560
rect -236 543 -182 560
rect -414 537 -182 543
rect -414 512 -385 537
rect -414 -512 -408 512
rect -391 -512 -385 512
rect -211 512 -182 537
rect -414 -537 -385 -512
rect -211 -512 -205 512
rect -188 -512 -182 512
rect -211 -537 -182 -512
rect -414 -543 -182 -537
rect -414 -560 -360 -543
rect -236 -560 -182 -543
rect -414 -566 -182 -560
rect -116 560 116 566
rect -116 543 -62 560
rect 62 543 116 560
rect -116 537 116 543
rect -116 512 -87 537
rect -116 -512 -110 512
rect -93 -512 -87 512
rect 87 512 116 537
rect -116 -537 -87 -512
rect 87 -512 93 512
rect 110 -512 116 512
rect 87 -537 116 -512
rect -116 -543 116 -537
rect -116 -560 -62 -543
rect 62 -560 116 -543
rect -116 -566 116 -560
rect 182 560 414 566
rect 182 543 236 560
rect 360 543 414 560
rect 182 537 414 543
rect 182 512 211 537
rect 182 -512 188 512
rect 205 -512 211 512
rect 385 512 414 537
rect 182 -537 211 -512
rect 385 -512 391 512
rect 408 -512 414 512
rect 385 -537 414 -512
rect 182 -543 414 -537
rect 182 -560 236 -543
rect 360 -560 414 -543
rect 182 -566 414 -560
rect 480 560 712 566
rect 480 543 534 560
rect 658 543 712 560
rect 480 537 712 543
rect 480 512 509 537
rect 480 -512 486 512
rect 503 -512 509 512
rect 683 512 712 537
rect 480 -537 509 -512
rect 683 -512 689 512
rect 706 -512 712 512
rect 683 -537 712 -512
rect 480 -543 712 -537
rect 480 -560 534 -543
rect 658 -560 712 -543
rect 480 -566 712 -560
<< mvpsubdiffcont >>
rect -763 648 763 665
rect -811 -617 -794 617
rect 794 -617 811 617
rect -763 -665 763 -648
<< mvnsubdiffcont >>
rect -658 543 -534 560
rect -706 -512 -689 512
rect -503 -512 -486 512
rect -658 -560 -534 -543
rect -360 543 -236 560
rect -408 -512 -391 512
rect -205 -512 -188 512
rect -360 -560 -236 -543
rect -62 543 62 560
rect -110 -512 -93 512
rect 93 -512 110 512
rect -62 -560 62 -543
rect 236 543 360 560
rect 188 -512 205 512
rect 391 -512 408 512
rect 236 -560 360 -543
rect 534 543 658 560
rect 486 -512 503 512
rect 689 -512 706 512
rect 534 -560 658 -543
<< mvpdiode >>
rect -646 494 -546 500
rect -646 -494 -640 494
rect -552 -494 -546 494
rect -646 -500 -546 -494
rect -348 494 -248 500
rect -348 -494 -342 494
rect -254 -494 -248 494
rect -348 -500 -248 -494
rect -50 494 50 500
rect -50 -494 -44 494
rect 44 -494 50 494
rect -50 -500 50 -494
rect 248 494 348 500
rect 248 -494 254 494
rect 342 -494 348 494
rect 248 -500 348 -494
rect 546 494 646 500
rect 546 -494 552 494
rect 640 -494 646 494
rect 546 -500 646 -494
<< mvpdiodec >>
rect -640 -494 -552 494
rect -342 -494 -254 494
rect -44 -494 44 494
rect 254 -494 342 494
rect 552 -494 640 494
<< locali >>
rect -811 648 -763 665
rect 763 648 811 665
rect -811 617 -794 648
rect 794 617 811 648
rect -706 543 -658 560
rect -534 543 -486 560
rect -706 512 -689 543
rect -503 512 -486 543
rect -640 494 -552 502
rect -640 -502 -552 -494
rect -706 -543 -689 -512
rect -503 -543 -486 -512
rect -706 -560 -658 -543
rect -534 -560 -486 -543
rect -408 543 -360 560
rect -236 543 -188 560
rect -408 512 -391 543
rect -205 512 -188 543
rect -342 494 -254 502
rect -342 -502 -254 -494
rect -408 -543 -391 -512
rect -205 -543 -188 -512
rect -408 -560 -360 -543
rect -236 -560 -188 -543
rect -110 543 -62 560
rect 62 543 110 560
rect -110 512 -93 543
rect 93 512 110 543
rect -44 494 44 502
rect -44 -502 44 -494
rect -110 -543 -93 -512
rect 93 -543 110 -512
rect -110 -560 -62 -543
rect 62 -560 110 -543
rect 188 543 236 560
rect 360 543 408 560
rect 188 512 205 543
rect 391 512 408 543
rect 254 494 342 502
rect 254 -502 342 -494
rect 188 -543 205 -512
rect 391 -543 408 -512
rect 188 -560 236 -543
rect 360 -560 408 -543
rect 486 543 534 560
rect 658 543 706 560
rect 486 512 503 543
rect 689 512 706 543
rect 552 494 640 502
rect 552 -502 640 -494
rect 486 -543 503 -512
rect 689 -543 706 -512
rect 486 -560 534 -543
rect 658 -560 706 -543
rect -811 -648 -794 -617
rect 794 -648 811 -617
rect -811 -665 -763 -648
rect 763 -665 811 -648
<< viali >>
rect -640 -494 -552 494
rect -342 -494 -254 494
rect -44 -494 44 494
rect 254 -494 342 494
rect 552 -494 640 494
<< metal1 >>
rect -643 494 -549 500
rect -643 -494 -640 494
rect -552 -494 -549 494
rect -643 -500 -549 -494
rect -345 494 -251 500
rect -345 -494 -342 494
rect -254 -494 -251 494
rect -345 -500 -251 -494
rect -47 494 47 500
rect -47 -494 -44 494
rect 44 -494 47 494
rect -47 -500 47 -494
rect 251 494 345 500
rect 251 -494 254 494
rect 342 -494 345 494
rect 251 -500 345 -494
rect 549 494 643 500
rect 549 -494 552 494
rect 640 -494 643 494
rect 549 -500 643 -494
<< properties >>
string FIXED_BBOX 494 -551 697 551
string gencell sky130_fd_pr__diode_pd2nw_11v0
string library sky130
string parameters w 1 l 10 area 10.0 peri 22.0 nx 5 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
