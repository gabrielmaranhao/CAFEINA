magic
tech sky130A
magscale 1 2
timestamp 1698888477
<< nwell >>
rect 806 -2412 2846 508
<< pmoshvt >>
rect 1017 68 1217 268
rect 1469 68 1669 268
rect 1727 68 1927 268
rect 1985 68 2185 268
rect 2437 68 2637 268
rect 1017 -235 1217 -35
rect 1469 -235 1669 -35
rect 1727 -235 1927 -35
rect 1985 -235 2185 -35
rect 2437 -235 2637 -35
rect 1017 -699 1217 -499
rect 1469 -699 1669 -499
rect 1727 -699 1927 -499
rect 1985 -699 2185 -499
rect 2437 -699 2637 -499
rect 1017 -1002 1217 -802
rect 1469 -1002 1669 -802
rect 1727 -1002 1927 -802
rect 1985 -1002 2185 -802
rect 2437 -1002 2637 -802
rect 1017 -1466 1217 -1266
rect 1469 -1466 1669 -1266
rect 1727 -1466 1927 -1266
rect 1985 -1466 2185 -1266
rect 2437 -1466 2637 -1266
rect 1017 -1769 1217 -1569
rect 1469 -1769 1669 -1569
rect 1727 -1769 1927 -1569
rect 1985 -1769 2185 -1569
rect 2437 -1769 2637 -1569
rect 1017 -2239 1217 -2039
rect 1469 -2239 1669 -2039
rect 1727 -2239 1927 -2039
rect 1985 -2239 2185 -2039
rect 2437 -2239 2637 -2039
<< pdiff >>
rect 959 253 1017 268
rect 959 219 971 253
rect 1005 219 1017 253
rect 959 185 1017 219
rect 959 151 971 185
rect 1005 151 1017 185
rect 959 117 1017 151
rect 959 83 971 117
rect 1005 83 1017 117
rect 959 68 1017 83
rect 1217 253 1275 268
rect 1217 219 1229 253
rect 1263 219 1275 253
rect 1217 185 1275 219
rect 1217 151 1229 185
rect 1263 151 1275 185
rect 1217 117 1275 151
rect 1217 83 1229 117
rect 1263 83 1275 117
rect 1217 68 1275 83
rect 1411 253 1469 268
rect 1411 219 1423 253
rect 1457 219 1469 253
rect 1411 185 1469 219
rect 1411 151 1423 185
rect 1457 151 1469 185
rect 1411 117 1469 151
rect 1411 83 1423 117
rect 1457 83 1469 117
rect 1411 68 1469 83
rect 1669 253 1727 268
rect 1669 219 1681 253
rect 1715 219 1727 253
rect 1669 185 1727 219
rect 1669 151 1681 185
rect 1715 151 1727 185
rect 1669 117 1727 151
rect 1669 83 1681 117
rect 1715 83 1727 117
rect 1669 68 1727 83
rect 1927 253 1985 268
rect 1927 219 1939 253
rect 1973 219 1985 253
rect 1927 185 1985 219
rect 1927 151 1939 185
rect 1973 151 1985 185
rect 1927 117 1985 151
rect 1927 83 1939 117
rect 1973 83 1985 117
rect 1927 68 1985 83
rect 2185 253 2243 268
rect 2185 219 2197 253
rect 2231 219 2243 253
rect 2185 185 2243 219
rect 2185 151 2197 185
rect 2231 151 2243 185
rect 2185 117 2243 151
rect 2185 83 2197 117
rect 2231 83 2243 117
rect 2185 68 2243 83
rect 2379 253 2437 268
rect 2379 219 2391 253
rect 2425 219 2437 253
rect 2379 185 2437 219
rect 2379 151 2391 185
rect 2425 151 2437 185
rect 2379 117 2437 151
rect 2379 83 2391 117
rect 2425 83 2437 117
rect 2379 68 2437 83
rect 2637 253 2695 268
rect 2637 219 2649 253
rect 2683 219 2695 253
rect 2637 185 2695 219
rect 2637 151 2649 185
rect 2683 151 2695 185
rect 2637 117 2695 151
rect 2637 83 2649 117
rect 2683 83 2695 117
rect 2637 68 2695 83
rect 959 -50 1017 -35
rect 959 -84 971 -50
rect 1005 -84 1017 -50
rect 959 -118 1017 -84
rect 959 -152 971 -118
rect 1005 -152 1017 -118
rect 959 -186 1017 -152
rect 959 -220 971 -186
rect 1005 -220 1017 -186
rect 959 -235 1017 -220
rect 1217 -50 1275 -35
rect 1217 -84 1229 -50
rect 1263 -84 1275 -50
rect 1217 -118 1275 -84
rect 1217 -152 1229 -118
rect 1263 -152 1275 -118
rect 1217 -186 1275 -152
rect 1217 -220 1229 -186
rect 1263 -220 1275 -186
rect 1217 -235 1275 -220
rect 1411 -50 1469 -35
rect 1411 -84 1423 -50
rect 1457 -84 1469 -50
rect 1411 -118 1469 -84
rect 1411 -152 1423 -118
rect 1457 -152 1469 -118
rect 1411 -186 1469 -152
rect 1411 -220 1423 -186
rect 1457 -220 1469 -186
rect 1411 -235 1469 -220
rect 1669 -50 1727 -35
rect 1669 -84 1681 -50
rect 1715 -84 1727 -50
rect 1669 -118 1727 -84
rect 1669 -152 1681 -118
rect 1715 -152 1727 -118
rect 1669 -186 1727 -152
rect 1669 -220 1681 -186
rect 1715 -220 1727 -186
rect 1669 -235 1727 -220
rect 1927 -50 1985 -35
rect 1927 -84 1939 -50
rect 1973 -84 1985 -50
rect 1927 -118 1985 -84
rect 1927 -152 1939 -118
rect 1973 -152 1985 -118
rect 1927 -186 1985 -152
rect 1927 -220 1939 -186
rect 1973 -220 1985 -186
rect 1927 -235 1985 -220
rect 2185 -50 2243 -35
rect 2185 -84 2197 -50
rect 2231 -84 2243 -50
rect 2185 -118 2243 -84
rect 2185 -152 2197 -118
rect 2231 -152 2243 -118
rect 2185 -186 2243 -152
rect 2185 -220 2197 -186
rect 2231 -220 2243 -186
rect 2185 -235 2243 -220
rect 2379 -50 2437 -35
rect 2379 -84 2391 -50
rect 2425 -84 2437 -50
rect 2379 -118 2437 -84
rect 2379 -152 2391 -118
rect 2425 -152 2437 -118
rect 2379 -186 2437 -152
rect 2379 -220 2391 -186
rect 2425 -220 2437 -186
rect 2379 -235 2437 -220
rect 2637 -50 2695 -35
rect 2637 -84 2649 -50
rect 2683 -84 2695 -50
rect 2637 -118 2695 -84
rect 2637 -152 2649 -118
rect 2683 -152 2695 -118
rect 2637 -186 2695 -152
rect 2637 -220 2649 -186
rect 2683 -220 2695 -186
rect 2637 -235 2695 -220
rect 959 -514 1017 -499
rect 959 -548 971 -514
rect 1005 -548 1017 -514
rect 959 -582 1017 -548
rect 959 -616 971 -582
rect 1005 -616 1017 -582
rect 959 -650 1017 -616
rect 959 -684 971 -650
rect 1005 -684 1017 -650
rect 959 -699 1017 -684
rect 1217 -514 1275 -499
rect 1217 -548 1229 -514
rect 1263 -548 1275 -514
rect 1217 -582 1275 -548
rect 1217 -616 1229 -582
rect 1263 -616 1275 -582
rect 1217 -650 1275 -616
rect 1217 -684 1229 -650
rect 1263 -684 1275 -650
rect 1217 -699 1275 -684
rect 1411 -514 1469 -499
rect 1411 -548 1423 -514
rect 1457 -548 1469 -514
rect 1411 -582 1469 -548
rect 1411 -616 1423 -582
rect 1457 -616 1469 -582
rect 1411 -650 1469 -616
rect 1411 -684 1423 -650
rect 1457 -684 1469 -650
rect 1411 -699 1469 -684
rect 1669 -514 1727 -499
rect 1669 -548 1681 -514
rect 1715 -548 1727 -514
rect 1669 -582 1727 -548
rect 1669 -616 1681 -582
rect 1715 -616 1727 -582
rect 1669 -650 1727 -616
rect 1669 -684 1681 -650
rect 1715 -684 1727 -650
rect 1669 -699 1727 -684
rect 1927 -514 1985 -499
rect 1927 -548 1939 -514
rect 1973 -548 1985 -514
rect 1927 -582 1985 -548
rect 1927 -616 1939 -582
rect 1973 -616 1985 -582
rect 1927 -650 1985 -616
rect 1927 -684 1939 -650
rect 1973 -684 1985 -650
rect 1927 -699 1985 -684
rect 2185 -514 2243 -499
rect 2185 -548 2197 -514
rect 2231 -548 2243 -514
rect 2185 -582 2243 -548
rect 2185 -616 2197 -582
rect 2231 -616 2243 -582
rect 2185 -650 2243 -616
rect 2185 -684 2197 -650
rect 2231 -684 2243 -650
rect 2185 -699 2243 -684
rect 2379 -514 2437 -499
rect 2379 -548 2391 -514
rect 2425 -548 2437 -514
rect 2379 -582 2437 -548
rect 2379 -616 2391 -582
rect 2425 -616 2437 -582
rect 2379 -650 2437 -616
rect 2379 -684 2391 -650
rect 2425 -684 2437 -650
rect 2379 -699 2437 -684
rect 2637 -514 2695 -499
rect 2637 -548 2649 -514
rect 2683 -548 2695 -514
rect 2637 -582 2695 -548
rect 2637 -616 2649 -582
rect 2683 -616 2695 -582
rect 2637 -650 2695 -616
rect 2637 -684 2649 -650
rect 2683 -684 2695 -650
rect 2637 -699 2695 -684
rect 959 -817 1017 -802
rect 959 -851 971 -817
rect 1005 -851 1017 -817
rect 959 -885 1017 -851
rect 959 -919 971 -885
rect 1005 -919 1017 -885
rect 959 -953 1017 -919
rect 959 -987 971 -953
rect 1005 -987 1017 -953
rect 959 -1002 1017 -987
rect 1217 -817 1275 -802
rect 1217 -851 1229 -817
rect 1263 -851 1275 -817
rect 1217 -885 1275 -851
rect 1217 -919 1229 -885
rect 1263 -919 1275 -885
rect 1217 -953 1275 -919
rect 1217 -987 1229 -953
rect 1263 -987 1275 -953
rect 1217 -1002 1275 -987
rect 1411 -817 1469 -802
rect 1411 -851 1423 -817
rect 1457 -851 1469 -817
rect 1411 -885 1469 -851
rect 1411 -919 1423 -885
rect 1457 -919 1469 -885
rect 1411 -953 1469 -919
rect 1411 -987 1423 -953
rect 1457 -987 1469 -953
rect 1411 -1002 1469 -987
rect 1669 -817 1727 -802
rect 1669 -851 1681 -817
rect 1715 -851 1727 -817
rect 1669 -885 1727 -851
rect 1669 -919 1681 -885
rect 1715 -919 1727 -885
rect 1669 -953 1727 -919
rect 1669 -987 1681 -953
rect 1715 -987 1727 -953
rect 1669 -1002 1727 -987
rect 1927 -817 1985 -802
rect 1927 -851 1939 -817
rect 1973 -851 1985 -817
rect 1927 -885 1985 -851
rect 1927 -919 1939 -885
rect 1973 -919 1985 -885
rect 1927 -953 1985 -919
rect 1927 -987 1939 -953
rect 1973 -987 1985 -953
rect 1927 -1002 1985 -987
rect 2185 -817 2243 -802
rect 2185 -851 2197 -817
rect 2231 -851 2243 -817
rect 2185 -885 2243 -851
rect 2185 -919 2197 -885
rect 2231 -919 2243 -885
rect 2185 -953 2243 -919
rect 2185 -987 2197 -953
rect 2231 -987 2243 -953
rect 2185 -1002 2243 -987
rect 2379 -817 2437 -802
rect 2379 -851 2391 -817
rect 2425 -851 2437 -817
rect 2379 -885 2437 -851
rect 2379 -919 2391 -885
rect 2425 -919 2437 -885
rect 2379 -953 2437 -919
rect 2379 -987 2391 -953
rect 2425 -987 2437 -953
rect 2379 -1002 2437 -987
rect 2637 -817 2695 -802
rect 2637 -851 2649 -817
rect 2683 -851 2695 -817
rect 2637 -885 2695 -851
rect 2637 -919 2649 -885
rect 2683 -919 2695 -885
rect 2637 -953 2695 -919
rect 2637 -987 2649 -953
rect 2683 -987 2695 -953
rect 2637 -1002 2695 -987
rect 959 -1281 1017 -1266
rect 959 -1315 971 -1281
rect 1005 -1315 1017 -1281
rect 959 -1349 1017 -1315
rect 959 -1383 971 -1349
rect 1005 -1383 1017 -1349
rect 959 -1417 1017 -1383
rect 959 -1451 971 -1417
rect 1005 -1451 1017 -1417
rect 959 -1466 1017 -1451
rect 1217 -1281 1275 -1266
rect 1217 -1315 1229 -1281
rect 1263 -1315 1275 -1281
rect 1217 -1349 1275 -1315
rect 1217 -1383 1229 -1349
rect 1263 -1383 1275 -1349
rect 1217 -1417 1275 -1383
rect 1217 -1451 1229 -1417
rect 1263 -1451 1275 -1417
rect 1217 -1466 1275 -1451
rect 1411 -1281 1469 -1266
rect 1411 -1315 1423 -1281
rect 1457 -1315 1469 -1281
rect 1411 -1349 1469 -1315
rect 1411 -1383 1423 -1349
rect 1457 -1383 1469 -1349
rect 1411 -1417 1469 -1383
rect 1411 -1451 1423 -1417
rect 1457 -1451 1469 -1417
rect 1411 -1466 1469 -1451
rect 1669 -1281 1727 -1266
rect 1669 -1315 1681 -1281
rect 1715 -1315 1727 -1281
rect 1669 -1349 1727 -1315
rect 1669 -1383 1681 -1349
rect 1715 -1383 1727 -1349
rect 1669 -1417 1727 -1383
rect 1669 -1451 1681 -1417
rect 1715 -1451 1727 -1417
rect 1669 -1466 1727 -1451
rect 1927 -1281 1985 -1266
rect 1927 -1315 1939 -1281
rect 1973 -1315 1985 -1281
rect 1927 -1349 1985 -1315
rect 1927 -1383 1939 -1349
rect 1973 -1383 1985 -1349
rect 1927 -1417 1985 -1383
rect 1927 -1451 1939 -1417
rect 1973 -1451 1985 -1417
rect 1927 -1466 1985 -1451
rect 2185 -1281 2243 -1266
rect 2185 -1315 2197 -1281
rect 2231 -1315 2243 -1281
rect 2185 -1349 2243 -1315
rect 2185 -1383 2197 -1349
rect 2231 -1383 2243 -1349
rect 2185 -1417 2243 -1383
rect 2185 -1451 2197 -1417
rect 2231 -1451 2243 -1417
rect 2185 -1466 2243 -1451
rect 2379 -1281 2437 -1266
rect 2379 -1315 2391 -1281
rect 2425 -1315 2437 -1281
rect 2379 -1349 2437 -1315
rect 2379 -1383 2391 -1349
rect 2425 -1383 2437 -1349
rect 2379 -1417 2437 -1383
rect 2379 -1451 2391 -1417
rect 2425 -1451 2437 -1417
rect 2379 -1466 2437 -1451
rect 2637 -1281 2695 -1266
rect 2637 -1315 2649 -1281
rect 2683 -1315 2695 -1281
rect 2637 -1349 2695 -1315
rect 2637 -1383 2649 -1349
rect 2683 -1383 2695 -1349
rect 2637 -1417 2695 -1383
rect 2637 -1451 2649 -1417
rect 2683 -1451 2695 -1417
rect 2637 -1466 2695 -1451
rect 959 -1584 1017 -1569
rect 959 -1618 971 -1584
rect 1005 -1618 1017 -1584
rect 959 -1652 1017 -1618
rect 959 -1686 971 -1652
rect 1005 -1686 1017 -1652
rect 959 -1720 1017 -1686
rect 959 -1754 971 -1720
rect 1005 -1754 1017 -1720
rect 959 -1769 1017 -1754
rect 1217 -1584 1275 -1569
rect 1217 -1618 1229 -1584
rect 1263 -1618 1275 -1584
rect 1217 -1652 1275 -1618
rect 1217 -1686 1229 -1652
rect 1263 -1686 1275 -1652
rect 1217 -1720 1275 -1686
rect 1217 -1754 1229 -1720
rect 1263 -1754 1275 -1720
rect 1217 -1769 1275 -1754
rect 1411 -1584 1469 -1569
rect 1411 -1618 1423 -1584
rect 1457 -1618 1469 -1584
rect 1411 -1652 1469 -1618
rect 1411 -1686 1423 -1652
rect 1457 -1686 1469 -1652
rect 1411 -1720 1469 -1686
rect 1411 -1754 1423 -1720
rect 1457 -1754 1469 -1720
rect 1411 -1769 1469 -1754
rect 1669 -1584 1727 -1569
rect 1669 -1618 1681 -1584
rect 1715 -1618 1727 -1584
rect 1669 -1652 1727 -1618
rect 1669 -1686 1681 -1652
rect 1715 -1686 1727 -1652
rect 1669 -1720 1727 -1686
rect 1669 -1754 1681 -1720
rect 1715 -1754 1727 -1720
rect 1669 -1769 1727 -1754
rect 1927 -1584 1985 -1569
rect 1927 -1618 1939 -1584
rect 1973 -1618 1985 -1584
rect 1927 -1652 1985 -1618
rect 1927 -1686 1939 -1652
rect 1973 -1686 1985 -1652
rect 1927 -1720 1985 -1686
rect 1927 -1754 1939 -1720
rect 1973 -1754 1985 -1720
rect 1927 -1769 1985 -1754
rect 2185 -1584 2243 -1569
rect 2185 -1618 2197 -1584
rect 2231 -1618 2243 -1584
rect 2185 -1652 2243 -1618
rect 2185 -1686 2197 -1652
rect 2231 -1686 2243 -1652
rect 2185 -1720 2243 -1686
rect 2185 -1754 2197 -1720
rect 2231 -1754 2243 -1720
rect 2185 -1769 2243 -1754
rect 2379 -1584 2437 -1569
rect 2379 -1618 2391 -1584
rect 2425 -1618 2437 -1584
rect 2379 -1652 2437 -1618
rect 2379 -1686 2391 -1652
rect 2425 -1686 2437 -1652
rect 2379 -1720 2437 -1686
rect 2379 -1754 2391 -1720
rect 2425 -1754 2437 -1720
rect 2379 -1769 2437 -1754
rect 2637 -1584 2695 -1569
rect 2637 -1618 2649 -1584
rect 2683 -1618 2695 -1584
rect 2637 -1652 2695 -1618
rect 2637 -1686 2649 -1652
rect 2683 -1686 2695 -1652
rect 2637 -1720 2695 -1686
rect 2637 -1754 2649 -1720
rect 2683 -1754 2695 -1720
rect 2637 -1769 2695 -1754
rect 959 -2054 1017 -2039
rect 959 -2088 971 -2054
rect 1005 -2088 1017 -2054
rect 959 -2122 1017 -2088
rect 959 -2156 971 -2122
rect 1005 -2156 1017 -2122
rect 959 -2190 1017 -2156
rect 959 -2224 971 -2190
rect 1005 -2224 1017 -2190
rect 959 -2239 1017 -2224
rect 1217 -2054 1275 -2039
rect 1217 -2088 1229 -2054
rect 1263 -2088 1275 -2054
rect 1217 -2122 1275 -2088
rect 1217 -2156 1229 -2122
rect 1263 -2156 1275 -2122
rect 1217 -2190 1275 -2156
rect 1217 -2224 1229 -2190
rect 1263 -2224 1275 -2190
rect 1217 -2239 1275 -2224
rect 1411 -2054 1469 -2039
rect 1411 -2088 1423 -2054
rect 1457 -2088 1469 -2054
rect 1411 -2122 1469 -2088
rect 1411 -2156 1423 -2122
rect 1457 -2156 1469 -2122
rect 1411 -2190 1469 -2156
rect 1411 -2224 1423 -2190
rect 1457 -2224 1469 -2190
rect 1411 -2239 1469 -2224
rect 1669 -2054 1727 -2039
rect 1669 -2088 1681 -2054
rect 1715 -2088 1727 -2054
rect 1669 -2122 1727 -2088
rect 1669 -2156 1681 -2122
rect 1715 -2156 1727 -2122
rect 1669 -2190 1727 -2156
rect 1669 -2224 1681 -2190
rect 1715 -2224 1727 -2190
rect 1669 -2239 1727 -2224
rect 1927 -2054 1985 -2039
rect 1927 -2088 1939 -2054
rect 1973 -2088 1985 -2054
rect 1927 -2122 1985 -2088
rect 1927 -2156 1939 -2122
rect 1973 -2156 1985 -2122
rect 1927 -2190 1985 -2156
rect 1927 -2224 1939 -2190
rect 1973 -2224 1985 -2190
rect 1927 -2239 1985 -2224
rect 2185 -2054 2243 -2039
rect 2185 -2088 2197 -2054
rect 2231 -2088 2243 -2054
rect 2185 -2122 2243 -2088
rect 2185 -2156 2197 -2122
rect 2231 -2156 2243 -2122
rect 2185 -2190 2243 -2156
rect 2185 -2224 2197 -2190
rect 2231 -2224 2243 -2190
rect 2185 -2239 2243 -2224
rect 2379 -2054 2437 -2039
rect 2379 -2088 2391 -2054
rect 2425 -2088 2437 -2054
rect 2379 -2122 2437 -2088
rect 2379 -2156 2391 -2122
rect 2425 -2156 2437 -2122
rect 2379 -2190 2437 -2156
rect 2379 -2224 2391 -2190
rect 2425 -2224 2437 -2190
rect 2379 -2239 2437 -2224
rect 2637 -2054 2695 -2039
rect 2637 -2088 2649 -2054
rect 2683 -2088 2695 -2054
rect 2637 -2122 2695 -2088
rect 2637 -2156 2649 -2122
rect 2683 -2156 2695 -2122
rect 2637 -2190 2695 -2156
rect 2637 -2224 2649 -2190
rect 2683 -2224 2695 -2190
rect 2637 -2239 2695 -2224
<< pdiffc >>
rect 971 219 1005 253
rect 971 151 1005 185
rect 971 83 1005 117
rect 1229 219 1263 253
rect 1229 151 1263 185
rect 1229 83 1263 117
rect 1423 219 1457 253
rect 1423 151 1457 185
rect 1423 83 1457 117
rect 1681 219 1715 253
rect 1681 151 1715 185
rect 1681 83 1715 117
rect 1939 219 1973 253
rect 1939 151 1973 185
rect 1939 83 1973 117
rect 2197 219 2231 253
rect 2197 151 2231 185
rect 2197 83 2231 117
rect 2391 219 2425 253
rect 2391 151 2425 185
rect 2391 83 2425 117
rect 2649 219 2683 253
rect 2649 151 2683 185
rect 2649 83 2683 117
rect 971 -84 1005 -50
rect 971 -152 1005 -118
rect 971 -220 1005 -186
rect 1229 -84 1263 -50
rect 1229 -152 1263 -118
rect 1229 -220 1263 -186
rect 1423 -84 1457 -50
rect 1423 -152 1457 -118
rect 1423 -220 1457 -186
rect 1681 -84 1715 -50
rect 1681 -152 1715 -118
rect 1681 -220 1715 -186
rect 1939 -84 1973 -50
rect 1939 -152 1973 -118
rect 1939 -220 1973 -186
rect 2197 -84 2231 -50
rect 2197 -152 2231 -118
rect 2197 -220 2231 -186
rect 2391 -84 2425 -50
rect 2391 -152 2425 -118
rect 2391 -220 2425 -186
rect 2649 -84 2683 -50
rect 2649 -152 2683 -118
rect 2649 -220 2683 -186
rect 971 -548 1005 -514
rect 971 -616 1005 -582
rect 971 -684 1005 -650
rect 1229 -548 1263 -514
rect 1229 -616 1263 -582
rect 1229 -684 1263 -650
rect 1423 -548 1457 -514
rect 1423 -616 1457 -582
rect 1423 -684 1457 -650
rect 1681 -548 1715 -514
rect 1681 -616 1715 -582
rect 1681 -684 1715 -650
rect 1939 -548 1973 -514
rect 1939 -616 1973 -582
rect 1939 -684 1973 -650
rect 2197 -548 2231 -514
rect 2197 -616 2231 -582
rect 2197 -684 2231 -650
rect 2391 -548 2425 -514
rect 2391 -616 2425 -582
rect 2391 -684 2425 -650
rect 2649 -548 2683 -514
rect 2649 -616 2683 -582
rect 2649 -684 2683 -650
rect 971 -851 1005 -817
rect 971 -919 1005 -885
rect 971 -987 1005 -953
rect 1229 -851 1263 -817
rect 1229 -919 1263 -885
rect 1229 -987 1263 -953
rect 1423 -851 1457 -817
rect 1423 -919 1457 -885
rect 1423 -987 1457 -953
rect 1681 -851 1715 -817
rect 1681 -919 1715 -885
rect 1681 -987 1715 -953
rect 1939 -851 1973 -817
rect 1939 -919 1973 -885
rect 1939 -987 1973 -953
rect 2197 -851 2231 -817
rect 2197 -919 2231 -885
rect 2197 -987 2231 -953
rect 2391 -851 2425 -817
rect 2391 -919 2425 -885
rect 2391 -987 2425 -953
rect 2649 -851 2683 -817
rect 2649 -919 2683 -885
rect 2649 -987 2683 -953
rect 971 -1315 1005 -1281
rect 971 -1383 1005 -1349
rect 971 -1451 1005 -1417
rect 1229 -1315 1263 -1281
rect 1229 -1383 1263 -1349
rect 1229 -1451 1263 -1417
rect 1423 -1315 1457 -1281
rect 1423 -1383 1457 -1349
rect 1423 -1451 1457 -1417
rect 1681 -1315 1715 -1281
rect 1681 -1383 1715 -1349
rect 1681 -1451 1715 -1417
rect 1939 -1315 1973 -1281
rect 1939 -1383 1973 -1349
rect 1939 -1451 1973 -1417
rect 2197 -1315 2231 -1281
rect 2197 -1383 2231 -1349
rect 2197 -1451 2231 -1417
rect 2391 -1315 2425 -1281
rect 2391 -1383 2425 -1349
rect 2391 -1451 2425 -1417
rect 2649 -1315 2683 -1281
rect 2649 -1383 2683 -1349
rect 2649 -1451 2683 -1417
rect 971 -1618 1005 -1584
rect 971 -1686 1005 -1652
rect 971 -1754 1005 -1720
rect 1229 -1618 1263 -1584
rect 1229 -1686 1263 -1652
rect 1229 -1754 1263 -1720
rect 1423 -1618 1457 -1584
rect 1423 -1686 1457 -1652
rect 1423 -1754 1457 -1720
rect 1681 -1618 1715 -1584
rect 1681 -1686 1715 -1652
rect 1681 -1754 1715 -1720
rect 1939 -1618 1973 -1584
rect 1939 -1686 1973 -1652
rect 1939 -1754 1973 -1720
rect 2197 -1618 2231 -1584
rect 2197 -1686 2231 -1652
rect 2197 -1754 2231 -1720
rect 2391 -1618 2425 -1584
rect 2391 -1686 2425 -1652
rect 2391 -1754 2425 -1720
rect 2649 -1618 2683 -1584
rect 2649 -1686 2683 -1652
rect 2649 -1754 2683 -1720
rect 971 -2088 1005 -2054
rect 971 -2156 1005 -2122
rect 971 -2224 1005 -2190
rect 1229 -2088 1263 -2054
rect 1229 -2156 1263 -2122
rect 1229 -2224 1263 -2190
rect 1423 -2088 1457 -2054
rect 1423 -2156 1457 -2122
rect 1423 -2224 1457 -2190
rect 1681 -2088 1715 -2054
rect 1681 -2156 1715 -2122
rect 1681 -2224 1715 -2190
rect 1939 -2088 1973 -2054
rect 1939 -2156 1973 -2122
rect 1939 -2224 1973 -2190
rect 2197 -2088 2231 -2054
rect 2197 -2156 2231 -2122
rect 2197 -2224 2231 -2190
rect 2391 -2088 2425 -2054
rect 2391 -2156 2425 -2122
rect 2391 -2224 2425 -2190
rect 2649 -2088 2683 -2054
rect 2649 -2156 2683 -2122
rect 2649 -2224 2683 -2190
<< nsubdiff >>
rect 856 429 977 463
rect 1011 429 1045 463
rect 1079 429 1113 463
rect 1147 429 1181 463
rect 1215 429 1249 463
rect 1283 429 1317 463
rect 1351 429 1385 463
rect 1419 429 1453 463
rect 1487 429 1521 463
rect 1555 429 1589 463
rect 1623 429 1657 463
rect 1691 429 1725 463
rect 1759 429 1793 463
rect 1827 429 1861 463
rect 1895 429 1929 463
rect 1963 429 1997 463
rect 2031 429 2065 463
rect 2099 429 2133 463
rect 2167 429 2201 463
rect 2235 429 2269 463
rect 2303 429 2337 463
rect 2371 429 2405 463
rect 2439 429 2473 463
rect 2507 429 2541 463
rect 2575 429 2609 463
rect 2643 429 2793 463
rect 856 342 890 429
rect 856 274 890 308
rect 2759 342 2793 429
rect 2759 274 2793 308
rect 856 206 890 240
rect 856 138 890 172
rect 856 70 890 104
rect 2759 206 2793 240
rect 2759 138 2793 172
rect 2759 70 2793 104
rect 856 2 890 36
rect 2759 2 2793 36
rect 856 -66 890 -32
rect 856 -134 890 -100
rect 856 -202 890 -168
rect 2759 -66 2793 -32
rect 2759 -134 2793 -100
rect 2759 -202 2793 -168
rect 856 -270 890 -236
rect 856 -338 890 -304
rect 2759 -270 2793 -236
rect 856 -406 890 -372
rect 2759 -338 2793 -304
rect 856 -474 890 -440
rect 2759 -406 2793 -372
rect 2759 -474 2793 -440
rect 856 -542 890 -508
rect 856 -610 890 -576
rect 856 -678 890 -644
rect 2759 -542 2793 -508
rect 2759 -610 2793 -576
rect 2759 -678 2793 -644
rect 856 -746 890 -712
rect 2759 -746 2793 -712
rect 856 -814 890 -780
rect 856 -882 890 -848
rect 856 -950 890 -916
rect 856 -1018 890 -984
rect 2759 -814 2793 -780
rect 2759 -882 2793 -848
rect 2759 -950 2793 -916
rect 856 -1086 890 -1052
rect 2759 -1018 2793 -984
rect 2759 -1086 2793 -1052
rect 856 -1154 890 -1120
rect 2759 -1154 2793 -1120
rect 856 -1222 890 -1188
rect 856 -1290 890 -1256
rect 2759 -1222 2793 -1188
rect 856 -1358 890 -1324
rect 856 -1426 890 -1392
rect 856 -1494 890 -1460
rect 2759 -1290 2793 -1256
rect 2759 -1358 2793 -1324
rect 2759 -1426 2793 -1392
rect 856 -1562 890 -1528
rect 2759 -1494 2793 -1460
rect 2759 -1562 2793 -1528
rect 856 -1630 890 -1596
rect 856 -1698 890 -1664
rect 856 -1766 890 -1732
rect 2759 -1630 2793 -1596
rect 2759 -1698 2793 -1664
rect 2759 -1766 2793 -1732
rect 856 -1834 890 -1800
rect 2759 -1834 2793 -1800
rect 856 -1902 890 -1868
rect 856 -1970 890 -1936
rect 2759 -1902 2793 -1868
rect 856 -2038 890 -2004
rect 2759 -1970 2793 -1936
rect 2759 -2038 2793 -2004
rect 856 -2106 890 -2072
rect 856 -2174 890 -2140
rect 856 -2310 890 -2208
rect 2759 -2106 2793 -2072
rect 2759 -2174 2793 -2140
rect 2759 -2310 2793 -2208
rect 856 -2344 977 -2310
rect 1011 -2344 1045 -2310
rect 1079 -2344 1113 -2310
rect 1147 -2344 1181 -2310
rect 1215 -2344 1249 -2310
rect 1283 -2344 1317 -2310
rect 1351 -2344 1385 -2310
rect 1419 -2344 1453 -2310
rect 1487 -2344 1521 -2310
rect 1555 -2344 1589 -2310
rect 1623 -2344 1657 -2310
rect 1691 -2344 1725 -2310
rect 1759 -2344 1793 -2310
rect 1827 -2344 1861 -2310
rect 1895 -2344 1929 -2310
rect 1963 -2344 1997 -2310
rect 2031 -2344 2065 -2310
rect 2099 -2344 2133 -2310
rect 2167 -2344 2201 -2310
rect 2235 -2344 2269 -2310
rect 2303 -2344 2337 -2310
rect 2371 -2344 2405 -2310
rect 2439 -2344 2473 -2310
rect 2507 -2344 2541 -2310
rect 2575 -2344 2609 -2310
rect 2643 -2344 2793 -2310
<< nsubdiffcont >>
rect 977 429 1011 463
rect 1045 429 1079 463
rect 1113 429 1147 463
rect 1181 429 1215 463
rect 1249 429 1283 463
rect 1317 429 1351 463
rect 1385 429 1419 463
rect 1453 429 1487 463
rect 1521 429 1555 463
rect 1589 429 1623 463
rect 1657 429 1691 463
rect 1725 429 1759 463
rect 1793 429 1827 463
rect 1861 429 1895 463
rect 1929 429 1963 463
rect 1997 429 2031 463
rect 2065 429 2099 463
rect 2133 429 2167 463
rect 2201 429 2235 463
rect 2269 429 2303 463
rect 2337 429 2371 463
rect 2405 429 2439 463
rect 2473 429 2507 463
rect 2541 429 2575 463
rect 2609 429 2643 463
rect 856 308 890 342
rect 856 240 890 274
rect 2759 308 2793 342
rect 856 172 890 206
rect 856 104 890 138
rect 856 36 890 70
rect 2759 240 2793 274
rect 2759 172 2793 206
rect 2759 104 2793 138
rect 856 -32 890 2
rect 2759 36 2793 70
rect 2759 -32 2793 2
rect 856 -100 890 -66
rect 856 -168 890 -134
rect 856 -236 890 -202
rect 2759 -100 2793 -66
rect 2759 -168 2793 -134
rect 856 -304 890 -270
rect 2759 -236 2793 -202
rect 2759 -304 2793 -270
rect 856 -372 890 -338
rect 2759 -372 2793 -338
rect 856 -440 890 -406
rect 856 -508 890 -474
rect 2759 -440 2793 -406
rect 856 -576 890 -542
rect 856 -644 890 -610
rect 856 -712 890 -678
rect 2759 -508 2793 -474
rect 2759 -576 2793 -542
rect 2759 -644 2793 -610
rect 2759 -712 2793 -678
rect 856 -780 890 -746
rect 2759 -780 2793 -746
rect 856 -848 890 -814
rect 856 -916 890 -882
rect 856 -984 890 -950
rect 2759 -848 2793 -814
rect 2759 -916 2793 -882
rect 2759 -984 2793 -950
rect 856 -1052 890 -1018
rect 856 -1120 890 -1086
rect 2759 -1052 2793 -1018
rect 856 -1188 890 -1154
rect 2759 -1120 2793 -1086
rect 856 -1256 890 -1222
rect 2759 -1188 2793 -1154
rect 2759 -1256 2793 -1222
rect 856 -1324 890 -1290
rect 856 -1392 890 -1358
rect 856 -1460 890 -1426
rect 2759 -1324 2793 -1290
rect 2759 -1392 2793 -1358
rect 2759 -1460 2793 -1426
rect 856 -1528 890 -1494
rect 2759 -1528 2793 -1494
rect 856 -1596 890 -1562
rect 856 -1664 890 -1630
rect 856 -1732 890 -1698
rect 856 -1800 890 -1766
rect 2759 -1596 2793 -1562
rect 2759 -1664 2793 -1630
rect 2759 -1732 2793 -1698
rect 856 -1868 890 -1834
rect 2759 -1800 2793 -1766
rect 856 -1936 890 -1902
rect 2759 -1868 2793 -1834
rect 2759 -1936 2793 -1902
rect 856 -2004 890 -1970
rect 856 -2072 890 -2038
rect 2759 -2004 2793 -1970
rect 856 -2140 890 -2106
rect 856 -2208 890 -2174
rect 2759 -2072 2793 -2038
rect 2759 -2140 2793 -2106
rect 2759 -2208 2793 -2174
rect 977 -2344 1011 -2310
rect 1045 -2344 1079 -2310
rect 1113 -2344 1147 -2310
rect 1181 -2344 1215 -2310
rect 1249 -2344 1283 -2310
rect 1317 -2344 1351 -2310
rect 1385 -2344 1419 -2310
rect 1453 -2344 1487 -2310
rect 1521 -2344 1555 -2310
rect 1589 -2344 1623 -2310
rect 1657 -2344 1691 -2310
rect 1725 -2344 1759 -2310
rect 1793 -2344 1827 -2310
rect 1861 -2344 1895 -2310
rect 1929 -2344 1963 -2310
rect 1997 -2344 2031 -2310
rect 2065 -2344 2099 -2310
rect 2133 -2344 2167 -2310
rect 2201 -2344 2235 -2310
rect 2269 -2344 2303 -2310
rect 2337 -2344 2371 -2310
rect 2405 -2344 2439 -2310
rect 2473 -2344 2507 -2310
rect 2541 -2344 2575 -2310
rect 2609 -2344 2643 -2310
<< poly >>
rect 1017 349 1217 365
rect 1017 315 1066 349
rect 1100 315 1134 349
rect 1168 315 1217 349
rect 1017 268 1217 315
rect 1469 349 1669 365
rect 1469 315 1518 349
rect 1552 315 1586 349
rect 1620 315 1669 349
rect 1469 268 1669 315
rect 1727 349 1927 365
rect 1727 315 1776 349
rect 1810 315 1844 349
rect 1878 315 1927 349
rect 1727 268 1927 315
rect 1985 349 2185 365
rect 1985 315 2034 349
rect 2068 315 2102 349
rect 2136 315 2185 349
rect 1985 268 2185 315
rect 2437 349 2637 365
rect 2437 315 2486 349
rect 2520 315 2554 349
rect 2588 315 2637 349
rect 2437 268 2637 315
rect 1017 42 1217 68
rect 1469 42 1669 68
rect 1727 42 1927 68
rect 1985 42 2185 68
rect 2437 42 2637 68
rect 1017 -35 1217 -9
rect 1469 -35 1669 -9
rect 1727 -35 1927 -9
rect 1985 -35 2185 -9
rect 2437 -35 2637 -9
rect 1017 -282 1217 -235
rect 1017 -316 1066 -282
rect 1100 -316 1134 -282
rect 1168 -316 1217 -282
rect 1017 -332 1217 -316
rect 1469 -282 1669 -235
rect 1469 -316 1518 -282
rect 1552 -316 1586 -282
rect 1620 -316 1669 -282
rect 1469 -332 1669 -316
rect 1727 -282 1927 -235
rect 1727 -316 1776 -282
rect 1810 -316 1844 -282
rect 1878 -316 1927 -282
rect 1727 -332 1927 -316
rect 1985 -282 2185 -235
rect 1985 -316 2034 -282
rect 2068 -316 2102 -282
rect 2136 -316 2185 -282
rect 1985 -332 2185 -316
rect 2437 -282 2637 -235
rect 2437 -316 2486 -282
rect 2520 -316 2554 -282
rect 2588 -316 2637 -282
rect 2437 -332 2637 -316
rect 1017 -418 1217 -402
rect 1017 -452 1066 -418
rect 1100 -452 1134 -418
rect 1168 -452 1217 -418
rect 1017 -499 1217 -452
rect 1469 -418 1669 -402
rect 1469 -452 1518 -418
rect 1552 -452 1586 -418
rect 1620 -452 1669 -418
rect 1469 -499 1669 -452
rect 1727 -418 1927 -402
rect 1727 -452 1776 -418
rect 1810 -452 1844 -418
rect 1878 -452 1927 -418
rect 1727 -499 1927 -452
rect 1985 -418 2185 -402
rect 1985 -452 2034 -418
rect 2068 -452 2102 -418
rect 2136 -452 2185 -418
rect 1985 -499 2185 -452
rect 2437 -418 2637 -402
rect 2437 -452 2486 -418
rect 2520 -452 2554 -418
rect 2588 -452 2637 -418
rect 2437 -499 2637 -452
rect 1017 -725 1217 -699
rect 1469 -725 1669 -699
rect 1727 -725 1927 -699
rect 1985 -725 2185 -699
rect 2437 -725 2637 -699
rect 1017 -802 1217 -776
rect 1469 -802 1669 -776
rect 1727 -802 1927 -776
rect 1985 -802 2185 -776
rect 2437 -802 2637 -776
rect 1017 -1049 1217 -1002
rect 1017 -1083 1066 -1049
rect 1100 -1083 1134 -1049
rect 1168 -1083 1217 -1049
rect 1017 -1099 1217 -1083
rect 1469 -1049 1669 -1002
rect 1469 -1083 1518 -1049
rect 1552 -1083 1586 -1049
rect 1620 -1083 1669 -1049
rect 1469 -1099 1669 -1083
rect 1727 -1049 1927 -1002
rect 1727 -1083 1776 -1049
rect 1810 -1083 1844 -1049
rect 1878 -1083 1927 -1049
rect 1727 -1099 1927 -1083
rect 1985 -1049 2185 -1002
rect 1985 -1083 2034 -1049
rect 2068 -1083 2102 -1049
rect 2136 -1083 2185 -1049
rect 1985 -1099 2185 -1083
rect 2437 -1049 2637 -1002
rect 2437 -1083 2486 -1049
rect 2520 -1083 2554 -1049
rect 2588 -1083 2637 -1049
rect 2437 -1099 2637 -1083
rect 1017 -1185 1217 -1169
rect 1017 -1219 1066 -1185
rect 1100 -1219 1134 -1185
rect 1168 -1219 1217 -1185
rect 1017 -1266 1217 -1219
rect 1469 -1185 1669 -1169
rect 1469 -1219 1518 -1185
rect 1552 -1219 1586 -1185
rect 1620 -1219 1669 -1185
rect 1469 -1266 1669 -1219
rect 1727 -1185 1927 -1169
rect 1727 -1219 1776 -1185
rect 1810 -1219 1844 -1185
rect 1878 -1219 1927 -1185
rect 1727 -1266 1927 -1219
rect 1985 -1185 2185 -1169
rect 1985 -1219 2034 -1185
rect 2068 -1219 2102 -1185
rect 2136 -1219 2185 -1185
rect 1985 -1266 2185 -1219
rect 2437 -1185 2637 -1169
rect 2437 -1219 2486 -1185
rect 2520 -1219 2554 -1185
rect 2588 -1219 2637 -1185
rect 2437 -1266 2637 -1219
rect 1017 -1492 1217 -1466
rect 1469 -1492 1669 -1466
rect 1727 -1492 1927 -1466
rect 1985 -1492 2185 -1466
rect 2437 -1492 2637 -1466
rect 1017 -1569 1217 -1543
rect 1469 -1569 1669 -1543
rect 1727 -1569 1927 -1543
rect 1985 -1569 2185 -1543
rect 2437 -1569 2637 -1543
rect 1017 -1816 1217 -1769
rect 1017 -1850 1066 -1816
rect 1100 -1850 1134 -1816
rect 1168 -1850 1217 -1816
rect 1017 -1866 1217 -1850
rect 1469 -1816 1669 -1769
rect 1469 -1850 1518 -1816
rect 1552 -1850 1586 -1816
rect 1620 -1850 1669 -1816
rect 1469 -1866 1669 -1850
rect 1727 -1816 1927 -1769
rect 1727 -1850 1776 -1816
rect 1810 -1850 1844 -1816
rect 1878 -1850 1927 -1816
rect 1727 -1866 1927 -1850
rect 1985 -1816 2185 -1769
rect 1985 -1850 2034 -1816
rect 2068 -1850 2102 -1816
rect 2136 -1850 2185 -1816
rect 1985 -1866 2185 -1850
rect 2437 -1816 2637 -1769
rect 2437 -1850 2486 -1816
rect 2520 -1850 2554 -1816
rect 2588 -1850 2637 -1816
rect 2437 -1866 2637 -1850
rect 1017 -1958 1217 -1942
rect 1017 -1992 1066 -1958
rect 1100 -1992 1134 -1958
rect 1168 -1992 1217 -1958
rect 1017 -2039 1217 -1992
rect 1469 -1958 1669 -1942
rect 1469 -1992 1518 -1958
rect 1552 -1992 1586 -1958
rect 1620 -1992 1669 -1958
rect 1469 -2039 1669 -1992
rect 1727 -1958 1927 -1942
rect 1727 -1992 1776 -1958
rect 1810 -1992 1844 -1958
rect 1878 -1992 1927 -1958
rect 1727 -2039 1927 -1992
rect 1985 -1958 2185 -1942
rect 1985 -1992 2034 -1958
rect 2068 -1992 2102 -1958
rect 2136 -1992 2185 -1958
rect 1985 -2039 2185 -1992
rect 2437 -1958 2637 -1942
rect 2437 -1992 2486 -1958
rect 2520 -1992 2554 -1958
rect 2588 -1992 2637 -1958
rect 2437 -2039 2637 -1992
rect 1017 -2265 1217 -2239
rect 1469 -2265 1669 -2239
rect 1727 -2265 1927 -2239
rect 1985 -2265 2185 -2239
rect 2437 -2265 2637 -2239
<< polycont >>
rect 1066 315 1100 349
rect 1134 315 1168 349
rect 1518 315 1552 349
rect 1586 315 1620 349
rect 1776 315 1810 349
rect 1844 315 1878 349
rect 2034 315 2068 349
rect 2102 315 2136 349
rect 2486 315 2520 349
rect 2554 315 2588 349
rect 1066 -316 1100 -282
rect 1134 -316 1168 -282
rect 1518 -316 1552 -282
rect 1586 -316 1620 -282
rect 1776 -316 1810 -282
rect 1844 -316 1878 -282
rect 2034 -316 2068 -282
rect 2102 -316 2136 -282
rect 2486 -316 2520 -282
rect 2554 -316 2588 -282
rect 1066 -452 1100 -418
rect 1134 -452 1168 -418
rect 1518 -452 1552 -418
rect 1586 -452 1620 -418
rect 1776 -452 1810 -418
rect 1844 -452 1878 -418
rect 2034 -452 2068 -418
rect 2102 -452 2136 -418
rect 2486 -452 2520 -418
rect 2554 -452 2588 -418
rect 1066 -1083 1100 -1049
rect 1134 -1083 1168 -1049
rect 1518 -1083 1552 -1049
rect 1586 -1083 1620 -1049
rect 1776 -1083 1810 -1049
rect 1844 -1083 1878 -1049
rect 2034 -1083 2068 -1049
rect 2102 -1083 2136 -1049
rect 2486 -1083 2520 -1049
rect 2554 -1083 2588 -1049
rect 1066 -1219 1100 -1185
rect 1134 -1219 1168 -1185
rect 1518 -1219 1552 -1185
rect 1586 -1219 1620 -1185
rect 1776 -1219 1810 -1185
rect 1844 -1219 1878 -1185
rect 2034 -1219 2068 -1185
rect 2102 -1219 2136 -1185
rect 2486 -1219 2520 -1185
rect 2554 -1219 2588 -1185
rect 1066 -1850 1100 -1816
rect 1134 -1850 1168 -1816
rect 1518 -1850 1552 -1816
rect 1586 -1850 1620 -1816
rect 1776 -1850 1810 -1816
rect 1844 -1850 1878 -1816
rect 2034 -1850 2068 -1816
rect 2102 -1850 2136 -1816
rect 2486 -1850 2520 -1816
rect 2554 -1850 2588 -1816
rect 1066 -1992 1100 -1958
rect 1134 -1992 1168 -1958
rect 1518 -1992 1552 -1958
rect 1586 -1992 1620 -1958
rect 1776 -1992 1810 -1958
rect 1844 -1992 1878 -1958
rect 2034 -1992 2068 -1958
rect 2102 -1992 2136 -1958
rect 2486 -1992 2520 -1958
rect 2554 -1992 2588 -1958
<< locali >>
rect 856 429 977 463
rect 1036 429 1045 463
rect 1108 429 1113 463
rect 1180 429 1181 463
rect 1215 429 1218 463
rect 1283 429 1290 463
rect 1351 429 1362 463
rect 1419 429 1434 463
rect 1487 429 1506 463
rect 1555 429 1578 463
rect 1623 429 1650 463
rect 1691 429 1722 463
rect 1759 429 1793 463
rect 1828 429 1861 463
rect 1900 429 1929 463
rect 1972 429 1997 463
rect 2044 429 2065 463
rect 2116 429 2133 463
rect 2188 429 2201 463
rect 2260 429 2269 463
rect 2332 429 2337 463
rect 2404 429 2405 463
rect 2439 429 2442 463
rect 2507 429 2514 463
rect 2575 429 2586 463
rect 2643 429 2793 463
rect 856 342 890 429
rect 1017 315 1064 349
rect 1100 315 1134 349
rect 1170 315 1217 349
rect 1469 315 1516 349
rect 1552 315 1586 349
rect 1622 315 1669 349
rect 1727 315 1774 349
rect 1810 315 1844 349
rect 1880 315 1927 349
rect 1985 315 2032 349
rect 2068 315 2102 349
rect 2138 315 2185 349
rect 2437 315 2484 349
rect 2520 315 2554 349
rect 2590 315 2637 349
rect 2759 342 2793 429
rect 856 274 890 282
rect 2759 274 2793 282
rect 856 206 890 210
rect 856 100 890 104
rect 971 253 1005 272
rect 971 185 1005 187
rect 971 149 1005 151
rect 971 64 1005 83
rect 1229 253 1263 272
rect 1229 185 1263 187
rect 1229 149 1263 151
rect 1229 64 1263 83
rect 1423 253 1457 272
rect 1423 185 1457 187
rect 1423 149 1457 151
rect 1423 64 1457 83
rect 1681 253 1715 272
rect 1681 185 1715 187
rect 1681 149 1715 151
rect 1681 64 1715 83
rect 1939 253 1973 272
rect 1939 185 1973 187
rect 1939 149 1973 151
rect 1939 64 1973 83
rect 2197 253 2231 272
rect 2197 185 2231 187
rect 2197 149 2231 151
rect 2197 64 2231 83
rect 2391 253 2425 272
rect 2391 185 2425 187
rect 2391 149 2425 151
rect 2391 64 2425 83
rect 2649 253 2683 272
rect 2649 185 2683 187
rect 2649 149 2683 151
rect 2649 64 2683 83
rect 2759 206 2793 210
rect 2759 100 2793 104
rect 856 28 890 36
rect 2759 28 2793 36
rect 856 -44 890 -32
rect 856 -116 890 -100
rect 856 -188 890 -168
rect 856 -260 890 -236
rect 971 -50 1005 -31
rect 971 -118 1005 -116
rect 971 -154 1005 -152
rect 971 -239 1005 -220
rect 1229 -50 1263 -31
rect 1229 -118 1263 -116
rect 1229 -154 1263 -152
rect 1229 -239 1263 -220
rect 1423 -50 1457 -31
rect 1423 -118 1457 -116
rect 1423 -154 1457 -152
rect 1423 -239 1457 -220
rect 1681 -50 1715 -31
rect 1681 -118 1715 -116
rect 1681 -154 1715 -152
rect 1681 -239 1715 -220
rect 1939 -50 1973 -31
rect 1939 -118 1973 -116
rect 1939 -154 1973 -152
rect 1939 -239 1973 -220
rect 2197 -50 2231 -31
rect 2197 -118 2231 -116
rect 2197 -154 2231 -152
rect 2197 -239 2231 -220
rect 2391 -50 2425 -31
rect 2391 -118 2425 -116
rect 2391 -154 2425 -152
rect 2391 -239 2425 -220
rect 2649 -50 2683 -31
rect 2649 -118 2683 -116
rect 2649 -154 2683 -152
rect 2649 -239 2683 -220
rect 2759 -44 2793 -32
rect 2759 -116 2793 -100
rect 2759 -188 2793 -168
rect 2759 -260 2793 -236
rect 856 -332 890 -304
rect 1017 -316 1064 -282
rect 1100 -316 1134 -282
rect 1170 -316 1217 -282
rect 1469 -316 1516 -282
rect 1552 -316 1586 -282
rect 1622 -316 1669 -282
rect 1727 -316 1774 -282
rect 1810 -316 1844 -282
rect 1880 -316 1927 -282
rect 1985 -316 2032 -282
rect 2068 -316 2102 -282
rect 2138 -316 2185 -282
rect 2437 -316 2484 -282
rect 2520 -316 2554 -282
rect 2590 -316 2637 -282
rect 856 -404 890 -372
rect 2759 -332 2793 -304
rect 2759 -404 2793 -372
rect 856 -474 890 -440
rect 1017 -452 1064 -418
rect 1100 -452 1134 -418
rect 1170 -452 1217 -418
rect 1469 -452 1516 -418
rect 1552 -452 1586 -418
rect 1622 -452 1669 -418
rect 1727 -452 1774 -418
rect 1810 -452 1844 -418
rect 1880 -452 1927 -418
rect 1985 -452 2032 -418
rect 2068 -452 2102 -418
rect 2138 -452 2185 -418
rect 2437 -452 2484 -418
rect 2520 -452 2554 -418
rect 2590 -452 2637 -418
rect 2759 -474 2793 -440
rect 856 -542 890 -510
rect 856 -610 890 -582
rect 856 -678 890 -654
rect 971 -514 1005 -495
rect 971 -582 1005 -580
rect 971 -618 1005 -616
rect 971 -703 1005 -684
rect 1229 -514 1263 -495
rect 1229 -582 1263 -580
rect 1229 -618 1263 -616
rect 1229 -703 1263 -684
rect 1423 -514 1457 -495
rect 1423 -582 1457 -580
rect 1423 -618 1457 -616
rect 1423 -703 1457 -684
rect 1681 -514 1715 -495
rect 1681 -582 1715 -580
rect 1681 -618 1715 -616
rect 1681 -703 1715 -684
rect 1939 -514 1973 -495
rect 1939 -582 1973 -580
rect 1939 -618 1973 -616
rect 1939 -703 1973 -684
rect 2197 -514 2231 -495
rect 2197 -582 2231 -580
rect 2197 -618 2231 -616
rect 2197 -703 2231 -684
rect 2391 -514 2425 -495
rect 2391 -582 2425 -580
rect 2391 -618 2425 -616
rect 2391 -703 2425 -684
rect 2649 -514 2683 -495
rect 2649 -582 2683 -580
rect 2649 -618 2683 -616
rect 2649 -703 2683 -684
rect 2759 -542 2793 -510
rect 2759 -610 2793 -582
rect 2759 -678 2793 -654
rect 856 -746 890 -726
rect 2759 -746 2793 -726
rect 856 -814 890 -798
rect 856 -882 890 -870
rect 856 -950 890 -942
rect 971 -817 1005 -798
rect 971 -885 1005 -883
rect 971 -921 1005 -919
rect 971 -1006 1005 -987
rect 1229 -817 1263 -798
rect 1229 -885 1263 -883
rect 1229 -921 1263 -919
rect 1229 -1006 1263 -987
rect 1423 -817 1457 -798
rect 1423 -885 1457 -883
rect 1423 -921 1457 -919
rect 1423 -1006 1457 -987
rect 1681 -817 1715 -798
rect 1681 -885 1715 -883
rect 1681 -921 1715 -919
rect 1681 -1006 1715 -987
rect 1939 -817 1973 -798
rect 1939 -885 1973 -883
rect 1939 -921 1973 -919
rect 1939 -1006 1973 -987
rect 2197 -817 2231 -798
rect 2197 -885 2231 -883
rect 2197 -921 2231 -919
rect 2197 -1006 2231 -987
rect 2391 -817 2425 -798
rect 2391 -885 2425 -883
rect 2391 -921 2425 -919
rect 2391 -1006 2425 -987
rect 2649 -817 2683 -798
rect 2649 -885 2683 -883
rect 2649 -921 2683 -919
rect 2649 -1006 2683 -987
rect 2759 -814 2793 -798
rect 2759 -882 2793 -870
rect 2759 -950 2793 -942
rect 856 -1018 890 -1014
rect 2759 -1018 2793 -1014
rect 1017 -1083 1064 -1049
rect 1100 -1083 1134 -1049
rect 1170 -1083 1217 -1049
rect 1469 -1083 1516 -1049
rect 1552 -1083 1586 -1049
rect 1622 -1083 1669 -1049
rect 1727 -1083 1774 -1049
rect 1810 -1083 1844 -1049
rect 1880 -1083 1927 -1049
rect 1985 -1083 2032 -1049
rect 2068 -1083 2102 -1049
rect 2138 -1083 2185 -1049
rect 2437 -1083 2484 -1049
rect 2520 -1083 2554 -1049
rect 2590 -1083 2637 -1049
rect 856 -1124 890 -1120
rect 2759 -1124 2793 -1120
rect 856 -1196 890 -1188
rect 1017 -1219 1064 -1185
rect 1100 -1219 1134 -1185
rect 1170 -1219 1217 -1185
rect 1469 -1219 1516 -1185
rect 1552 -1219 1586 -1185
rect 1622 -1219 1669 -1185
rect 1727 -1219 1774 -1185
rect 1810 -1219 1844 -1185
rect 1880 -1219 1927 -1185
rect 1985 -1219 2032 -1185
rect 2068 -1219 2102 -1185
rect 2138 -1219 2185 -1185
rect 2437 -1219 2484 -1185
rect 2520 -1219 2554 -1185
rect 2590 -1219 2637 -1185
rect 2759 -1196 2793 -1188
rect 856 -1268 890 -1256
rect 856 -1340 890 -1324
rect 856 -1412 890 -1392
rect 856 -1484 890 -1460
rect 971 -1281 1005 -1262
rect 971 -1349 1005 -1347
rect 971 -1385 1005 -1383
rect 971 -1470 1005 -1451
rect 1229 -1281 1263 -1262
rect 1229 -1349 1263 -1347
rect 1229 -1385 1263 -1383
rect 1229 -1470 1263 -1451
rect 1423 -1281 1457 -1262
rect 1423 -1349 1457 -1347
rect 1423 -1385 1457 -1383
rect 1423 -1470 1457 -1451
rect 1681 -1281 1715 -1262
rect 1681 -1349 1715 -1347
rect 1681 -1385 1715 -1383
rect 1681 -1470 1715 -1451
rect 1939 -1281 1973 -1262
rect 1939 -1349 1973 -1347
rect 1939 -1385 1973 -1383
rect 1939 -1470 1973 -1451
rect 2197 -1281 2231 -1262
rect 2197 -1349 2231 -1347
rect 2197 -1385 2231 -1383
rect 2197 -1470 2231 -1451
rect 2391 -1281 2425 -1262
rect 2391 -1349 2425 -1347
rect 2391 -1385 2425 -1383
rect 2391 -1470 2425 -1451
rect 2649 -1281 2683 -1262
rect 2649 -1349 2683 -1347
rect 2649 -1385 2683 -1383
rect 2649 -1470 2683 -1451
rect 2759 -1268 2793 -1256
rect 2759 -1340 2793 -1324
rect 2759 -1412 2793 -1392
rect 856 -1556 890 -1528
rect 2759 -1484 2793 -1460
rect 2759 -1556 2793 -1528
rect 856 -1628 890 -1596
rect 856 -1698 890 -1664
rect 856 -1766 890 -1734
rect 971 -1584 1005 -1565
rect 971 -1652 1005 -1650
rect 971 -1688 1005 -1686
rect 971 -1773 1005 -1754
rect 1229 -1584 1263 -1565
rect 1229 -1652 1263 -1650
rect 1229 -1688 1263 -1686
rect 1229 -1773 1263 -1754
rect 1423 -1584 1457 -1565
rect 1423 -1652 1457 -1650
rect 1423 -1688 1457 -1686
rect 1423 -1773 1457 -1754
rect 1681 -1584 1715 -1565
rect 1681 -1652 1715 -1650
rect 1681 -1688 1715 -1686
rect 1681 -1773 1715 -1754
rect 1939 -1584 1973 -1565
rect 1939 -1652 1973 -1650
rect 1939 -1688 1973 -1686
rect 1939 -1773 1973 -1754
rect 2197 -1584 2231 -1565
rect 2197 -1652 2231 -1650
rect 2197 -1688 2231 -1686
rect 2197 -1773 2231 -1754
rect 2391 -1584 2425 -1565
rect 2391 -1652 2425 -1650
rect 2391 -1688 2425 -1686
rect 2391 -1773 2425 -1754
rect 2649 -1584 2683 -1565
rect 2649 -1652 2683 -1650
rect 2649 -1688 2683 -1686
rect 2649 -1773 2683 -1754
rect 2759 -1628 2793 -1596
rect 2759 -1698 2793 -1664
rect 2759 -1766 2793 -1734
rect 856 -1834 890 -1806
rect 1017 -1850 1064 -1816
rect 1100 -1850 1134 -1816
rect 1170 -1850 1217 -1816
rect 1469 -1850 1516 -1816
rect 1552 -1850 1586 -1816
rect 1622 -1850 1669 -1816
rect 1727 -1850 1774 -1816
rect 1810 -1850 1844 -1816
rect 1880 -1850 1927 -1816
rect 1985 -1850 2032 -1816
rect 2068 -1850 2102 -1816
rect 2138 -1850 2185 -1816
rect 2437 -1850 2484 -1816
rect 2520 -1850 2554 -1816
rect 2590 -1850 2637 -1816
rect 2759 -1834 2793 -1806
rect 856 -1902 890 -1878
rect 856 -1970 890 -1950
rect 2759 -1902 2793 -1878
rect 1017 -1992 1064 -1958
rect 1100 -1992 1134 -1958
rect 1170 -1992 1217 -1958
rect 1469 -1992 1516 -1958
rect 1552 -1992 1586 -1958
rect 1622 -1992 1669 -1958
rect 1727 -1992 1774 -1958
rect 1810 -1992 1844 -1958
rect 1880 -1992 1927 -1958
rect 1985 -1992 2032 -1958
rect 2068 -1992 2102 -1958
rect 2138 -1992 2185 -1958
rect 2437 -1992 2484 -1958
rect 2520 -1992 2554 -1958
rect 2590 -1992 2637 -1958
rect 2759 -1970 2793 -1950
rect 856 -2038 890 -2022
rect 856 -2106 890 -2094
rect 856 -2174 890 -2166
rect 856 -2310 890 -2208
rect 971 -2054 1005 -2035
rect 971 -2122 1005 -2120
rect 971 -2158 1005 -2156
rect 971 -2243 1005 -2224
rect 1229 -2054 1263 -2035
rect 1229 -2122 1263 -2120
rect 1229 -2158 1263 -2156
rect 1229 -2243 1263 -2224
rect 1423 -2054 1457 -2035
rect 1423 -2122 1457 -2120
rect 1423 -2158 1457 -2156
rect 1423 -2243 1457 -2224
rect 1681 -2054 1715 -2035
rect 1681 -2122 1715 -2120
rect 1681 -2158 1715 -2156
rect 1681 -2243 1715 -2224
rect 1939 -2054 1973 -2035
rect 1939 -2122 1973 -2120
rect 1939 -2158 1973 -2156
rect 1939 -2243 1973 -2224
rect 2197 -2054 2231 -2035
rect 2197 -2122 2231 -2120
rect 2197 -2158 2231 -2156
rect 2197 -2243 2231 -2224
rect 2391 -2054 2425 -2035
rect 2391 -2122 2425 -2120
rect 2391 -2158 2425 -2156
rect 2391 -2243 2425 -2224
rect 2649 -2054 2683 -2035
rect 2649 -2122 2683 -2120
rect 2649 -2158 2683 -2156
rect 2649 -2243 2683 -2224
rect 2759 -2038 2793 -2022
rect 2759 -2106 2793 -2094
rect 2759 -2174 2793 -2166
rect 2759 -2310 2793 -2208
rect 856 -2344 977 -2310
rect 1036 -2344 1045 -2310
rect 1108 -2344 1113 -2310
rect 1180 -2344 1181 -2310
rect 1215 -2344 1218 -2310
rect 1283 -2344 1290 -2310
rect 1351 -2344 1362 -2310
rect 1419 -2344 1434 -2310
rect 1487 -2344 1506 -2310
rect 1555 -2344 1578 -2310
rect 1623 -2344 1650 -2310
rect 1691 -2344 1722 -2310
rect 1759 -2344 1793 -2310
rect 1828 -2344 1861 -2310
rect 1900 -2344 1929 -2310
rect 1972 -2344 1997 -2310
rect 2044 -2344 2065 -2310
rect 2116 -2344 2133 -2310
rect 2188 -2344 2201 -2310
rect 2260 -2344 2269 -2310
rect 2332 -2344 2337 -2310
rect 2404 -2344 2405 -2310
rect 2439 -2344 2442 -2310
rect 2507 -2344 2514 -2310
rect 2575 -2344 2586 -2310
rect 2643 -2344 2793 -2310
<< viali >>
rect 1002 429 1011 463
rect 1011 429 1036 463
rect 1074 429 1079 463
rect 1079 429 1108 463
rect 1146 429 1147 463
rect 1147 429 1180 463
rect 1218 429 1249 463
rect 1249 429 1252 463
rect 1290 429 1317 463
rect 1317 429 1324 463
rect 1362 429 1385 463
rect 1385 429 1396 463
rect 1434 429 1453 463
rect 1453 429 1468 463
rect 1506 429 1521 463
rect 1521 429 1540 463
rect 1578 429 1589 463
rect 1589 429 1612 463
rect 1650 429 1657 463
rect 1657 429 1684 463
rect 1722 429 1725 463
rect 1725 429 1756 463
rect 1794 429 1827 463
rect 1827 429 1828 463
rect 1866 429 1895 463
rect 1895 429 1900 463
rect 1938 429 1963 463
rect 1963 429 1972 463
rect 2010 429 2031 463
rect 2031 429 2044 463
rect 2082 429 2099 463
rect 2099 429 2116 463
rect 2154 429 2167 463
rect 2167 429 2188 463
rect 2226 429 2235 463
rect 2235 429 2260 463
rect 2298 429 2303 463
rect 2303 429 2332 463
rect 2370 429 2371 463
rect 2371 429 2404 463
rect 2442 429 2473 463
rect 2473 429 2476 463
rect 2514 429 2541 463
rect 2541 429 2548 463
rect 2586 429 2609 463
rect 2609 429 2620 463
rect 856 308 890 316
rect 1064 315 1066 349
rect 1066 315 1098 349
rect 1136 315 1168 349
rect 1168 315 1170 349
rect 1516 315 1518 349
rect 1518 315 1550 349
rect 1588 315 1620 349
rect 1620 315 1622 349
rect 1774 315 1776 349
rect 1776 315 1808 349
rect 1846 315 1878 349
rect 1878 315 1880 349
rect 2032 315 2034 349
rect 2034 315 2066 349
rect 2104 315 2136 349
rect 2136 315 2138 349
rect 2484 315 2486 349
rect 2486 315 2518 349
rect 2556 315 2588 349
rect 2588 315 2590 349
rect 856 282 890 308
rect 2759 308 2793 316
rect 2759 282 2793 308
rect 856 240 890 244
rect 856 210 890 240
rect 856 138 890 172
rect 856 70 890 100
rect 856 66 890 70
rect 971 219 1005 221
rect 971 187 1005 219
rect 971 117 1005 149
rect 971 115 1005 117
rect 1229 219 1263 221
rect 1229 187 1263 219
rect 1229 117 1263 149
rect 1229 115 1263 117
rect 1423 219 1457 221
rect 1423 187 1457 219
rect 1423 117 1457 149
rect 1423 115 1457 117
rect 1681 219 1715 221
rect 1681 187 1715 219
rect 1681 117 1715 149
rect 1681 115 1715 117
rect 1939 219 1973 221
rect 1939 187 1973 219
rect 1939 117 1973 149
rect 1939 115 1973 117
rect 2197 219 2231 221
rect 2197 187 2231 219
rect 2197 117 2231 149
rect 2197 115 2231 117
rect 2391 219 2425 221
rect 2391 187 2425 219
rect 2391 117 2425 149
rect 2391 115 2425 117
rect 2649 219 2683 221
rect 2649 187 2683 219
rect 2649 117 2683 149
rect 2649 115 2683 117
rect 2759 240 2793 244
rect 2759 210 2793 240
rect 2759 138 2793 172
rect 2759 70 2793 100
rect 2759 66 2793 70
rect 856 2 890 28
rect 856 -6 890 2
rect 2759 2 2793 28
rect 2759 -6 2793 2
rect 856 -66 890 -44
rect 856 -78 890 -66
rect 856 -134 890 -116
rect 856 -150 890 -134
rect 856 -202 890 -188
rect 856 -222 890 -202
rect 971 -84 1005 -82
rect 971 -116 1005 -84
rect 971 -186 1005 -154
rect 971 -188 1005 -186
rect 1229 -84 1263 -82
rect 1229 -116 1263 -84
rect 1229 -186 1263 -154
rect 1229 -188 1263 -186
rect 1423 -84 1457 -82
rect 1423 -116 1457 -84
rect 1423 -186 1457 -154
rect 1423 -188 1457 -186
rect 1681 -84 1715 -82
rect 1681 -116 1715 -84
rect 1681 -186 1715 -154
rect 1681 -188 1715 -186
rect 1939 -84 1973 -82
rect 1939 -116 1973 -84
rect 1939 -186 1973 -154
rect 1939 -188 1973 -186
rect 2197 -84 2231 -82
rect 2197 -116 2231 -84
rect 2197 -186 2231 -154
rect 2197 -188 2231 -186
rect 2391 -84 2425 -82
rect 2391 -116 2425 -84
rect 2391 -186 2425 -154
rect 2391 -188 2425 -186
rect 2649 -84 2683 -82
rect 2649 -116 2683 -84
rect 2649 -186 2683 -154
rect 2649 -188 2683 -186
rect 2759 -66 2793 -44
rect 2759 -78 2793 -66
rect 2759 -134 2793 -116
rect 2759 -150 2793 -134
rect 2759 -202 2793 -188
rect 2759 -222 2793 -202
rect 856 -270 890 -260
rect 856 -294 890 -270
rect 2759 -270 2793 -260
rect 1064 -316 1066 -282
rect 1066 -316 1098 -282
rect 1136 -316 1168 -282
rect 1168 -316 1170 -282
rect 1516 -316 1518 -282
rect 1518 -316 1550 -282
rect 1588 -316 1620 -282
rect 1620 -316 1622 -282
rect 1774 -316 1776 -282
rect 1776 -316 1808 -282
rect 1846 -316 1878 -282
rect 1878 -316 1880 -282
rect 2032 -316 2034 -282
rect 2034 -316 2066 -282
rect 2104 -316 2136 -282
rect 2136 -316 2138 -282
rect 2484 -316 2486 -282
rect 2486 -316 2518 -282
rect 2556 -316 2588 -282
rect 2588 -316 2590 -282
rect 2759 -294 2793 -270
rect 856 -338 890 -332
rect 856 -366 890 -338
rect 856 -406 890 -404
rect 856 -438 890 -406
rect 2759 -338 2793 -332
rect 2759 -366 2793 -338
rect 2759 -406 2793 -404
rect 1064 -452 1066 -418
rect 1066 -452 1098 -418
rect 1136 -452 1168 -418
rect 1168 -452 1170 -418
rect 1516 -452 1518 -418
rect 1518 -452 1550 -418
rect 1588 -452 1620 -418
rect 1620 -452 1622 -418
rect 1774 -452 1776 -418
rect 1776 -452 1808 -418
rect 1846 -452 1878 -418
rect 1878 -452 1880 -418
rect 2032 -452 2034 -418
rect 2034 -452 2066 -418
rect 2104 -452 2136 -418
rect 2136 -452 2138 -418
rect 2484 -452 2486 -418
rect 2486 -452 2518 -418
rect 2556 -452 2588 -418
rect 2588 -452 2590 -418
rect 2759 -438 2793 -406
rect 856 -508 890 -476
rect 856 -510 890 -508
rect 856 -576 890 -548
rect 856 -582 890 -576
rect 856 -644 890 -620
rect 856 -654 890 -644
rect 856 -712 890 -692
rect 971 -548 1005 -546
rect 971 -580 1005 -548
rect 971 -650 1005 -618
rect 971 -652 1005 -650
rect 1229 -548 1263 -546
rect 1229 -580 1263 -548
rect 1229 -650 1263 -618
rect 1229 -652 1263 -650
rect 1423 -548 1457 -546
rect 1423 -580 1457 -548
rect 1423 -650 1457 -618
rect 1423 -652 1457 -650
rect 1681 -548 1715 -546
rect 1681 -580 1715 -548
rect 1681 -650 1715 -618
rect 1681 -652 1715 -650
rect 1939 -548 1973 -546
rect 1939 -580 1973 -548
rect 1939 -650 1973 -618
rect 1939 -652 1973 -650
rect 2197 -548 2231 -546
rect 2197 -580 2231 -548
rect 2197 -650 2231 -618
rect 2197 -652 2231 -650
rect 2391 -548 2425 -546
rect 2391 -580 2425 -548
rect 2391 -650 2425 -618
rect 2391 -652 2425 -650
rect 2649 -548 2683 -546
rect 2649 -580 2683 -548
rect 2649 -650 2683 -618
rect 2649 -652 2683 -650
rect 2759 -508 2793 -476
rect 2759 -510 2793 -508
rect 2759 -576 2793 -548
rect 2759 -582 2793 -576
rect 2759 -644 2793 -620
rect 2759 -654 2793 -644
rect 856 -726 890 -712
rect 856 -780 890 -764
rect 856 -798 890 -780
rect 2759 -712 2793 -692
rect 2759 -726 2793 -712
rect 2759 -780 2793 -764
rect 2759 -798 2793 -780
rect 856 -848 890 -836
rect 856 -870 890 -848
rect 856 -916 890 -908
rect 856 -942 890 -916
rect 856 -984 890 -980
rect 856 -1014 890 -984
rect 971 -851 1005 -849
rect 971 -883 1005 -851
rect 971 -953 1005 -921
rect 971 -955 1005 -953
rect 1229 -851 1263 -849
rect 1229 -883 1263 -851
rect 1229 -953 1263 -921
rect 1229 -955 1263 -953
rect 1423 -851 1457 -849
rect 1423 -883 1457 -851
rect 1423 -953 1457 -921
rect 1423 -955 1457 -953
rect 1681 -851 1715 -849
rect 1681 -883 1715 -851
rect 1681 -953 1715 -921
rect 1681 -955 1715 -953
rect 1939 -851 1973 -849
rect 1939 -883 1973 -851
rect 1939 -953 1973 -921
rect 1939 -955 1973 -953
rect 2197 -851 2231 -849
rect 2197 -883 2231 -851
rect 2197 -953 2231 -921
rect 2197 -955 2231 -953
rect 2391 -851 2425 -849
rect 2391 -883 2425 -851
rect 2391 -953 2425 -921
rect 2391 -955 2425 -953
rect 2649 -851 2683 -849
rect 2649 -883 2683 -851
rect 2649 -953 2683 -921
rect 2649 -955 2683 -953
rect 2759 -848 2793 -836
rect 2759 -870 2793 -848
rect 2759 -916 2793 -908
rect 2759 -942 2793 -916
rect 2759 -984 2793 -980
rect 2759 -1014 2793 -984
rect 856 -1086 890 -1052
rect 1064 -1083 1066 -1049
rect 1066 -1083 1098 -1049
rect 1136 -1083 1168 -1049
rect 1168 -1083 1170 -1049
rect 1516 -1083 1518 -1049
rect 1518 -1083 1550 -1049
rect 1588 -1083 1620 -1049
rect 1620 -1083 1622 -1049
rect 1774 -1083 1776 -1049
rect 1776 -1083 1808 -1049
rect 1846 -1083 1878 -1049
rect 1878 -1083 1880 -1049
rect 2032 -1083 2034 -1049
rect 2034 -1083 2066 -1049
rect 2104 -1083 2136 -1049
rect 2136 -1083 2138 -1049
rect 2484 -1083 2486 -1049
rect 2486 -1083 2518 -1049
rect 2556 -1083 2588 -1049
rect 2588 -1083 2590 -1049
rect 856 -1154 890 -1124
rect 856 -1158 890 -1154
rect 2759 -1086 2793 -1052
rect 2759 -1154 2793 -1124
rect 2759 -1158 2793 -1154
rect 856 -1222 890 -1196
rect 1064 -1219 1066 -1185
rect 1066 -1219 1098 -1185
rect 1136 -1219 1168 -1185
rect 1168 -1219 1170 -1185
rect 1516 -1219 1518 -1185
rect 1518 -1219 1550 -1185
rect 1588 -1219 1620 -1185
rect 1620 -1219 1622 -1185
rect 1774 -1219 1776 -1185
rect 1776 -1219 1808 -1185
rect 1846 -1219 1878 -1185
rect 1878 -1219 1880 -1185
rect 2032 -1219 2034 -1185
rect 2034 -1219 2066 -1185
rect 2104 -1219 2136 -1185
rect 2136 -1219 2138 -1185
rect 2484 -1219 2486 -1185
rect 2486 -1219 2518 -1185
rect 2556 -1219 2588 -1185
rect 2588 -1219 2590 -1185
rect 856 -1230 890 -1222
rect 2759 -1222 2793 -1196
rect 2759 -1230 2793 -1222
rect 856 -1290 890 -1268
rect 856 -1302 890 -1290
rect 856 -1358 890 -1340
rect 856 -1374 890 -1358
rect 856 -1426 890 -1412
rect 856 -1446 890 -1426
rect 971 -1315 1005 -1313
rect 971 -1347 1005 -1315
rect 971 -1417 1005 -1385
rect 971 -1419 1005 -1417
rect 1229 -1315 1263 -1313
rect 1229 -1347 1263 -1315
rect 1229 -1417 1263 -1385
rect 1229 -1419 1263 -1417
rect 1423 -1315 1457 -1313
rect 1423 -1347 1457 -1315
rect 1423 -1417 1457 -1385
rect 1423 -1419 1457 -1417
rect 1681 -1315 1715 -1313
rect 1681 -1347 1715 -1315
rect 1681 -1417 1715 -1385
rect 1681 -1419 1715 -1417
rect 1939 -1315 1973 -1313
rect 1939 -1347 1973 -1315
rect 1939 -1417 1973 -1385
rect 1939 -1419 1973 -1417
rect 2197 -1315 2231 -1313
rect 2197 -1347 2231 -1315
rect 2197 -1417 2231 -1385
rect 2197 -1419 2231 -1417
rect 2391 -1315 2425 -1313
rect 2391 -1347 2425 -1315
rect 2391 -1417 2425 -1385
rect 2391 -1419 2425 -1417
rect 2649 -1315 2683 -1313
rect 2649 -1347 2683 -1315
rect 2649 -1417 2683 -1385
rect 2649 -1419 2683 -1417
rect 2759 -1290 2793 -1268
rect 2759 -1302 2793 -1290
rect 2759 -1358 2793 -1340
rect 2759 -1374 2793 -1358
rect 2759 -1426 2793 -1412
rect 2759 -1446 2793 -1426
rect 856 -1494 890 -1484
rect 856 -1518 890 -1494
rect 856 -1562 890 -1556
rect 856 -1590 890 -1562
rect 2759 -1494 2793 -1484
rect 2759 -1518 2793 -1494
rect 2759 -1562 2793 -1556
rect 856 -1630 890 -1628
rect 856 -1662 890 -1630
rect 856 -1732 890 -1700
rect 856 -1734 890 -1732
rect 856 -1800 890 -1772
rect 971 -1618 1005 -1616
rect 971 -1650 1005 -1618
rect 971 -1720 1005 -1688
rect 971 -1722 1005 -1720
rect 1229 -1618 1263 -1616
rect 1229 -1650 1263 -1618
rect 1229 -1720 1263 -1688
rect 1229 -1722 1263 -1720
rect 1423 -1618 1457 -1616
rect 1423 -1650 1457 -1618
rect 1423 -1720 1457 -1688
rect 1423 -1722 1457 -1720
rect 1681 -1618 1715 -1616
rect 1681 -1650 1715 -1618
rect 1681 -1720 1715 -1688
rect 1681 -1722 1715 -1720
rect 1939 -1618 1973 -1616
rect 1939 -1650 1973 -1618
rect 1939 -1720 1973 -1688
rect 1939 -1722 1973 -1720
rect 2197 -1618 2231 -1616
rect 2197 -1650 2231 -1618
rect 2197 -1720 2231 -1688
rect 2197 -1722 2231 -1720
rect 2391 -1618 2425 -1616
rect 2391 -1650 2425 -1618
rect 2391 -1720 2425 -1688
rect 2391 -1722 2425 -1720
rect 2649 -1618 2683 -1616
rect 2649 -1650 2683 -1618
rect 2649 -1720 2683 -1688
rect 2649 -1722 2683 -1720
rect 2759 -1590 2793 -1562
rect 2759 -1630 2793 -1628
rect 2759 -1662 2793 -1630
rect 2759 -1732 2793 -1700
rect 2759 -1734 2793 -1732
rect 856 -1806 890 -1800
rect 2759 -1800 2793 -1772
rect 2759 -1806 2793 -1800
rect 856 -1868 890 -1844
rect 1064 -1850 1066 -1816
rect 1066 -1850 1098 -1816
rect 1136 -1850 1168 -1816
rect 1168 -1850 1170 -1816
rect 1516 -1850 1518 -1816
rect 1518 -1850 1550 -1816
rect 1588 -1850 1620 -1816
rect 1620 -1850 1622 -1816
rect 1774 -1850 1776 -1816
rect 1776 -1850 1808 -1816
rect 1846 -1850 1878 -1816
rect 1878 -1850 1880 -1816
rect 2032 -1850 2034 -1816
rect 2034 -1850 2066 -1816
rect 2104 -1850 2136 -1816
rect 2136 -1850 2138 -1816
rect 2484 -1850 2486 -1816
rect 2486 -1850 2518 -1816
rect 2556 -1850 2588 -1816
rect 2588 -1850 2590 -1816
rect 856 -1878 890 -1868
rect 856 -1936 890 -1916
rect 856 -1950 890 -1936
rect 2759 -1868 2793 -1844
rect 2759 -1878 2793 -1868
rect 2759 -1936 2793 -1916
rect 2759 -1950 2793 -1936
rect 856 -2004 890 -1988
rect 1064 -1992 1066 -1958
rect 1066 -1992 1098 -1958
rect 1136 -1992 1168 -1958
rect 1168 -1992 1170 -1958
rect 1516 -1992 1518 -1958
rect 1518 -1992 1550 -1958
rect 1588 -1992 1620 -1958
rect 1620 -1992 1622 -1958
rect 1774 -1992 1776 -1958
rect 1776 -1992 1808 -1958
rect 1846 -1992 1878 -1958
rect 1878 -1992 1880 -1958
rect 2032 -1992 2034 -1958
rect 2034 -1992 2066 -1958
rect 2104 -1992 2136 -1958
rect 2136 -1992 2138 -1958
rect 2484 -1992 2486 -1958
rect 2486 -1992 2518 -1958
rect 2556 -1992 2588 -1958
rect 2588 -1992 2590 -1958
rect 856 -2022 890 -2004
rect 2759 -2004 2793 -1988
rect 2759 -2022 2793 -2004
rect 856 -2072 890 -2060
rect 856 -2094 890 -2072
rect 856 -2140 890 -2132
rect 856 -2166 890 -2140
rect 971 -2088 1005 -2086
rect 971 -2120 1005 -2088
rect 971 -2190 1005 -2158
rect 971 -2192 1005 -2190
rect 1229 -2088 1263 -2086
rect 1229 -2120 1263 -2088
rect 1229 -2190 1263 -2158
rect 1229 -2192 1263 -2190
rect 1423 -2088 1457 -2086
rect 1423 -2120 1457 -2088
rect 1423 -2190 1457 -2158
rect 1423 -2192 1457 -2190
rect 1681 -2088 1715 -2086
rect 1681 -2120 1715 -2088
rect 1681 -2190 1715 -2158
rect 1681 -2192 1715 -2190
rect 1939 -2088 1973 -2086
rect 1939 -2120 1973 -2088
rect 1939 -2190 1973 -2158
rect 1939 -2192 1973 -2190
rect 2197 -2088 2231 -2086
rect 2197 -2120 2231 -2088
rect 2197 -2190 2231 -2158
rect 2197 -2192 2231 -2190
rect 2391 -2088 2425 -2086
rect 2391 -2120 2425 -2088
rect 2391 -2190 2425 -2158
rect 2391 -2192 2425 -2190
rect 2649 -2088 2683 -2086
rect 2649 -2120 2683 -2088
rect 2649 -2190 2683 -2158
rect 2649 -2192 2683 -2190
rect 2759 -2072 2793 -2060
rect 2759 -2094 2793 -2072
rect 2759 -2140 2793 -2132
rect 2759 -2166 2793 -2140
rect 1002 -2344 1011 -2310
rect 1011 -2344 1036 -2310
rect 1074 -2344 1079 -2310
rect 1079 -2344 1108 -2310
rect 1146 -2344 1147 -2310
rect 1147 -2344 1180 -2310
rect 1218 -2344 1249 -2310
rect 1249 -2344 1252 -2310
rect 1290 -2344 1317 -2310
rect 1317 -2344 1324 -2310
rect 1362 -2344 1385 -2310
rect 1385 -2344 1396 -2310
rect 1434 -2344 1453 -2310
rect 1453 -2344 1468 -2310
rect 1506 -2344 1521 -2310
rect 1521 -2344 1540 -2310
rect 1578 -2344 1589 -2310
rect 1589 -2344 1612 -2310
rect 1650 -2344 1657 -2310
rect 1657 -2344 1684 -2310
rect 1722 -2344 1725 -2310
rect 1725 -2344 1756 -2310
rect 1794 -2344 1827 -2310
rect 1827 -2344 1828 -2310
rect 1866 -2344 1895 -2310
rect 1895 -2344 1900 -2310
rect 1938 -2344 1963 -2310
rect 1963 -2344 1972 -2310
rect 2010 -2344 2031 -2310
rect 2031 -2344 2044 -2310
rect 2082 -2344 2099 -2310
rect 2099 -2344 2116 -2310
rect 2154 -2344 2167 -2310
rect 2167 -2344 2188 -2310
rect 2226 -2344 2235 -2310
rect 2235 -2344 2260 -2310
rect 2298 -2344 2303 -2310
rect 2303 -2344 2332 -2310
rect 2370 -2344 2371 -2310
rect 2371 -2344 2404 -2310
rect 2442 -2344 2473 -2310
rect 2473 -2344 2476 -2310
rect 2514 -2344 2541 -2310
rect 2541 -2344 2548 -2310
rect 2586 -2344 2609 -2310
rect 2609 -2344 2620 -2310
<< metal1 >>
rect 831 463 2804 488
rect 831 429 1002 463
rect 1036 429 1074 463
rect 1108 429 1146 463
rect 1180 429 1218 463
rect 1252 429 1290 463
rect 1324 429 1362 463
rect 1396 429 1434 463
rect 1468 429 1506 463
rect 1540 429 1578 463
rect 1612 429 1650 463
rect 1684 429 1722 463
rect 1756 429 1794 463
rect 1828 429 1866 463
rect 1900 429 1938 463
rect 1972 429 2010 463
rect 2044 429 2082 463
rect 2116 429 2154 463
rect 2188 429 2226 463
rect 2260 429 2298 463
rect 2332 429 2370 463
rect 2404 429 2442 463
rect 2476 429 2514 463
rect 2548 429 2586 463
rect 2620 429 2804 463
rect 831 349 2804 429
rect 831 316 1064 349
rect 831 282 856 316
rect 890 315 1064 316
rect 1098 315 1136 349
rect 1170 315 1516 349
rect 1550 315 1588 349
rect 1622 315 1774 349
rect 1808 315 1846 349
rect 1880 315 2032 349
rect 2066 315 2104 349
rect 2138 315 2484 349
rect 2518 315 2556 349
rect 2590 316 2804 349
rect 2590 315 2759 316
rect 890 282 2759 315
rect 2793 282 2804 316
rect 831 244 2804 282
rect 831 210 856 244
rect 890 221 2759 244
rect 890 210 971 221
rect 831 187 971 210
rect 1005 187 1229 221
rect 1263 187 1423 221
rect 1457 187 1681 221
rect 1715 187 1939 221
rect 1973 187 2197 221
rect 2231 187 2391 221
rect 2425 187 2649 221
rect 2683 210 2759 221
rect 2793 210 2804 244
rect 2683 187 2804 210
rect 831 172 2804 187
rect 831 138 856 172
rect 890 149 2759 172
rect 890 138 971 149
rect 831 115 971 138
rect 1005 115 1229 149
rect 1263 115 1423 149
rect 1457 115 1681 149
rect 1715 115 1939 149
rect 1973 115 2197 149
rect 2231 115 2391 149
rect 2425 115 2649 149
rect 2683 138 2759 149
rect 2793 138 2804 172
rect 2683 115 2804 138
rect 831 100 2804 115
rect 831 66 856 100
rect 890 68 2759 100
rect 890 66 1269 68
rect 831 28 1269 66
rect 831 -6 856 28
rect 890 -6 1269 28
rect 831 -35 1269 -6
rect 2385 66 2759 68
rect 2793 66 2804 100
rect 2385 28 2804 66
rect 2385 -6 2759 28
rect 2793 -6 2804 28
rect 831 -44 1463 -35
rect 831 -78 856 -44
rect 890 -78 1463 -44
rect 831 -82 1463 -78
rect 831 -116 971 -82
rect 1005 -116 1229 -82
rect 1263 -116 1423 -82
rect 1457 -116 1463 -82
rect 831 -150 856 -116
rect 890 -150 1463 -116
rect 831 -154 1463 -150
rect 831 -188 971 -154
rect 1005 -188 1229 -154
rect 1263 -188 1423 -154
rect 1457 -188 1463 -154
rect 831 -222 856 -188
rect 890 -222 1463 -188
rect 831 -235 1463 -222
rect 1675 -82 1721 -35
rect 1675 -116 1681 -82
rect 1715 -116 1721 -82
rect 1675 -154 1721 -116
rect 1675 -188 1681 -154
rect 1715 -188 1721 -154
rect 1675 -235 1721 -188
rect 1933 -82 1979 -35
rect 1933 -116 1939 -82
rect 1973 -116 1979 -82
rect 1933 -154 1979 -116
rect 1933 -188 1939 -154
rect 1973 -188 1979 -154
rect 1933 -235 1979 -188
rect 2191 -82 2311 -35
rect 2191 -116 2197 -82
rect 2231 -116 2311 -82
rect 2191 -154 2311 -116
rect 2191 -188 2197 -154
rect 2231 -188 2311 -154
rect 831 -260 1386 -235
rect 831 -294 856 -260
rect 890 -282 1386 -260
rect 2191 -276 2311 -188
rect 890 -294 1064 -282
rect 831 -316 1064 -294
rect 1098 -316 1136 -282
rect 1170 -316 1386 -282
rect 831 -332 1386 -316
rect 831 -366 856 -332
rect 890 -366 1386 -332
rect 831 -404 1386 -366
rect 831 -438 856 -404
rect 890 -418 1386 -404
rect 890 -438 1064 -418
rect 831 -452 1064 -438
rect 1098 -452 1136 -418
rect 1170 -452 1386 -418
rect 831 -476 1386 -452
rect 1473 -282 2311 -276
rect 1473 -306 1516 -282
rect 1550 -306 1588 -282
rect 1622 -306 1774 -282
rect 1808 -306 1846 -282
rect 1880 -306 2032 -282
rect 2066 -306 2104 -282
rect 2138 -306 2311 -282
rect 1473 -358 1502 -306
rect 1554 -358 1566 -306
rect 1622 -316 1630 -306
rect 1618 -358 1630 -316
rect 1682 -358 1736 -306
rect 1788 -358 1800 -316
rect 1852 -358 1864 -316
rect 1916 -358 1976 -306
rect 2028 -316 2032 -306
rect 2028 -358 2040 -316
rect 2092 -358 2104 -306
rect 2156 -358 2311 -306
rect 1473 -376 2311 -358
rect 1473 -428 1502 -376
rect 1554 -428 1566 -376
rect 1618 -418 1630 -376
rect 1622 -428 1630 -418
rect 1682 -428 1736 -376
rect 1788 -418 1800 -376
rect 1852 -418 1864 -376
rect 1916 -428 1976 -376
rect 2028 -418 2040 -376
rect 2028 -428 2032 -418
rect 2092 -428 2104 -376
rect 2156 -428 2311 -376
rect 1473 -452 1516 -428
rect 1550 -452 1588 -428
rect 1622 -452 1774 -428
rect 1808 -452 1846 -428
rect 1880 -452 2032 -428
rect 2066 -452 2104 -428
rect 2138 -452 2311 -428
rect 1473 -458 2311 -452
rect 831 -510 856 -476
rect 890 -499 1386 -476
rect 890 -510 1463 -499
rect 831 -546 1463 -510
rect 831 -548 971 -546
rect 831 -582 856 -548
rect 890 -580 971 -548
rect 1005 -580 1229 -546
rect 1263 -580 1423 -546
rect 1457 -580 1463 -546
rect 890 -582 1463 -580
rect 831 -618 1463 -582
rect 831 -620 971 -618
rect 831 -654 856 -620
rect 890 -652 971 -620
rect 1005 -652 1229 -618
rect 1263 -652 1423 -618
rect 1457 -652 1463 -618
rect 890 -654 1463 -652
rect 831 -692 1463 -654
rect 831 -726 856 -692
rect 890 -699 1463 -692
rect 1675 -546 1721 -499
rect 1675 -580 1681 -546
rect 1715 -580 1721 -546
rect 1675 -618 1721 -580
rect 1675 -652 1681 -618
rect 1715 -652 1721 -618
rect 1675 -699 1721 -652
rect 1933 -546 1979 -499
rect 1933 -580 1939 -546
rect 1973 -580 1979 -546
rect 1933 -618 1979 -580
rect 1933 -652 1939 -618
rect 1973 -652 1979 -618
rect 1933 -699 1979 -652
rect 2191 -546 2311 -458
rect 2191 -580 2197 -546
rect 2231 -580 2311 -546
rect 2191 -618 2311 -580
rect 2191 -652 2197 -618
rect 2231 -652 2311 -618
rect 890 -726 1386 -699
rect 831 -764 1386 -726
rect 831 -798 856 -764
rect 890 -798 1386 -764
rect 831 -802 1386 -798
rect 831 -836 1463 -802
rect 831 -870 856 -836
rect 890 -849 1463 -836
rect 890 -870 971 -849
rect 831 -883 971 -870
rect 1005 -883 1229 -849
rect 1263 -883 1423 -849
rect 1457 -883 1463 -849
rect 831 -908 1463 -883
rect 831 -942 856 -908
rect 890 -921 1463 -908
rect 890 -942 971 -921
rect 831 -955 971 -942
rect 1005 -955 1229 -921
rect 1263 -955 1423 -921
rect 1457 -955 1463 -921
rect 831 -980 1463 -955
rect 831 -1014 856 -980
rect 890 -1002 1463 -980
rect 1675 -849 1721 -802
rect 1675 -883 1681 -849
rect 1715 -883 1721 -849
rect 1675 -921 1721 -883
rect 1675 -955 1681 -921
rect 1715 -955 1721 -921
rect 1675 -1002 1721 -955
rect 1933 -849 1979 -802
rect 1933 -883 1939 -849
rect 1973 -883 1979 -849
rect 1933 -921 1979 -883
rect 1933 -955 1939 -921
rect 1973 -955 1979 -921
rect 1933 -1002 1979 -955
rect 2191 -849 2311 -652
rect 2191 -883 2197 -849
rect 2231 -883 2311 -849
rect 2191 -921 2311 -883
rect 2191 -955 2197 -921
rect 2231 -955 2311 -921
rect 890 -1014 1386 -1002
rect 831 -1049 1386 -1014
rect 2191 -1043 2311 -955
rect 831 -1052 1064 -1049
rect 831 -1086 856 -1052
rect 890 -1083 1064 -1052
rect 1098 -1083 1136 -1049
rect 1170 -1083 1386 -1049
rect 890 -1086 1386 -1083
rect 831 -1124 1386 -1086
rect 831 -1158 856 -1124
rect 890 -1158 1386 -1124
rect 831 -1185 1386 -1158
rect 831 -1196 1064 -1185
rect 831 -1230 856 -1196
rect 890 -1219 1064 -1196
rect 1098 -1219 1136 -1185
rect 1170 -1219 1386 -1185
rect 890 -1230 1386 -1219
rect 1473 -1049 2311 -1043
rect 1473 -1073 1516 -1049
rect 1550 -1073 1588 -1049
rect 1622 -1073 1774 -1049
rect 1808 -1073 1846 -1049
rect 1880 -1073 2032 -1049
rect 2066 -1073 2104 -1049
rect 2138 -1073 2311 -1049
rect 1473 -1125 1502 -1073
rect 1554 -1125 1566 -1073
rect 1622 -1083 1630 -1073
rect 1618 -1125 1630 -1083
rect 1682 -1125 1736 -1073
rect 1788 -1125 1800 -1083
rect 1852 -1125 1864 -1083
rect 1916 -1125 1976 -1073
rect 2028 -1083 2032 -1073
rect 2028 -1125 2040 -1083
rect 2092 -1125 2104 -1073
rect 2156 -1125 2311 -1073
rect 1473 -1143 2311 -1125
rect 1473 -1195 1502 -1143
rect 1554 -1195 1566 -1143
rect 1618 -1185 1630 -1143
rect 1622 -1195 1630 -1185
rect 1682 -1195 1736 -1143
rect 1788 -1185 1800 -1143
rect 1852 -1185 1864 -1143
rect 1916 -1195 1976 -1143
rect 2028 -1185 2040 -1143
rect 2028 -1195 2032 -1185
rect 2092 -1195 2104 -1143
rect 2156 -1195 2311 -1143
rect 1473 -1219 1516 -1195
rect 1550 -1219 1588 -1195
rect 1622 -1219 1774 -1195
rect 1808 -1219 1846 -1195
rect 1880 -1219 2032 -1195
rect 2066 -1219 2104 -1195
rect 2138 -1219 2311 -1195
rect 1473 -1225 2311 -1219
rect 831 -1266 1386 -1230
rect 831 -1268 1463 -1266
rect 831 -1302 856 -1268
rect 890 -1302 1463 -1268
rect 831 -1313 1463 -1302
rect 831 -1340 971 -1313
rect 831 -1374 856 -1340
rect 890 -1347 971 -1340
rect 1005 -1347 1229 -1313
rect 1263 -1347 1423 -1313
rect 1457 -1347 1463 -1313
rect 890 -1374 1463 -1347
rect 831 -1385 1463 -1374
rect 831 -1412 971 -1385
rect 831 -1446 856 -1412
rect 890 -1419 971 -1412
rect 1005 -1419 1229 -1385
rect 1263 -1419 1423 -1385
rect 1457 -1419 1463 -1385
rect 890 -1446 1463 -1419
rect 831 -1466 1463 -1446
rect 1675 -1313 1721 -1266
rect 1675 -1347 1681 -1313
rect 1715 -1347 1721 -1313
rect 1675 -1385 1721 -1347
rect 1675 -1419 1681 -1385
rect 1715 -1419 1721 -1385
rect 1675 -1466 1721 -1419
rect 1933 -1313 1979 -1266
rect 1933 -1347 1939 -1313
rect 1973 -1347 1979 -1313
rect 1933 -1385 1979 -1347
rect 1933 -1419 1939 -1385
rect 1973 -1419 1979 -1385
rect 1933 -1466 1979 -1419
rect 2191 -1313 2311 -1225
rect 2191 -1347 2197 -1313
rect 2231 -1347 2311 -1313
rect 2191 -1385 2311 -1347
rect 2191 -1419 2197 -1385
rect 2231 -1419 2311 -1385
rect 831 -1484 1386 -1466
rect 831 -1518 856 -1484
rect 890 -1518 1386 -1484
rect 831 -1556 1386 -1518
rect 831 -1590 856 -1556
rect 890 -1569 1386 -1556
rect 890 -1590 1463 -1569
rect 831 -1616 1463 -1590
rect 831 -1628 971 -1616
rect 831 -1662 856 -1628
rect 890 -1650 971 -1628
rect 1005 -1650 1229 -1616
rect 1263 -1650 1423 -1616
rect 1457 -1650 1463 -1616
rect 890 -1662 1463 -1650
rect 831 -1688 1463 -1662
rect 831 -1700 971 -1688
rect 831 -1734 856 -1700
rect 890 -1722 971 -1700
rect 1005 -1722 1229 -1688
rect 1263 -1722 1423 -1688
rect 1457 -1722 1463 -1688
rect 890 -1734 1463 -1722
rect 831 -1769 1463 -1734
rect 1675 -1616 1721 -1569
rect 1675 -1650 1681 -1616
rect 1715 -1650 1721 -1616
rect 1675 -1688 1721 -1650
rect 1675 -1722 1681 -1688
rect 1715 -1722 1721 -1688
rect 1675 -1769 1721 -1722
rect 1933 -1616 1979 -1569
rect 1933 -1650 1939 -1616
rect 1973 -1650 1979 -1616
rect 1933 -1688 1979 -1650
rect 1933 -1722 1939 -1688
rect 1973 -1722 1979 -1688
rect 1933 -1769 1979 -1722
rect 2191 -1616 2311 -1419
rect 2191 -1650 2197 -1616
rect 2231 -1650 2311 -1616
rect 2191 -1688 2311 -1650
rect 2191 -1722 2197 -1688
rect 2231 -1722 2311 -1688
rect 831 -1772 1269 -1769
rect 831 -1806 856 -1772
rect 890 -1806 1269 -1772
rect 831 -1816 1269 -1806
rect 2191 -1810 2311 -1722
rect 831 -1844 1064 -1816
rect 831 -1878 856 -1844
rect 890 -1850 1064 -1844
rect 1098 -1850 1136 -1816
rect 1170 -1850 1269 -1816
rect 890 -1878 1269 -1850
rect 831 -1916 1269 -1878
rect 1473 -1816 2311 -1810
rect 1473 -1818 1516 -1816
rect 1550 -1818 1588 -1816
rect 1622 -1818 1774 -1816
rect 1808 -1818 1846 -1816
rect 1880 -1818 2032 -1816
rect 2066 -1818 2104 -1816
rect 2138 -1818 2311 -1816
rect 1473 -1870 1502 -1818
rect 1554 -1870 1566 -1818
rect 1622 -1850 1630 -1818
rect 1618 -1870 1630 -1850
rect 1682 -1870 1736 -1818
rect 1788 -1870 1800 -1850
rect 1852 -1870 1864 -1850
rect 1916 -1870 1976 -1818
rect 2028 -1850 2032 -1818
rect 2028 -1870 2040 -1850
rect 2092 -1870 2104 -1818
rect 2156 -1870 2311 -1818
rect 1473 -1880 2311 -1870
rect 2385 -44 2804 -6
rect 2385 -78 2759 -44
rect 2793 -78 2804 -44
rect 2385 -82 2804 -78
rect 2385 -116 2391 -82
rect 2425 -116 2649 -82
rect 2683 -116 2804 -82
rect 2385 -150 2759 -116
rect 2793 -150 2804 -116
rect 2385 -154 2804 -150
rect 2385 -188 2391 -154
rect 2425 -188 2649 -154
rect 2683 -188 2804 -154
rect 2385 -222 2759 -188
rect 2793 -222 2804 -188
rect 2385 -260 2804 -222
rect 2385 -282 2759 -260
rect 2385 -316 2484 -282
rect 2518 -316 2556 -282
rect 2590 -294 2759 -282
rect 2793 -294 2804 -260
rect 2590 -316 2804 -294
rect 2385 -332 2804 -316
rect 2385 -366 2759 -332
rect 2793 -366 2804 -332
rect 2385 -404 2804 -366
rect 2385 -418 2759 -404
rect 2385 -452 2484 -418
rect 2518 -452 2556 -418
rect 2590 -438 2759 -418
rect 2793 -438 2804 -404
rect 2590 -452 2804 -438
rect 2385 -476 2804 -452
rect 2385 -510 2759 -476
rect 2793 -510 2804 -476
rect 2385 -546 2804 -510
rect 2385 -580 2391 -546
rect 2425 -580 2649 -546
rect 2683 -548 2804 -546
rect 2683 -580 2759 -548
rect 2385 -582 2759 -580
rect 2793 -582 2804 -548
rect 2385 -618 2804 -582
rect 2385 -652 2391 -618
rect 2425 -652 2649 -618
rect 2683 -620 2804 -618
rect 2683 -652 2759 -620
rect 2385 -654 2759 -652
rect 2793 -654 2804 -620
rect 2385 -692 2804 -654
rect 2385 -726 2759 -692
rect 2793 -726 2804 -692
rect 2385 -764 2804 -726
rect 2385 -798 2759 -764
rect 2793 -798 2804 -764
rect 2385 -836 2804 -798
rect 2385 -849 2759 -836
rect 2385 -883 2391 -849
rect 2425 -883 2649 -849
rect 2683 -870 2759 -849
rect 2793 -870 2804 -836
rect 2683 -883 2804 -870
rect 2385 -908 2804 -883
rect 2385 -921 2759 -908
rect 2385 -955 2391 -921
rect 2425 -955 2649 -921
rect 2683 -942 2759 -921
rect 2793 -942 2804 -908
rect 2683 -955 2804 -942
rect 2385 -980 2804 -955
rect 2385 -1014 2759 -980
rect 2793 -1014 2804 -980
rect 2385 -1049 2804 -1014
rect 2385 -1083 2484 -1049
rect 2518 -1083 2556 -1049
rect 2590 -1052 2804 -1049
rect 2590 -1083 2759 -1052
rect 2385 -1086 2759 -1083
rect 2793 -1086 2804 -1052
rect 2385 -1124 2804 -1086
rect 2385 -1158 2759 -1124
rect 2793 -1158 2804 -1124
rect 2385 -1185 2804 -1158
rect 2385 -1219 2484 -1185
rect 2518 -1219 2556 -1185
rect 2590 -1196 2804 -1185
rect 2590 -1219 2759 -1196
rect 2385 -1230 2759 -1219
rect 2793 -1230 2804 -1196
rect 2385 -1268 2804 -1230
rect 2385 -1302 2759 -1268
rect 2793 -1302 2804 -1268
rect 2385 -1313 2804 -1302
rect 2385 -1347 2391 -1313
rect 2425 -1347 2649 -1313
rect 2683 -1340 2804 -1313
rect 2683 -1347 2759 -1340
rect 2385 -1374 2759 -1347
rect 2793 -1374 2804 -1340
rect 2385 -1385 2804 -1374
rect 2385 -1419 2391 -1385
rect 2425 -1419 2649 -1385
rect 2683 -1412 2804 -1385
rect 2683 -1419 2759 -1412
rect 2385 -1446 2759 -1419
rect 2793 -1446 2804 -1412
rect 2385 -1484 2804 -1446
rect 2385 -1518 2759 -1484
rect 2793 -1518 2804 -1484
rect 2385 -1556 2804 -1518
rect 2385 -1590 2759 -1556
rect 2793 -1590 2804 -1556
rect 2385 -1616 2804 -1590
rect 2385 -1650 2391 -1616
rect 2425 -1650 2649 -1616
rect 2683 -1628 2804 -1616
rect 2683 -1650 2759 -1628
rect 2385 -1662 2759 -1650
rect 2793 -1662 2804 -1628
rect 2385 -1688 2804 -1662
rect 2385 -1722 2391 -1688
rect 2425 -1722 2649 -1688
rect 2683 -1700 2804 -1688
rect 2683 -1722 2759 -1700
rect 2385 -1734 2759 -1722
rect 2793 -1734 2804 -1700
rect 2385 -1772 2804 -1734
rect 2385 -1806 2759 -1772
rect 2793 -1806 2804 -1772
rect 2385 -1816 2804 -1806
rect 2385 -1850 2484 -1816
rect 2518 -1850 2556 -1816
rect 2590 -1844 2804 -1816
rect 2590 -1850 2759 -1844
rect 2385 -1878 2759 -1850
rect 2793 -1878 2804 -1844
rect 831 -1950 856 -1916
rect 890 -1950 1269 -1916
rect 831 -1952 1269 -1950
rect 2385 -1916 2804 -1878
rect 2385 -1950 2759 -1916
rect 2793 -1950 2804 -1916
rect 2385 -1952 2804 -1950
rect 831 -1958 2804 -1952
rect 831 -1988 1064 -1958
rect 831 -2022 856 -1988
rect 890 -1992 1064 -1988
rect 1098 -1992 1136 -1958
rect 1170 -1992 1516 -1958
rect 1550 -1992 1588 -1958
rect 1622 -1992 1774 -1958
rect 1808 -1992 1846 -1958
rect 1880 -1992 2032 -1958
rect 2066 -1992 2104 -1958
rect 2138 -1992 2484 -1958
rect 2518 -1992 2556 -1958
rect 2590 -1988 2804 -1958
rect 2590 -1992 2759 -1988
rect 890 -2022 2759 -1992
rect 2793 -2022 2804 -1988
rect 831 -2060 2804 -2022
rect 831 -2094 856 -2060
rect 890 -2086 2759 -2060
rect 890 -2094 971 -2086
rect 831 -2120 971 -2094
rect 1005 -2120 1229 -2086
rect 1263 -2120 1423 -2086
rect 1457 -2120 1681 -2086
rect 1715 -2120 1939 -2086
rect 1973 -2120 2197 -2086
rect 2231 -2120 2391 -2086
rect 2425 -2120 2649 -2086
rect 2683 -2094 2759 -2086
rect 2793 -2094 2804 -2060
rect 2683 -2120 2804 -2094
rect 831 -2132 2804 -2120
rect 831 -2166 856 -2132
rect 890 -2158 2759 -2132
rect 890 -2166 971 -2158
rect 831 -2192 971 -2166
rect 1005 -2192 1229 -2158
rect 1263 -2192 1423 -2158
rect 1457 -2192 1681 -2158
rect 1715 -2192 1939 -2158
rect 1973 -2192 2197 -2158
rect 2231 -2192 2391 -2158
rect 2425 -2192 2649 -2158
rect 2683 -2166 2759 -2158
rect 2793 -2166 2804 -2132
rect 2683 -2192 2804 -2166
rect 831 -2310 2804 -2192
rect 831 -2344 1002 -2310
rect 1036 -2344 1074 -2310
rect 1108 -2344 1146 -2310
rect 1180 -2344 1218 -2310
rect 1252 -2344 1290 -2310
rect 1324 -2344 1362 -2310
rect 1396 -2344 1434 -2310
rect 1468 -2344 1506 -2310
rect 1540 -2344 1578 -2310
rect 1612 -2344 1650 -2310
rect 1684 -2344 1722 -2310
rect 1756 -2344 1794 -2310
rect 1828 -2344 1866 -2310
rect 1900 -2344 1938 -2310
rect 1972 -2344 2010 -2310
rect 2044 -2344 2082 -2310
rect 2116 -2344 2154 -2310
rect 2188 -2344 2226 -2310
rect 2260 -2344 2298 -2310
rect 2332 -2344 2370 -2310
rect 2404 -2344 2442 -2310
rect 2476 -2344 2514 -2310
rect 2548 -2344 2586 -2310
rect 2620 -2344 2804 -2310
rect 831 -2369 2804 -2344
<< via1 >>
rect 1502 -316 1516 -306
rect 1516 -316 1550 -306
rect 1550 -316 1554 -306
rect 1502 -358 1554 -316
rect 1566 -316 1588 -306
rect 1588 -316 1618 -306
rect 1566 -358 1618 -316
rect 1630 -358 1682 -306
rect 1736 -316 1774 -306
rect 1774 -316 1788 -306
rect 1800 -316 1808 -306
rect 1808 -316 1846 -306
rect 1846 -316 1852 -306
rect 1864 -316 1880 -306
rect 1880 -316 1916 -306
rect 1736 -358 1788 -316
rect 1800 -358 1852 -316
rect 1864 -358 1916 -316
rect 1976 -358 2028 -306
rect 2040 -316 2066 -306
rect 2066 -316 2092 -306
rect 2040 -358 2092 -316
rect 2104 -316 2138 -306
rect 2138 -316 2156 -306
rect 2104 -358 2156 -316
rect 1502 -418 1554 -376
rect 1502 -428 1516 -418
rect 1516 -428 1550 -418
rect 1550 -428 1554 -418
rect 1566 -418 1618 -376
rect 1566 -428 1588 -418
rect 1588 -428 1618 -418
rect 1630 -428 1682 -376
rect 1736 -418 1788 -376
rect 1800 -418 1852 -376
rect 1864 -418 1916 -376
rect 1736 -428 1774 -418
rect 1774 -428 1788 -418
rect 1800 -428 1808 -418
rect 1808 -428 1846 -418
rect 1846 -428 1852 -418
rect 1864 -428 1880 -418
rect 1880 -428 1916 -418
rect 1976 -428 2028 -376
rect 2040 -418 2092 -376
rect 2040 -428 2066 -418
rect 2066 -428 2092 -418
rect 2104 -418 2156 -376
rect 2104 -428 2138 -418
rect 2138 -428 2156 -418
rect 1502 -1083 1516 -1073
rect 1516 -1083 1550 -1073
rect 1550 -1083 1554 -1073
rect 1502 -1125 1554 -1083
rect 1566 -1083 1588 -1073
rect 1588 -1083 1618 -1073
rect 1566 -1125 1618 -1083
rect 1630 -1125 1682 -1073
rect 1736 -1083 1774 -1073
rect 1774 -1083 1788 -1073
rect 1800 -1083 1808 -1073
rect 1808 -1083 1846 -1073
rect 1846 -1083 1852 -1073
rect 1864 -1083 1880 -1073
rect 1880 -1083 1916 -1073
rect 1736 -1125 1788 -1083
rect 1800 -1125 1852 -1083
rect 1864 -1125 1916 -1083
rect 1976 -1125 2028 -1073
rect 2040 -1083 2066 -1073
rect 2066 -1083 2092 -1073
rect 2040 -1125 2092 -1083
rect 2104 -1083 2138 -1073
rect 2138 -1083 2156 -1073
rect 2104 -1125 2156 -1083
rect 1502 -1185 1554 -1143
rect 1502 -1195 1516 -1185
rect 1516 -1195 1550 -1185
rect 1550 -1195 1554 -1185
rect 1566 -1185 1618 -1143
rect 1566 -1195 1588 -1185
rect 1588 -1195 1618 -1185
rect 1630 -1195 1682 -1143
rect 1736 -1185 1788 -1143
rect 1800 -1185 1852 -1143
rect 1864 -1185 1916 -1143
rect 1736 -1195 1774 -1185
rect 1774 -1195 1788 -1185
rect 1800 -1195 1808 -1185
rect 1808 -1195 1846 -1185
rect 1846 -1195 1852 -1185
rect 1864 -1195 1880 -1185
rect 1880 -1195 1916 -1185
rect 1976 -1195 2028 -1143
rect 2040 -1185 2092 -1143
rect 2040 -1195 2066 -1185
rect 2066 -1195 2092 -1185
rect 2104 -1185 2156 -1143
rect 2104 -1195 2138 -1185
rect 2138 -1195 2156 -1185
rect 1502 -1850 1516 -1818
rect 1516 -1850 1550 -1818
rect 1550 -1850 1554 -1818
rect 1502 -1870 1554 -1850
rect 1566 -1850 1588 -1818
rect 1588 -1850 1618 -1818
rect 1566 -1870 1618 -1850
rect 1630 -1870 1682 -1818
rect 1736 -1850 1774 -1818
rect 1774 -1850 1788 -1818
rect 1800 -1850 1808 -1818
rect 1808 -1850 1846 -1818
rect 1846 -1850 1852 -1818
rect 1864 -1850 1880 -1818
rect 1880 -1850 1916 -1818
rect 1736 -1870 1788 -1850
rect 1800 -1870 1852 -1850
rect 1864 -1870 1916 -1850
rect 1976 -1870 2028 -1818
rect 2040 -1850 2066 -1818
rect 2066 -1850 2092 -1818
rect 2040 -1870 2092 -1850
rect 2104 -1850 2138 -1818
rect 2138 -1850 2156 -1818
rect 2104 -1870 2156 -1850
<< metal2 >>
rect 1493 -306 2481 -298
rect 1493 -358 1502 -306
rect 1554 -358 1566 -306
rect 1618 -358 1630 -306
rect 1682 -358 1736 -306
rect 1788 -358 1800 -306
rect 1852 -358 1864 -306
rect 1916 -358 1976 -306
rect 2028 -358 2040 -306
rect 2092 -358 2104 -306
rect 2156 -339 2481 -306
rect 2156 -358 2221 -339
rect 1493 -376 2221 -358
rect 1493 -428 1502 -376
rect 1554 -428 1566 -376
rect 1618 -428 1630 -376
rect 1682 -428 1736 -376
rect 1788 -428 1800 -376
rect 1852 -428 1864 -376
rect 1916 -428 1976 -376
rect 2028 -428 2040 -376
rect 2092 -428 2104 -376
rect 2156 -395 2221 -376
rect 2277 -395 2301 -339
rect 2357 -395 2381 -339
rect 2437 -395 2481 -339
rect 2156 -428 2481 -395
rect 1493 -438 2481 -428
rect 1493 -1073 2481 -1065
rect 1493 -1125 1502 -1073
rect 1554 -1125 1566 -1073
rect 1618 -1125 1630 -1073
rect 1682 -1125 1736 -1073
rect 1788 -1125 1800 -1073
rect 1852 -1125 1864 -1073
rect 1916 -1125 1976 -1073
rect 2028 -1125 2040 -1073
rect 2092 -1125 2104 -1073
rect 2156 -1106 2481 -1073
rect 2156 -1125 2221 -1106
rect 1493 -1143 2221 -1125
rect 1493 -1195 1502 -1143
rect 1554 -1195 1566 -1143
rect 1618 -1195 1630 -1143
rect 1682 -1195 1736 -1143
rect 1788 -1195 1800 -1143
rect 1852 -1195 1864 -1143
rect 1916 -1195 1976 -1143
rect 2028 -1195 2040 -1143
rect 2092 -1195 2104 -1143
rect 2156 -1162 2221 -1143
rect 2277 -1162 2301 -1106
rect 2357 -1162 2381 -1106
rect 2437 -1162 2481 -1106
rect 2156 -1195 2481 -1162
rect 1493 -1205 2481 -1195
rect 1493 -1818 2481 -1810
rect 1493 -1870 1502 -1818
rect 1554 -1870 1566 -1818
rect 1618 -1870 1630 -1818
rect 1682 -1870 1736 -1818
rect 1788 -1870 1800 -1818
rect 1852 -1870 1864 -1818
rect 1916 -1870 1976 -1818
rect 2028 -1870 2040 -1818
rect 2092 -1870 2104 -1818
rect 2156 -1832 2481 -1818
rect 2156 -1870 2221 -1832
rect 1493 -1888 2221 -1870
rect 2277 -1888 2301 -1832
rect 2357 -1888 2381 -1832
rect 2437 -1888 2481 -1832
rect 1493 -1911 2481 -1888
<< via2 >>
rect 2221 -395 2277 -339
rect 2301 -395 2357 -339
rect 2381 -395 2437 -339
rect 2221 -1162 2277 -1106
rect 2301 -1162 2357 -1106
rect 2381 -1162 2437 -1106
rect 2221 -1888 2277 -1832
rect 2301 -1888 2357 -1832
rect 2381 -1888 2437 -1832
<< metal3 >>
rect 2181 -339 2481 -317
rect 2181 -395 2221 -339
rect 2277 -395 2301 -339
rect 2357 -395 2381 -339
rect 2437 -395 2481 -339
rect 2181 -1106 2481 -395
rect 2181 -1162 2221 -1106
rect 2277 -1162 2301 -1106
rect 2357 -1162 2381 -1106
rect 2437 -1162 2481 -1106
rect 2181 -1832 2481 -1162
rect 2181 -1888 2221 -1832
rect 2277 -1888 2301 -1832
rect 2357 -1888 2381 -1832
rect 2437 -1888 2481 -1832
rect 2181 -1911 2481 -1888
<< labels >>
flabel metal3 s 2227 -1811 2446 -458 2 FreeSans 3126 0 0 0 VB4
port 1 nsew
flabel metal1 s 877 -2094 1181 443 2 FreeSans 3126 0 0 0 AVDD
port 2 nsew
<< end >>
